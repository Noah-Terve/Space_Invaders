library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alien_sprite is
  port(
    clk : in std_logic;
    xaddr : in unsigned(8 downto 0);
    yaddr : in unsigned(7 downto 0);
	rgb : out std_logic_vector(5 downto 0)
  );
end alien_sprite;

architecture synth of alien_sprite is
    signal addr : std_logic_vector(16 downto 0);         
    begin
        process(clk) is begin
            if rising_edge(clk) then
                case addr is
                    when "00000000000000000" => rgb <= "000000";
					when "00000000000000001" => rgb <= "000000";
					when "00000000000000010" => rgb <= "000000";
					when "00000000000000011" => rgb <= "000000";
					when "00000000000000100" => rgb <= "000000";
					when "00000000000000101" => rgb <= "000000";
					when "00000000000000110" => rgb <= "000000";
					when "00000000000000111" => rgb <= "000000";
					when "00000000000001000" => rgb <= "000000";
					when "00000000000001001" => rgb <= "000000";
					when "00000000000001010" => rgb <= "000000";
					when "00000000000001011" => rgb <= "000000";
					when "00000000000001100" => rgb <= "000000";
					when "00000000000001101" => rgb <= "000000";
					when "00000000000001110" => rgb <= "000000";
					when "00000000000001111" => rgb <= "000000";
					when "00000000000010000" => rgb <= "000000";
					when "00000000000010001" => rgb <= "000000";
					when "00000000000010010" => rgb <= "000000";
					when "00000000000010011" => rgb <= "000000";
					when "00000000000010100" => rgb <= "000000";
					when "00000000000010101" => rgb <= "000000";
					when "00000000000010110" => rgb <= "000000";
					when "00000000000010111" => rgb <= "000000";
					when "00000000000011000" => rgb <= "000000";
					when "00000000000011001" => rgb <= "000000";
					when "00000000000011010" => rgb <= "000000";
					when "00000000000011011" => rgb <= "000000";
					when "00000000000011100" => rgb <= "000000";
					when "00000000000011101" => rgb <= "000000";
					when "00000000000011110" => rgb <= "000000";
					when "00000000000011111" => rgb <= "000000";
					when "00000000000100000" => rgb <= "000000";
					when "00000000000100001" => rgb <= "000000";
					when "00000000000100010" => rgb <= "000000";
					when "00000000000100011" => rgb <= "000000";
					when "00000000000100100" => rgb <= "000000";
					when "00000000000100101" => rgb <= "000000";
					when "00000000000100110" => rgb <= "000000";
					when "00000000000100111" => rgb <= "000000";
					when "00000000000101000" => rgb <= "000000";
					when "00000000000101001" => rgb <= "000000";
					when "00000000000101010" => rgb <= "000000";
					when "00000000000101011" => rgb <= "000000";
					when "00000000000101100" => rgb <= "000000";
					when "00000000000101101" => rgb <= "000000";
					when "00000000000101110" => rgb <= "000000";
					when "00000000000101111" => rgb <= "000000";
					when "00000000000110000" => rgb <= "000000";
					when "00000000000110001" => rgb <= "000000";
					when "00000000000110010" => rgb <= "000000";
					when "00000000000110011" => rgb <= "000000";
					when "00000000000110100" => rgb <= "000000";
					when "00000000000110101" => rgb <= "000000";
					when "00000000000110110" => rgb <= "000000";
					when "00000000000110111" => rgb <= "000000";
					when "00000000000111000" => rgb <= "000000";
					when "00000000000111001" => rgb <= "000000";
					when "00000000000111010" => rgb <= "000000";
					when "00000000000111011" => rgb <= "000000";
					when "00000000000111100" => rgb <= "000000";
					when "00000000000111101" => rgb <= "000000";
					when "00000000000111110" => rgb <= "000000";
					when "00000000000111111" => rgb <= "000000";
					when "00000000001000000" => rgb <= "000000";
					when "00000000001000001" => rgb <= "000000";
					when "00000000001000010" => rgb <= "000000";
					when "00000000001000011" => rgb <= "000000";
					when "00000000001000100" => rgb <= "000000";
					when "00000000001000101" => rgb <= "000000";
					when "00000000001000110" => rgb <= "000000";
					when "00000000001000111" => rgb <= "000000";
					when "00000000001001000" => rgb <= "000000";
					when "00000000001001001" => rgb <= "000000";
					when "00000000001001010" => rgb <= "000000";
					when "00000000001001011" => rgb <= "000000";
					when "00000000001001100" => rgb <= "000000";
					when "00000000001001101" => rgb <= "000000";
					when "00000000001001110" => rgb <= "000000";
					when "00000000001001111" => rgb <= "000000";
					when "00000000001010000" => rgb <= "000000";
					when "00000000001010001" => rgb <= "000000";
					when "00000000001010010" => rgb <= "000000";
					when "00000000001010011" => rgb <= "000000";
					when "00000000001010100" => rgb <= "000000";
					when "00000000001010101" => rgb <= "000000";
					when "00000000001010110" => rgb <= "000000";
					when "00000000001010111" => rgb <= "000000";
					when "00000000001011000" => rgb <= "000000";
					when "00000000001011001" => rgb <= "000000";
					when "00000000001011010" => rgb <= "000000";
					when "00000000001011011" => rgb <= "000000";
					when "00000000001011100" => rgb <= "000000";
					when "00000000001011101" => rgb <= "000000";
					when "00000000001011110" => rgb <= "000000";
					when "00000000001011111" => rgb <= "000000";
					when "00000000001100000" => rgb <= "000000";
					when "00000000001100001" => rgb <= "000000";
					when "00000000001100010" => rgb <= "000000";
					when "00000000001100011" => rgb <= "000000";
					when "00000000001100100" => rgb <= "000000";
					when "00000000001100101" => rgb <= "000000";
					when "00000000001100110" => rgb <= "000000";
					when "00000000001100111" => rgb <= "000000";
					when "00000000001101000" => rgb <= "000000";
					when "00000000001101001" => rgb <= "000000";
					when "00000000001101010" => rgb <= "000000";
					when "00000000001101011" => rgb <= "000000";
					when "00000000001101100" => rgb <= "000000";
					when "00000000001101101" => rgb <= "000000";
					when "00000000001101110" => rgb <= "000000";
					when "00000000001101111" => rgb <= "000000";
					when "00000000001110000" => rgb <= "000000";
					when "00000000001110001" => rgb <= "000000";
					when "00000000001110010" => rgb <= "000000";
					when "00000000001110011" => rgb <= "000000";
					when "00000000001110100" => rgb <= "000000";
					when "00000000001110101" => rgb <= "000000";
					when "00000000001110110" => rgb <= "000000";
					when "00000000001110111" => rgb <= "000000";
					when "00000000001111000" => rgb <= "000000";
					when "00000000001111001" => rgb <= "000000";
					when "00000000001111010" => rgb <= "000000";
					when "00000000001111011" => rgb <= "000000";
					when "00000000001111100" => rgb <= "000000";
					when "00000000001111101" => rgb <= "000000";
					when "00000000001111110" => rgb <= "000000";
					when "00000000001111111" => rgb <= "000000";
					when "00000000010000000" => rgb <= "000000";
					when "00000000010000001" => rgb <= "000000";
					when "00000000010000010" => rgb <= "000000";
					when "00000000010000011" => rgb <= "000000";
					when "00000000010000100" => rgb <= "000000";
					when "00000000010000101" => rgb <= "000000";
					when "00000000010000110" => rgb <= "000000";
					when "00000000010000111" => rgb <= "000000";
					when "00000000010001000" => rgb <= "000000";
					when "00000000010001001" => rgb <= "000000";
					when "00000000010001010" => rgb <= "000000";
					when "00000000010001011" => rgb <= "000000";
					when "00000000010001100" => rgb <= "000000";
					when "00000000010001101" => rgb <= "000000";
					when "00000000010001110" => rgb <= "000000";
					when "00000000010001111" => rgb <= "000000";
					when "00000000010010000" => rgb <= "000000";
					when "00000000010010001" => rgb <= "000000";
					when "00000000010010010" => rgb <= "000000";
					when "00000000010010011" => rgb <= "000000";
					when "00000000010010100" => rgb <= "000000";
					when "00000000010010101" => rgb <= "000000";
					when "00000000010010110" => rgb <= "000000";
					when "00000000010010111" => rgb <= "000000";
					when "00000000010011000" => rgb <= "000000";
					when "00000000010011001" => rgb <= "000000";
					when "00000000010011010" => rgb <= "000000";
					when "00000000010011011" => rgb <= "000000";
					when "00000000010011100" => rgb <= "000000";
					when "00000000010011101" => rgb <= "000000";
					when "00000000010011110" => rgb <= "000000";
					when "00000000010011111" => rgb <= "000000";
					when "00000000010100000" => rgb <= "000000";
					when "00000000010100001" => rgb <= "000000";
					when "00000000010100010" => rgb <= "000000";
					when "00000000010100011" => rgb <= "000000";
					when "00000000010100100" => rgb <= "000000";
					when "00000000010100101" => rgb <= "000000";
					when "00000000010100110" => rgb <= "000000";
					when "00000000010100111" => rgb <= "000000";
					when "00000000010101000" => rgb <= "000000";
					when "00000000010101001" => rgb <= "000000";
					when "00000000010101010" => rgb <= "000000";
					when "00000000010101011" => rgb <= "000000";
					when "00000000010101100" => rgb <= "000000";
					when "00000000010101101" => rgb <= "000000";
					when "00000000010101110" => rgb <= "000000";
					when "00000000010101111" => rgb <= "000000";
					when "00000000010110000" => rgb <= "000000";
					when "00000000010110001" => rgb <= "000000";
					when "00000000010110010" => rgb <= "000000";
					when "00000000010110011" => rgb <= "000000";
					when "00000000010110100" => rgb <= "000000";
					when "00000000010110101" => rgb <= "000000";
					when "00000000010110110" => rgb <= "000000";
					when "00000000010110111" => rgb <= "000000";
					when "00000000010111000" => rgb <= "000000";
					when "00000000010111001" => rgb <= "000000";
					when "00000000010111010" => rgb <= "000000";
					when "00000000010111011" => rgb <= "000000";
					when "00000000010111100" => rgb <= "000000";
					when "00000000010111101" => rgb <= "000000";
					when "00000000010111110" => rgb <= "000000";
					when "00000000010111111" => rgb <= "000000";
					when "00000000011000000" => rgb <= "000000";
					when "00000000011000001" => rgb <= "000000";
					when "00000000011000010" => rgb <= "000000";
					when "00000000011000011" => rgb <= "000000";
					when "00000000011000100" => rgb <= "000000";
					when "00000000011000101" => rgb <= "000000";
					when "00000000011000110" => rgb <= "000000";
					when "00000000011000111" => rgb <= "000000";
					when "00000000011001000" => rgb <= "000000";
					when "00000000011001001" => rgb <= "000000";
					when "00000000011001010" => rgb <= "000000";
					when "00000000011001011" => rgb <= "000000";
					when "00000000011001100" => rgb <= "000000";
					when "00000000011001101" => rgb <= "000000";
					when "00000000011001110" => rgb <= "000000";
					when "00000000011001111" => rgb <= "000000";
					when "00000000011010000" => rgb <= "000000";
					when "00000000011010001" => rgb <= "000000";
					when "00000000011010010" => rgb <= "000000";
					when "00000000011010011" => rgb <= "000000";
					when "00000000011010100" => rgb <= "000000";
					when "00000000011010101" => rgb <= "000000";
					when "00000000011010110" => rgb <= "000000";
					when "00000000011010111" => rgb <= "000000";
					when "00000000011011000" => rgb <= "000000";
					when "00000000011011001" => rgb <= "000000";
					when "00000000011011010" => rgb <= "000000";
					when "00000000011011011" => rgb <= "000000";
					when "00000000011011100" => rgb <= "000000";
					when "00000000011011101" => rgb <= "000000";
					when "00000000011011110" => rgb <= "000000";
					when "00000000011011111" => rgb <= "000000";
					when "00000000011100000" => rgb <= "000000";
					when "00000000011100001" => rgb <= "000000";
					when "00000000011100010" => rgb <= "000000";
					when "00000000011100011" => rgb <= "000000";
					when "00000000011100100" => rgb <= "000000";
					when "00000000011100101" => rgb <= "000000";
					when "00000000011100110" => rgb <= "000000";
					when "00000000011100111" => rgb <= "000000";
					when "00000000011101000" => rgb <= "000000";
					when "00000000011101001" => rgb <= "000000";
					when "00000000011101010" => rgb <= "000000";
					when "00000000011101011" => rgb <= "000000";
					when "00000000011101100" => rgb <= "000000";
					when "00000000011101101" => rgb <= "000000";
					when "00000000011101110" => rgb <= "000000";
					when "00000000011101111" => rgb <= "000000";
					when "00000000011110000" => rgb <= "000000";
					when "00000000011110001" => rgb <= "000000";
					when "00000000011110010" => rgb <= "000000";
					when "00000000011110011" => rgb <= "000000";
					when "00000000011110100" => rgb <= "000000";
					when "00000000011110101" => rgb <= "000000";
					when "00000000011110110" => rgb <= "000000";
					when "00000000011110111" => rgb <= "000000";
					when "00000000011111000" => rgb <= "000000";
					when "00000000011111001" => rgb <= "000000";
					when "00000000011111010" => rgb <= "000000";
					when "00000000011111011" => rgb <= "000000";
					when "00000000011111100" => rgb <= "000000";
					when "00000000011111101" => rgb <= "000000";
					when "00000000011111110" => rgb <= "000000";
					when "00000000011111111" => rgb <= "000000";
					when "00000000100000000" => rgb <= "000000";
					when "00000000100000001" => rgb <= "000000";
					when "00000000100000010" => rgb <= "000000";
					when "00000000100000011" => rgb <= "000000";
					when "00000000100000100" => rgb <= "000000";
					when "00000000100000101" => rgb <= "000000";
					when "00000000100000110" => rgb <= "000000";
					when "00000000100000111" => rgb <= "000000";
					when "00000000100001000" => rgb <= "000000";
					when "00000000100001001" => rgb <= "000000";
					when "00000000100001010" => rgb <= "000000";
					when "00000000100001011" => rgb <= "000000";
					when "00000000100001100" => rgb <= "000000";
					when "00000000100001101" => rgb <= "000000";
					when "00000000100001110" => rgb <= "000000";
					when "00000000100001111" => rgb <= "000000";
					when "00000000100010000" => rgb <= "000000";
					when "00000000100010001" => rgb <= "000000";
					when "00000000100010010" => rgb <= "000000";
					when "00000000100010011" => rgb <= "000000";
					when "00000000100010100" => rgb <= "000000";
					when "00000000100010101" => rgb <= "000000";
					when "00000000100010110" => rgb <= "000000";
					when "00000000100010111" => rgb <= "000000";
					when "00000000100011000" => rgb <= "000000";
					when "00000000100011001" => rgb <= "000000";
					when "00000000100011010" => rgb <= "000000";
					when "00000000100011011" => rgb <= "000000";
					when "00000000100011100" => rgb <= "000000";
					when "00000000100011101" => rgb <= "000000";
					when "00000000100011110" => rgb <= "000000";
					when "00000000100011111" => rgb <= "000000";
					when "00000000100100000" => rgb <= "000000";
					when "00000000100100001" => rgb <= "000000";
					when "00000000100100010" => rgb <= "000000";
					when "00000000100100011" => rgb <= "000000";
					when "00000000100100100" => rgb <= "000000";
					when "00000000100100101" => rgb <= "000000";
					when "00000000100100110" => rgb <= "000000";
					when "00000000100100111" => rgb <= "000000";
					when "00000000100101000" => rgb <= "000000";
					when "00000000100101001" => rgb <= "000000";
					when "00000000100101010" => rgb <= "000000";
					when "00000000100101011" => rgb <= "000000";
					when "00000000100101100" => rgb <= "000000";
					when "00000000100101101" => rgb <= "000000";
					when "00000000100101110" => rgb <= "000000";
					when "00000000100101111" => rgb <= "000000";
					when "00000000100110000" => rgb <= "000000";
					when "00000000100110001" => rgb <= "000000";
					when "00000000100110010" => rgb <= "000000";
					when "00000000100110011" => rgb <= "000000";
					when "00000000100110100" => rgb <= "000000";
					when "00000000100110101" => rgb <= "000000";
					when "00000000100110110" => rgb <= "000000";
					when "00000000100110111" => rgb <= "000000";
					when "00000000100111000" => rgb <= "000000";
					when "00000000100111001" => rgb <= "000000";
					when "00000000100111010" => rgb <= "000000";
					when "00000000100111011" => rgb <= "000000";
					when "00000000100111100" => rgb <= "000000";
					when "00000000100111101" => rgb <= "000000";
					when "00000000100111110" => rgb <= "000000";
					when "00000000100111111" => rgb <= "000000";
					when "00000001000000000" => rgb <= "000000";
					when "00000001000000001" => rgb <= "000000";
					when "00000001000000010" => rgb <= "000000";
					when "00000001000000011" => rgb <= "000000";
					when "00000001000000100" => rgb <= "000000";
					when "00000001000000101" => rgb <= "000000";
					when "00000001000000110" => rgb <= "000000";
					when "00000001000000111" => rgb <= "000000";
					when "00000001000001000" => rgb <= "000000";
					when "00000001000001001" => rgb <= "000000";
					when "00000001000001010" => rgb <= "000000";
					when "00000001000001011" => rgb <= "000000";
					when "00000001000001100" => rgb <= "000000";
					when "00000001000001101" => rgb <= "000000";
					when "00000001000001110" => rgb <= "000000";
					when "00000001000001111" => rgb <= "000000";
					when "00000001000010000" => rgb <= "000000";
					when "00000001000010001" => rgb <= "000000";
					when "00000001000010010" => rgb <= "000000";
					when "00000001000010011" => rgb <= "000000";
					when "00000001000010100" => rgb <= "000000";
					when "00000001000010101" => rgb <= "000000";
					when "00000001000010110" => rgb <= "000000";
					when "00000001000010111" => rgb <= "000000";
					when "00000001000011000" => rgb <= "000000";
					when "00000001000011001" => rgb <= "000000";
					when "00000001000011010" => rgb <= "000000";
					when "00000001000011011" => rgb <= "000000";
					when "00000001000011100" => rgb <= "000000";
					when "00000001000011101" => rgb <= "000000";
					when "00000001000011110" => rgb <= "000000";
					when "00000001000011111" => rgb <= "000000";
					when "00000001000100000" => rgb <= "000000";
					when "00000001000100001" => rgb <= "000000";
					when "00000001000100010" => rgb <= "000000";
					when "00000001000100011" => rgb <= "000000";
					when "00000001000100100" => rgb <= "000000";
					when "00000001000100101" => rgb <= "000000";
					when "00000001000100110" => rgb <= "000000";
					when "00000001000100111" => rgb <= "000000";
					when "00000001000101000" => rgb <= "000000";
					when "00000001000101001" => rgb <= "000000";
					when "00000001000101010" => rgb <= "000000";
					when "00000001000101011" => rgb <= "000000";
					when "00000001000101100" => rgb <= "000000";
					when "00000001000101101" => rgb <= "000000";
					when "00000001000101110" => rgb <= "000000";
					when "00000001000101111" => rgb <= "000000";
					when "00000001000110000" => rgb <= "000000";
					when "00000001000110001" => rgb <= "000000";
					when "00000001000110010" => rgb <= "000000";
					when "00000001000110011" => rgb <= "000000";
					when "00000001000110100" => rgb <= "000000";
					when "00000001000110101" => rgb <= "000000";
					when "00000001000110110" => rgb <= "000000";
					when "00000001000110111" => rgb <= "000000";
					when "00000001000111000" => rgb <= "000000";
					when "00000001000111001" => rgb <= "000000";
					when "00000001000111010" => rgb <= "000000";
					when "00000001000111011" => rgb <= "000000";
					when "00000001000111100" => rgb <= "000000";
					when "00000001000111101" => rgb <= "000000";
					when "00000001000111110" => rgb <= "000000";
					when "00000001000111111" => rgb <= "000000";
					when "00000001001000000" => rgb <= "000000";
					when "00000001001000001" => rgb <= "000000";
					when "00000001001000010" => rgb <= "000000";
					when "00000001001000011" => rgb <= "000000";
					when "00000001001000100" => rgb <= "000000";
					when "00000001001000101" => rgb <= "000000";
					when "00000001001000110" => rgb <= "000000";
					when "00000001001000111" => rgb <= "000000";
					when "00000001001001000" => rgb <= "000000";
					when "00000001001001001" => rgb <= "000000";
					when "00000001001001010" => rgb <= "000000";
					when "00000001001001011" => rgb <= "000000";
					when "00000001001001100" => rgb <= "000000";
					when "00000001001001101" => rgb <= "000000";
					when "00000001001001110" => rgb <= "000000";
					when "00000001001001111" => rgb <= "000000";
					when "00000001001010000" => rgb <= "000000";
					when "00000001001010001" => rgb <= "000000";
					when "00000001001010010" => rgb <= "000000";
					when "00000001001010011" => rgb <= "000000";
					when "00000001001010100" => rgb <= "000000";
					when "00000001001010101" => rgb <= "000000";
					when "00000001001010110" => rgb <= "000000";
					when "00000001001010111" => rgb <= "000000";
					when "00000001001011000" => rgb <= "000000";
					when "00000001001011001" => rgb <= "000000";
					when "00000001001011010" => rgb <= "000000";
					when "00000001001011011" => rgb <= "000000";
					when "00000001001011100" => rgb <= "000000";
					when "00000001001011101" => rgb <= "000000";
					when "00000001001011110" => rgb <= "000000";
					when "00000001001011111" => rgb <= "000000";
					when "00000001001100000" => rgb <= "000000";
					when "00000001001100001" => rgb <= "000000";
					when "00000001001100010" => rgb <= "000000";
					when "00000001001100011" => rgb <= "000000";
					when "00000001001100100" => rgb <= "000000";
					when "00000001001100101" => rgb <= "000000";
					when "00000001001100110" => rgb <= "000000";
					when "00000001001100111" => rgb <= "000000";
					when "00000001001101000" => rgb <= "000000";
					when "00000001001101001" => rgb <= "000000";
					when "00000001001101010" => rgb <= "000000";
					when "00000001001101011" => rgb <= "000000";
					when "00000001001101100" => rgb <= "000000";
					when "00000001001101101" => rgb <= "000000";
					when "00000001001101110" => rgb <= "000000";
					when "00000001001101111" => rgb <= "000000";
					when "00000001001110000" => rgb <= "000000";
					when "00000001001110001" => rgb <= "000000";
					when "00000001001110010" => rgb <= "000000";
					when "00000001001110011" => rgb <= "000000";
					when "00000001001110100" => rgb <= "000000";
					when "00000001001110101" => rgb <= "000000";
					when "00000001001110110" => rgb <= "000000";
					when "00000001001110111" => rgb <= "000000";
					when "00000001001111000" => rgb <= "000000";
					when "00000001001111001" => rgb <= "000000";
					when "00000001001111010" => rgb <= "000000";
					when "00000001001111011" => rgb <= "000000";
					when "00000001001111100" => rgb <= "000000";
					when "00000001001111101" => rgb <= "000000";
					when "00000001001111110" => rgb <= "000000";
					when "00000001001111111" => rgb <= "000000";
					when "00000001010000000" => rgb <= "000000";
					when "00000001010000001" => rgb <= "000000";
					when "00000001010000010" => rgb <= "000000";
					when "00000001010000011" => rgb <= "000000";
					when "00000001010000100" => rgb <= "000000";
					when "00000001010000101" => rgb <= "000000";
					when "00000001010000110" => rgb <= "000000";
					when "00000001010000111" => rgb <= "000000";
					when "00000001010001000" => rgb <= "000000";
					when "00000001010001001" => rgb <= "000000";
					when "00000001010001010" => rgb <= "000000";
					when "00000001010001011" => rgb <= "000000";
					when "00000001010001100" => rgb <= "000000";
					when "00000001010001101" => rgb <= "000000";
					when "00000001010001110" => rgb <= "000000";
					when "00000001010001111" => rgb <= "000000";
					when "00000001010010000" => rgb <= "000000";
					when "00000001010010001" => rgb <= "000000";
					when "00000001010010010" => rgb <= "000000";
					when "00000001010010011" => rgb <= "000000";
					when "00000001010010100" => rgb <= "000000";
					when "00000001010010101" => rgb <= "000000";
					when "00000001010010110" => rgb <= "000000";
					when "00000001010010111" => rgb <= "000000";
					when "00000001010011000" => rgb <= "000000";
					when "00000001010011001" => rgb <= "000000";
					when "00000001010011010" => rgb <= "000000";
					when "00000001010011011" => rgb <= "000000";
					when "00000001010011100" => rgb <= "000000";
					when "00000001010011101" => rgb <= "000000";
					when "00000001010011110" => rgb <= "000000";
					when "00000001010011111" => rgb <= "000000";
					when "00000001010100000" => rgb <= "000000";
					when "00000001010100001" => rgb <= "000000";
					when "00000001010100010" => rgb <= "000000";
					when "00000001010100011" => rgb <= "000000";
					when "00000001010100100" => rgb <= "000000";
					when "00000001010100101" => rgb <= "000000";
					when "00000001010100110" => rgb <= "000000";
					when "00000001010100111" => rgb <= "000000";
					when "00000001010101000" => rgb <= "000000";
					when "00000001010101001" => rgb <= "000000";
					when "00000001010101010" => rgb <= "000000";
					when "00000001010101011" => rgb <= "000000";
					when "00000001010101100" => rgb <= "000000";
					when "00000001010101101" => rgb <= "000000";
					when "00000001010101110" => rgb <= "000000";
					when "00000001010101111" => rgb <= "000000";
					when "00000001010110000" => rgb <= "000000";
					when "00000001010110001" => rgb <= "000000";
					when "00000001010110010" => rgb <= "000000";
					when "00000001010110011" => rgb <= "000000";
					when "00000001010110100" => rgb <= "000000";
					when "00000001010110101" => rgb <= "000000";
					when "00000001010110110" => rgb <= "000000";
					when "00000001010110111" => rgb <= "000000";
					when "00000001010111000" => rgb <= "000000";
					when "00000001010111001" => rgb <= "000000";
					when "00000001010111010" => rgb <= "000000";
					when "00000001010111011" => rgb <= "000000";
					when "00000001010111100" => rgb <= "000000";
					when "00000001010111101" => rgb <= "000000";
					when "00000001010111110" => rgb <= "000000";
					when "00000001010111111" => rgb <= "000000";
					when "00000001011000000" => rgb <= "000000";
					when "00000001011000001" => rgb <= "000000";
					when "00000001011000010" => rgb <= "000000";
					when "00000001011000011" => rgb <= "000000";
					when "00000001011000100" => rgb <= "000000";
					when "00000001011000101" => rgb <= "000000";
					when "00000001011000110" => rgb <= "000000";
					when "00000001011000111" => rgb <= "000000";
					when "00000001011001000" => rgb <= "000000";
					when "00000001011001001" => rgb <= "000000";
					when "00000001011001010" => rgb <= "000000";
					when "00000001011001011" => rgb <= "000000";
					when "00000001011001100" => rgb <= "000000";
					when "00000001011001101" => rgb <= "000000";
					when "00000001011001110" => rgb <= "000000";
					when "00000001011001111" => rgb <= "000000";
					when "00000001011010000" => rgb <= "000000";
					when "00000001011010001" => rgb <= "000000";
					when "00000001011010010" => rgb <= "000000";
					when "00000001011010011" => rgb <= "000000";
					when "00000001011010100" => rgb <= "000000";
					when "00000001011010101" => rgb <= "000000";
					when "00000001011010110" => rgb <= "000000";
					when "00000001011010111" => rgb <= "000000";
					when "00000001011011000" => rgb <= "000000";
					when "00000001011011001" => rgb <= "000000";
					when "00000001011011010" => rgb <= "000000";
					when "00000001011011011" => rgb <= "000000";
					when "00000001011011100" => rgb <= "000000";
					when "00000001011011101" => rgb <= "000000";
					when "00000001011011110" => rgb <= "000000";
					when "00000001011011111" => rgb <= "000000";
					when "00000001011100000" => rgb <= "000000";
					when "00000001011100001" => rgb <= "000000";
					when "00000001011100010" => rgb <= "000000";
					when "00000001011100011" => rgb <= "000000";
					when "00000001011100100" => rgb <= "000000";
					when "00000001011100101" => rgb <= "000000";
					when "00000001011100110" => rgb <= "000000";
					when "00000001011100111" => rgb <= "000000";
					when "00000001011101000" => rgb <= "000000";
					when "00000001011101001" => rgb <= "000000";
					when "00000001011101010" => rgb <= "000000";
					when "00000001011101011" => rgb <= "000000";
					when "00000001011101100" => rgb <= "000000";
					when "00000001011101101" => rgb <= "000000";
					when "00000001011101110" => rgb <= "000000";
					when "00000001011101111" => rgb <= "000000";
					when "00000001011110000" => rgb <= "000000";
					when "00000001011110001" => rgb <= "000000";
					when "00000001011110010" => rgb <= "000000";
					when "00000001011110011" => rgb <= "000000";
					when "00000001011110100" => rgb <= "000000";
					when "00000001011110101" => rgb <= "000000";
					when "00000001011110110" => rgb <= "000000";
					when "00000001011110111" => rgb <= "000000";
					when "00000001011111000" => rgb <= "000000";
					when "00000001011111001" => rgb <= "000000";
					when "00000001011111010" => rgb <= "000000";
					when "00000001011111011" => rgb <= "000000";
					when "00000001011111100" => rgb <= "000000";
					when "00000001011111101" => rgb <= "000000";
					when "00000001011111110" => rgb <= "000000";
					when "00000001011111111" => rgb <= "000000";
					when "00000001100000000" => rgb <= "000000";
					when "00000001100000001" => rgb <= "000000";
					when "00000001100000010" => rgb <= "000000";
					when "00000001100000011" => rgb <= "000000";
					when "00000001100000100" => rgb <= "000000";
					when "00000001100000101" => rgb <= "000000";
					when "00000001100000110" => rgb <= "000000";
					when "00000001100000111" => rgb <= "000000";
					when "00000001100001000" => rgb <= "000000";
					when "00000001100001001" => rgb <= "000000";
					when "00000001100001010" => rgb <= "000000";
					when "00000001100001011" => rgb <= "000000";
					when "00000001100001100" => rgb <= "000000";
					when "00000001100001101" => rgb <= "000000";
					when "00000001100001110" => rgb <= "000000";
					when "00000001100001111" => rgb <= "000000";
					when "00000001100010000" => rgb <= "000000";
					when "00000001100010001" => rgb <= "000000";
					when "00000001100010010" => rgb <= "000000";
					when "00000001100010011" => rgb <= "000000";
					when "00000001100010100" => rgb <= "000000";
					when "00000001100010101" => rgb <= "000000";
					when "00000001100010110" => rgb <= "000000";
					when "00000001100010111" => rgb <= "000000";
					when "00000001100011000" => rgb <= "000000";
					when "00000001100011001" => rgb <= "000000";
					when "00000001100011010" => rgb <= "000000";
					when "00000001100011011" => rgb <= "000000";
					when "00000001100011100" => rgb <= "000000";
					when "00000001100011101" => rgb <= "000000";
					when "00000001100011110" => rgb <= "000000";
					when "00000001100011111" => rgb <= "000000";
					when "00000001100100000" => rgb <= "000000";
					when "00000001100100001" => rgb <= "000000";
					when "00000001100100010" => rgb <= "000000";
					when "00000001100100011" => rgb <= "000000";
					when "00000001100100100" => rgb <= "000000";
					when "00000001100100101" => rgb <= "000000";
					when "00000001100100110" => rgb <= "000000";
					when "00000001100100111" => rgb <= "000000";
					when "00000001100101000" => rgb <= "000000";
					when "00000001100101001" => rgb <= "000000";
					when "00000001100101010" => rgb <= "000000";
					when "00000001100101011" => rgb <= "000000";
					when "00000001100101100" => rgb <= "000000";
					when "00000001100101101" => rgb <= "000000";
					when "00000001100101110" => rgb <= "000000";
					when "00000001100101111" => rgb <= "000000";
					when "00000001100110000" => rgb <= "000000";
					when "00000001100110001" => rgb <= "000000";
					when "00000001100110010" => rgb <= "000000";
					when "00000001100110011" => rgb <= "000000";
					when "00000001100110100" => rgb <= "000000";
					when "00000001100110101" => rgb <= "000000";
					when "00000001100110110" => rgb <= "000000";
					when "00000001100110111" => rgb <= "000000";
					when "00000001100111000" => rgb <= "000000";
					when "00000001100111001" => rgb <= "000000";
					when "00000001100111010" => rgb <= "000000";
					when "00000001100111011" => rgb <= "000000";
					when "00000001100111100" => rgb <= "000000";
					when "00000001100111101" => rgb <= "000000";
					when "00000001100111110" => rgb <= "000000";
					when "00000001100111111" => rgb <= "000000";
					when "00000010000000000" => rgb <= "000000";
					when "00000010000000001" => rgb <= "000000";
					when "00000010000000010" => rgb <= "000000";
					when "00000010000000011" => rgb <= "000000";
					when "00000010000000100" => rgb <= "000000";
					when "00000010000000101" => rgb <= "000000";
					when "00000010000000110" => rgb <= "000000";
					when "00000010000000111" => rgb <= "000000";
					when "00000010000001000" => rgb <= "000000";
					when "00000010000001001" => rgb <= "000000";
					when "00000010000001010" => rgb <= "000000";
					when "00000010000001011" => rgb <= "000000";
					when "00000010000001100" => rgb <= "000000";
					when "00000010000001101" => rgb <= "000000";
					when "00000010000001110" => rgb <= "000000";
					when "00000010000001111" => rgb <= "000000";
					when "00000010000010000" => rgb <= "000000";
					when "00000010000010001" => rgb <= "000000";
					when "00000010000010010" => rgb <= "000000";
					when "00000010000010011" => rgb <= "000000";
					when "00000010000010100" => rgb <= "000000";
					when "00000010000010101" => rgb <= "000000";
					when "00000010000010110" => rgb <= "000000";
					when "00000010000010111" => rgb <= "000000";
					when "00000010000011000" => rgb <= "000000";
					when "00000010000011001" => rgb <= "000000";
					when "00000010000011010" => rgb <= "000000";
					when "00000010000011011" => rgb <= "000000";
					when "00000010000011100" => rgb <= "000000";
					when "00000010000011101" => rgb <= "000000";
					when "00000010000011110" => rgb <= "000000";
					when "00000010000011111" => rgb <= "000000";
					when "00000010000100000" => rgb <= "000000";
					when "00000010000100001" => rgb <= "000000";
					when "00000010000100010" => rgb <= "000000";
					when "00000010000100011" => rgb <= "000000";
					when "00000010000100100" => rgb <= "000000";
					when "00000010000100101" => rgb <= "000000";
					when "00000010000100110" => rgb <= "000000";
					when "00000010000100111" => rgb <= "000000";
					when "00000010000101000" => rgb <= "000000";
					when "00000010000101001" => rgb <= "000000";
					when "00000010000101010" => rgb <= "000000";
					when "00000010000101011" => rgb <= "000000";
					when "00000010000101100" => rgb <= "000000";
					when "00000010000101101" => rgb <= "000000";
					when "00000010000101110" => rgb <= "000000";
					when "00000010000101111" => rgb <= "000000";
					when "00000010000110000" => rgb <= "000000";
					when "00000010000110001" => rgb <= "000000";
					when "00000010000110010" => rgb <= "000000";
					when "00000010000110011" => rgb <= "000000";
					when "00000010000110100" => rgb <= "000000";
					when "00000010000110101" => rgb <= "000000";
					when "00000010000110110" => rgb <= "000000";
					when "00000010000110111" => rgb <= "000000";
					when "00000010000111000" => rgb <= "000000";
					when "00000010000111001" => rgb <= "000000";
					when "00000010000111010" => rgb <= "000000";
					when "00000010000111011" => rgb <= "000000";
					when "00000010000111100" => rgb <= "000000";
					when "00000010000111101" => rgb <= "000000";
					when "00000010000111110" => rgb <= "000000";
					when "00000010000111111" => rgb <= "000000";
					when "00000010001000000" => rgb <= "000000";
					when "00000010001000001" => rgb <= "000000";
					when "00000010001000010" => rgb <= "000000";
					when "00000010001000011" => rgb <= "000000";
					when "00000010001000100" => rgb <= "000000";
					when "00000010001000101" => rgb <= "000000";
					when "00000010001000110" => rgb <= "000000";
					when "00000010001000111" => rgb <= "000000";
					when "00000010001001000" => rgb <= "000000";
					when "00000010001001001" => rgb <= "000000";
					when "00000010001001010" => rgb <= "000000";
					when "00000010001001011" => rgb <= "000000";
					when "00000010001001100" => rgb <= "000000";
					when "00000010001001101" => rgb <= "000000";
					when "00000010001001110" => rgb <= "000000";
					when "00000010001001111" => rgb <= "000000";
					when "00000010001010000" => rgb <= "000000";
					when "00000010001010001" => rgb <= "000000";
					when "00000010001010010" => rgb <= "000000";
					when "00000010001010011" => rgb <= "000000";
					when "00000010001010100" => rgb <= "000000";
					when "00000010001010101" => rgb <= "000000";
					when "00000010001010110" => rgb <= "000000";
					when "00000010001010111" => rgb <= "000000";
					when "00000010001011000" => rgb <= "000000";
					when "00000010001011001" => rgb <= "000000";
					when "00000010001011010" => rgb <= "000000";
					when "00000010001011011" => rgb <= "000000";
					when "00000010001011100" => rgb <= "000000";
					when "00000010001011101" => rgb <= "000000";
					when "00000010001011110" => rgb <= "000000";
					when "00000010001011111" => rgb <= "000000";
					when "00000010001100000" => rgb <= "000000";
					when "00000010001100001" => rgb <= "000000";
					when "00000010001100010" => rgb <= "000000";
					when "00000010001100011" => rgb <= "000000";
					when "00000010001100100" => rgb <= "000000";
					when "00000010001100101" => rgb <= "000000";
					when "00000010001100110" => rgb <= "000000";
					when "00000010001100111" => rgb <= "000000";
					when "00000010001101000" => rgb <= "000000";
					when "00000010001101001" => rgb <= "000000";
					when "00000010001101010" => rgb <= "000000";
					when "00000010001101011" => rgb <= "000000";
					when "00000010001101100" => rgb <= "000000";
					when "00000010001101101" => rgb <= "000000";
					when "00000010001101110" => rgb <= "000000";
					when "00000010001101111" => rgb <= "000000";
					when "00000010001110000" => rgb <= "000000";
					when "00000010001110001" => rgb <= "000000";
					when "00000010001110010" => rgb <= "000000";
					when "00000010001110011" => rgb <= "000000";
					when "00000010001110100" => rgb <= "000000";
					when "00000010001110101" => rgb <= "000000";
					when "00000010001110110" => rgb <= "000000";
					when "00000010001110111" => rgb <= "000000";
					when "00000010001111000" => rgb <= "000000";
					when "00000010001111001" => rgb <= "000000";
					when "00000010001111010" => rgb <= "000000";
					when "00000010001111011" => rgb <= "000000";
					when "00000010001111100" => rgb <= "000000";
					when "00000010001111101" => rgb <= "000000";
					when "00000010001111110" => rgb <= "000000";
					when "00000010001111111" => rgb <= "000000";
					when "00000010010000000" => rgb <= "000000";
					when "00000010010000001" => rgb <= "000000";
					when "00000010010000010" => rgb <= "000000";
					when "00000010010000011" => rgb <= "000000";
					when "00000010010000100" => rgb <= "000000";
					when "00000010010000101" => rgb <= "000000";
					when "00000010010000110" => rgb <= "000000";
					when "00000010010000111" => rgb <= "000000";
					when "00000010010001000" => rgb <= "000000";
					when "00000010010001001" => rgb <= "000000";
					when "00000010010001010" => rgb <= "000000";
					when "00000010010001011" => rgb <= "000000";
					when "00000010010001100" => rgb <= "000000";
					when "00000010010001101" => rgb <= "000000";
					when "00000010010001110" => rgb <= "000000";
					when "00000010010001111" => rgb <= "000000";
					when "00000010010010000" => rgb <= "000000";
					when "00000010010010001" => rgb <= "000000";
					when "00000010010010010" => rgb <= "000000";
					when "00000010010010011" => rgb <= "000000";
					when "00000010010010100" => rgb <= "000000";
					when "00000010010010101" => rgb <= "000000";
					when "00000010010010110" => rgb <= "000000";
					when "00000010010010111" => rgb <= "000000";
					when "00000010010011000" => rgb <= "000000";
					when "00000010010011001" => rgb <= "000000";
					when "00000010010011010" => rgb <= "000000";
					when "00000010010011011" => rgb <= "000000";
					when "00000010010011100" => rgb <= "000000";
					when "00000010010011101" => rgb <= "000000";
					when "00000010010011110" => rgb <= "000000";
					when "00000010010011111" => rgb <= "000000";
					when "00000010010100000" => rgb <= "000000";
					when "00000010010100001" => rgb <= "000000";
					when "00000010010100010" => rgb <= "000000";
					when "00000010010100011" => rgb <= "000000";
					when "00000010010100100" => rgb <= "000000";
					when "00000010010100101" => rgb <= "000000";
					when "00000010010100110" => rgb <= "000000";
					when "00000010010100111" => rgb <= "000000";
					when "00000010010101000" => rgb <= "000000";
					when "00000010010101001" => rgb <= "000000";
					when "00000010010101010" => rgb <= "000000";
					when "00000010010101011" => rgb <= "000000";
					when "00000010010101100" => rgb <= "000000";
					when "00000010010101101" => rgb <= "000000";
					when "00000010010101110" => rgb <= "000000";
					when "00000010010101111" => rgb <= "000000";
					when "00000010010110000" => rgb <= "000000";
					when "00000010010110001" => rgb <= "000000";
					when "00000010010110010" => rgb <= "000000";
					when "00000010010110011" => rgb <= "000000";
					when "00000010010110100" => rgb <= "000000";
					when "00000010010110101" => rgb <= "000000";
					when "00000010010110110" => rgb <= "000000";
					when "00000010010110111" => rgb <= "000000";
					when "00000010010111000" => rgb <= "000000";
					when "00000010010111001" => rgb <= "000000";
					when "00000010010111010" => rgb <= "000000";
					when "00000010010111011" => rgb <= "000000";
					when "00000010010111100" => rgb <= "000000";
					when "00000010010111101" => rgb <= "000000";
					when "00000010010111110" => rgb <= "000000";
					when "00000010010111111" => rgb <= "000000";
					when "00000010011000000" => rgb <= "000000";
					when "00000010011000001" => rgb <= "000000";
					when "00000010011000010" => rgb <= "000000";
					when "00000010011000011" => rgb <= "000000";
					when "00000010011000100" => rgb <= "000000";
					when "00000010011000101" => rgb <= "000000";
					when "00000010011000110" => rgb <= "000000";
					when "00000010011000111" => rgb <= "000000";
					when "00000010011001000" => rgb <= "000000";
					when "00000010011001001" => rgb <= "000000";
					when "00000010011001010" => rgb <= "000000";
					when "00000010011001011" => rgb <= "000000";
					when "00000010011001100" => rgb <= "000000";
					when "00000010011001101" => rgb <= "000000";
					when "00000010011001110" => rgb <= "000000";
					when "00000010011001111" => rgb <= "000000";
					when "00000010011010000" => rgb <= "000000";
					when "00000010011010001" => rgb <= "000000";
					when "00000010011010010" => rgb <= "000000";
					when "00000010011010011" => rgb <= "000000";
					when "00000010011010100" => rgb <= "000000";
					when "00000010011010101" => rgb <= "000000";
					when "00000010011010110" => rgb <= "000000";
					when "00000010011010111" => rgb <= "000000";
					when "00000010011011000" => rgb <= "000000";
					when "00000010011011001" => rgb <= "000000";
					when "00000010011011010" => rgb <= "000000";
					when "00000010011011011" => rgb <= "000000";
					when "00000010011011100" => rgb <= "000000";
					when "00000010011011101" => rgb <= "000000";
					when "00000010011011110" => rgb <= "000000";
					when "00000010011011111" => rgb <= "000000";
					when "00000010011100000" => rgb <= "000000";
					when "00000010011100001" => rgb <= "000000";
					when "00000010011100010" => rgb <= "000000";
					when "00000010011100011" => rgb <= "000000";
					when "00000010011100100" => rgb <= "000000";
					when "00000010011100101" => rgb <= "000000";
					when "00000010011100110" => rgb <= "000000";
					when "00000010011100111" => rgb <= "000000";
					when "00000010011101000" => rgb <= "000000";
					when "00000010011101001" => rgb <= "000000";
					when "00000010011101010" => rgb <= "000000";
					when "00000010011101011" => rgb <= "000000";
					when "00000010011101100" => rgb <= "000000";
					when "00000010011101101" => rgb <= "000000";
					when "00000010011101110" => rgb <= "000000";
					when "00000010011101111" => rgb <= "000000";
					when "00000010011110000" => rgb <= "000000";
					when "00000010011110001" => rgb <= "000000";
					when "00000010011110010" => rgb <= "000000";
					when "00000010011110011" => rgb <= "000000";
					when "00000010011110100" => rgb <= "000000";
					when "00000010011110101" => rgb <= "000000";
					when "00000010011110110" => rgb <= "000000";
					when "00000010011110111" => rgb <= "000000";
					when "00000010011111000" => rgb <= "000000";
					when "00000010011111001" => rgb <= "000000";
					when "00000010011111010" => rgb <= "000000";
					when "00000010011111011" => rgb <= "000000";
					when "00000010011111100" => rgb <= "000000";
					when "00000010011111101" => rgb <= "000000";
					when "00000010011111110" => rgb <= "000000";
					when "00000010011111111" => rgb <= "000000";
					when "00000010100000000" => rgb <= "000000";
					when "00000010100000001" => rgb <= "000000";
					when "00000010100000010" => rgb <= "000000";
					when "00000010100000011" => rgb <= "000000";
					when "00000010100000100" => rgb <= "000000";
					when "00000010100000101" => rgb <= "000000";
					when "00000010100000110" => rgb <= "000000";
					when "00000010100000111" => rgb <= "000000";
					when "00000010100001000" => rgb <= "000000";
					when "00000010100001001" => rgb <= "000000";
					when "00000010100001010" => rgb <= "000000";
					when "00000010100001011" => rgb <= "000000";
					when "00000010100001100" => rgb <= "000000";
					when "00000010100001101" => rgb <= "000000";
					when "00000010100001110" => rgb <= "000000";
					when "00000010100001111" => rgb <= "000000";
					when "00000010100010000" => rgb <= "000000";
					when "00000010100010001" => rgb <= "000000";
					when "00000010100010010" => rgb <= "000000";
					when "00000010100010011" => rgb <= "000000";
					when "00000010100010100" => rgb <= "000000";
					when "00000010100010101" => rgb <= "000000";
					when "00000010100010110" => rgb <= "000000";
					when "00000010100010111" => rgb <= "000000";
					when "00000010100011000" => rgb <= "000000";
					when "00000010100011001" => rgb <= "000000";
					when "00000010100011010" => rgb <= "000000";
					when "00000010100011011" => rgb <= "000000";
					when "00000010100011100" => rgb <= "000000";
					when "00000010100011101" => rgb <= "000000";
					when "00000010100011110" => rgb <= "000000";
					when "00000010100011111" => rgb <= "000000";
					when "00000010100100000" => rgb <= "000000";
					when "00000010100100001" => rgb <= "000000";
					when "00000010100100010" => rgb <= "000000";
					when "00000010100100011" => rgb <= "000000";
					when "00000010100100100" => rgb <= "000000";
					when "00000010100100101" => rgb <= "000000";
					when "00000010100100110" => rgb <= "000000";
					when "00000010100100111" => rgb <= "000000";
					when "00000010100101000" => rgb <= "000000";
					when "00000010100101001" => rgb <= "000000";
					when "00000010100101010" => rgb <= "000000";
					when "00000010100101011" => rgb <= "000000";
					when "00000010100101100" => rgb <= "000000";
					when "00000010100101101" => rgb <= "000000";
					when "00000010100101110" => rgb <= "000000";
					when "00000010100101111" => rgb <= "000000";
					when "00000010100110000" => rgb <= "000000";
					when "00000010100110001" => rgb <= "000000";
					when "00000010100110010" => rgb <= "000000";
					when "00000010100110011" => rgb <= "000000";
					when "00000010100110100" => rgb <= "000000";
					when "00000010100110101" => rgb <= "000000";
					when "00000010100110110" => rgb <= "000000";
					when "00000010100110111" => rgb <= "000000";
					when "00000010100111000" => rgb <= "000000";
					when "00000010100111001" => rgb <= "000000";
					when "00000010100111010" => rgb <= "000000";
					when "00000010100111011" => rgb <= "000000";
					when "00000010100111100" => rgb <= "000000";
					when "00000010100111101" => rgb <= "000000";
					when "00000010100111110" => rgb <= "000000";
					when "00000010100111111" => rgb <= "000000";
					when "00000011000000000" => rgb <= "000000";
					when "00000011000000001" => rgb <= "000000";
					when "00000011000000010" => rgb <= "000000";
					when "00000011000000011" => rgb <= "000000";
					when "00000011000000100" => rgb <= "000000";
					when "00000011000000101" => rgb <= "000000";
					when "00000011000000110" => rgb <= "000000";
					when "00000011000000111" => rgb <= "000000";
					when "00000011000001000" => rgb <= "000000";
					when "00000011000001001" => rgb <= "000000";
					when "00000011000001010" => rgb <= "000000";
					when "00000011000001011" => rgb <= "000000";
					when "00000011000001100" => rgb <= "000000";
					when "00000011000001101" => rgb <= "000000";
					when "00000011000001110" => rgb <= "000000";
					when "00000011000001111" => rgb <= "000000";
					when "00000011000010000" => rgb <= "000000";
					when "00000011000010001" => rgb <= "000000";
					when "00000011000010010" => rgb <= "000000";
					when "00000011000010011" => rgb <= "000000";
					when "00000011000010100" => rgb <= "000000";
					when "00000011000010101" => rgb <= "000000";
					when "00000011000010110" => rgb <= "000000";
					when "00000011000010111" => rgb <= "000000";
					when "00000011000011000" => rgb <= "000000";
					when "00000011000011001" => rgb <= "000000";
					when "00000011000011010" => rgb <= "000000";
					when "00000011000011011" => rgb <= "000000";
					when "00000011000011100" => rgb <= "000000";
					when "00000011000011101" => rgb <= "000000";
					when "00000011000011110" => rgb <= "000000";
					when "00000011000011111" => rgb <= "000000";
					when "00000011000100000" => rgb <= "000000";
					when "00000011000100001" => rgb <= "000000";
					when "00000011000100010" => rgb <= "000000";
					when "00000011000100011" => rgb <= "000000";
					when "00000011000100100" => rgb <= "000000";
					when "00000011000100101" => rgb <= "000000";
					when "00000011000100110" => rgb <= "000000";
					when "00000011000100111" => rgb <= "000000";
					when "00000011000101000" => rgb <= "000000";
					when "00000011000101001" => rgb <= "000000";
					when "00000011000101010" => rgb <= "000000";
					when "00000011000101011" => rgb <= "000000";
					when "00000011000101100" => rgb <= "000000";
					when "00000011000101101" => rgb <= "000000";
					when "00000011000101110" => rgb <= "000000";
					when "00000011000101111" => rgb <= "000000";
					when "00000011000110000" => rgb <= "000000";
					when "00000011000110001" => rgb <= "000000";
					when "00000011000110010" => rgb <= "000000";
					when "00000011000110011" => rgb <= "000000";
					when "00000011000110100" => rgb <= "000000";
					when "00000011000110101" => rgb <= "000000";
					when "00000011000110110" => rgb <= "000000";
					when "00000011000110111" => rgb <= "000000";
					when "00000011000111000" => rgb <= "000000";
					when "00000011000111001" => rgb <= "000000";
					when "00000011000111010" => rgb <= "000000";
					when "00000011000111011" => rgb <= "000000";
					when "00000011000111100" => rgb <= "000000";
					when "00000011000111101" => rgb <= "000000";
					when "00000011000111110" => rgb <= "000000";
					when "00000011000111111" => rgb <= "000000";
					when "00000011001000000" => rgb <= "000000";
					when "00000011001000001" => rgb <= "000000";
					when "00000011001000010" => rgb <= "000000";
					when "00000011001000011" => rgb <= "000000";
					when "00000011001000100" => rgb <= "000000";
					when "00000011001000101" => rgb <= "000000";
					when "00000011001000110" => rgb <= "000000";
					when "00000011001000111" => rgb <= "000000";
					when "00000011001001000" => rgb <= "000000";
					when "00000011001001001" => rgb <= "000000";
					when "00000011001001010" => rgb <= "000000";
					when "00000011001001011" => rgb <= "000000";
					when "00000011001001100" => rgb <= "000000";
					when "00000011001001101" => rgb <= "000000";
					when "00000011001001110" => rgb <= "000000";
					when "00000011001001111" => rgb <= "000000";
					when "00000011001010000" => rgb <= "000000";
					when "00000011001010001" => rgb <= "000000";
					when "00000011001010010" => rgb <= "000000";
					when "00000011001010011" => rgb <= "000000";
					when "00000011001010100" => rgb <= "000000";
					when "00000011001010101" => rgb <= "000000";
					when "00000011001010110" => rgb <= "000000";
					when "00000011001010111" => rgb <= "000000";
					when "00000011001011000" => rgb <= "000000";
					when "00000011001011001" => rgb <= "000000";
					when "00000011001011010" => rgb <= "000000";
					when "00000011001011011" => rgb <= "000000";
					when "00000011001011100" => rgb <= "000000";
					when "00000011001011101" => rgb <= "000000";
					when "00000011001011110" => rgb <= "000000";
					when "00000011001011111" => rgb <= "000000";
					when "00000011001100000" => rgb <= "000000";
					when "00000011001100001" => rgb <= "000000";
					when "00000011001100010" => rgb <= "000000";
					when "00000011001100011" => rgb <= "000000";
					when "00000011001100100" => rgb <= "000000";
					when "00000011001100101" => rgb <= "000000";
					when "00000011001100110" => rgb <= "000000";
					when "00000011001100111" => rgb <= "000000";
					when "00000011001101000" => rgb <= "000000";
					when "00000011001101001" => rgb <= "000000";
					when "00000011001101010" => rgb <= "000000";
					when "00000011001101011" => rgb <= "000000";
					when "00000011001101100" => rgb <= "000000";
					when "00000011001101101" => rgb <= "000000";
					when "00000011001101110" => rgb <= "000000";
					when "00000011001101111" => rgb <= "000000";
					when "00000011001110000" => rgb <= "000000";
					when "00000011001110001" => rgb <= "000000";
					when "00000011001110010" => rgb <= "000000";
					when "00000011001110011" => rgb <= "000000";
					when "00000011001110100" => rgb <= "000000";
					when "00000011001110101" => rgb <= "000000";
					when "00000011001110110" => rgb <= "000000";
					when "00000011001110111" => rgb <= "000000";
					when "00000011001111000" => rgb <= "000000";
					when "00000011001111001" => rgb <= "000000";
					when "00000011001111010" => rgb <= "000000";
					when "00000011001111011" => rgb <= "000000";
					when "00000011001111100" => rgb <= "000000";
					when "00000011001111101" => rgb <= "000000";
					when "00000011001111110" => rgb <= "000000";
					when "00000011001111111" => rgb <= "000000";
					when "00000011010000000" => rgb <= "000000";
					when "00000011010000001" => rgb <= "000000";
					when "00000011010000010" => rgb <= "000000";
					when "00000011010000011" => rgb <= "000000";
					when "00000011010000100" => rgb <= "000000";
					when "00000011010000101" => rgb <= "000000";
					when "00000011010000110" => rgb <= "000000";
					when "00000011010000111" => rgb <= "000000";
					when "00000011010001000" => rgb <= "000000";
					when "00000011010001001" => rgb <= "000000";
					when "00000011010001010" => rgb <= "000000";
					when "00000011010001011" => rgb <= "000000";
					when "00000011010001100" => rgb <= "000000";
					when "00000011010001101" => rgb <= "000000";
					when "00000011010001110" => rgb <= "000000";
					when "00000011010001111" => rgb <= "000000";
					when "00000011010010000" => rgb <= "000000";
					when "00000011010010001" => rgb <= "000000";
					when "00000011010010010" => rgb <= "000000";
					when "00000011010010011" => rgb <= "000000";
					when "00000011010010100" => rgb <= "000000";
					when "00000011010010101" => rgb <= "000000";
					when "00000011010010110" => rgb <= "000000";
					when "00000011010010111" => rgb <= "000000";
					when "00000011010011000" => rgb <= "000000";
					when "00000011010011001" => rgb <= "000000";
					when "00000011010011010" => rgb <= "000000";
					when "00000011010011011" => rgb <= "000000";
					when "00000011010011100" => rgb <= "000000";
					when "00000011010011101" => rgb <= "000000";
					when "00000011010011110" => rgb <= "000000";
					when "00000011010011111" => rgb <= "000000";
					when "00000011010100000" => rgb <= "000000";
					when "00000011010100001" => rgb <= "000000";
					when "00000011010100010" => rgb <= "000000";
					when "00000011010100011" => rgb <= "000000";
					when "00000011010100100" => rgb <= "000000";
					when "00000011010100101" => rgb <= "000000";
					when "00000011010100110" => rgb <= "000000";
					when "00000011010100111" => rgb <= "000000";
					when "00000011010101000" => rgb <= "000000";
					when "00000011010101001" => rgb <= "000000";
					when "00000011010101010" => rgb <= "000000";
					when "00000011010101011" => rgb <= "000000";
					when "00000011010101100" => rgb <= "000000";
					when "00000011010101101" => rgb <= "000000";
					when "00000011010101110" => rgb <= "000000";
					when "00000011010101111" => rgb <= "000000";
					when "00000011010110000" => rgb <= "000000";
					when "00000011010110001" => rgb <= "000000";
					when "00000011010110010" => rgb <= "000000";
					when "00000011010110011" => rgb <= "000000";
					when "00000011010110100" => rgb <= "000000";
					when "00000011010110101" => rgb <= "000000";
					when "00000011010110110" => rgb <= "000000";
					when "00000011010110111" => rgb <= "000000";
					when "00000011010111000" => rgb <= "000000";
					when "00000011010111001" => rgb <= "000000";
					when "00000011010111010" => rgb <= "000000";
					when "00000011010111011" => rgb <= "000000";
					when "00000011010111100" => rgb <= "000000";
					when "00000011010111101" => rgb <= "000000";
					when "00000011010111110" => rgb <= "000000";
					when "00000011010111111" => rgb <= "000000";
					when "00000011011000000" => rgb <= "000000";
					when "00000011011000001" => rgb <= "000000";
					when "00000011011000010" => rgb <= "000000";
					when "00000011011000011" => rgb <= "000000";
					when "00000011011000100" => rgb <= "000000";
					when "00000011011000101" => rgb <= "000000";
					when "00000011011000110" => rgb <= "000000";
					when "00000011011000111" => rgb <= "000000";
					when "00000011011001000" => rgb <= "000000";
					when "00000011011001001" => rgb <= "000000";
					when "00000011011001010" => rgb <= "000000";
					when "00000011011001011" => rgb <= "000000";
					when "00000011011001100" => rgb <= "000000";
					when "00000011011001101" => rgb <= "000000";
					when "00000011011001110" => rgb <= "000000";
					when "00000011011001111" => rgb <= "000000";
					when "00000011011010000" => rgb <= "000000";
					when "00000011011010001" => rgb <= "000000";
					when "00000011011010010" => rgb <= "000000";
					when "00000011011010011" => rgb <= "000000";
					when "00000011011010100" => rgb <= "000000";
					when "00000011011010101" => rgb <= "000000";
					when "00000011011010110" => rgb <= "000000";
					when "00000011011010111" => rgb <= "000000";
					when "00000011011011000" => rgb <= "000000";
					when "00000011011011001" => rgb <= "000000";
					when "00000011011011010" => rgb <= "000000";
					when "00000011011011011" => rgb <= "000000";
					when "00000011011011100" => rgb <= "000000";
					when "00000011011011101" => rgb <= "000000";
					when "00000011011011110" => rgb <= "000000";
					when "00000011011011111" => rgb <= "000000";
					when "00000011011100000" => rgb <= "000000";
					when "00000011011100001" => rgb <= "000000";
					when "00000011011100010" => rgb <= "000000";
					when "00000011011100011" => rgb <= "000000";
					when "00000011011100100" => rgb <= "000000";
					when "00000011011100101" => rgb <= "000000";
					when "00000011011100110" => rgb <= "000000";
					when "00000011011100111" => rgb <= "000000";
					when "00000011011101000" => rgb <= "000000";
					when "00000011011101001" => rgb <= "000000";
					when "00000011011101010" => rgb <= "000000";
					when "00000011011101011" => rgb <= "000000";
					when "00000011011101100" => rgb <= "000000";
					when "00000011011101101" => rgb <= "000000";
					when "00000011011101110" => rgb <= "000000";
					when "00000011011101111" => rgb <= "000000";
					when "00000011011110000" => rgb <= "000000";
					when "00000011011110001" => rgb <= "000000";
					when "00000011011110010" => rgb <= "000000";
					when "00000011011110011" => rgb <= "000000";
					when "00000011011110100" => rgb <= "000000";
					when "00000011011110101" => rgb <= "000000";
					when "00000011011110110" => rgb <= "000000";
					when "00000011011110111" => rgb <= "000000";
					when "00000011011111000" => rgb <= "000000";
					when "00000011011111001" => rgb <= "000000";
					when "00000011011111010" => rgb <= "000000";
					when "00000011011111011" => rgb <= "000000";
					when "00000011011111100" => rgb <= "000000";
					when "00000011011111101" => rgb <= "000000";
					when "00000011011111110" => rgb <= "000000";
					when "00000011011111111" => rgb <= "000000";
					when "00000011100000000" => rgb <= "000000";
					when "00000011100000001" => rgb <= "000000";
					when "00000011100000010" => rgb <= "000000";
					when "00000011100000011" => rgb <= "000000";
					when "00000011100000100" => rgb <= "000000";
					when "00000011100000101" => rgb <= "000000";
					when "00000011100000110" => rgb <= "000000";
					when "00000011100000111" => rgb <= "000000";
					when "00000011100001000" => rgb <= "000000";
					when "00000011100001001" => rgb <= "000000";
					when "00000011100001010" => rgb <= "000000";
					when "00000011100001011" => rgb <= "000000";
					when "00000011100001100" => rgb <= "000000";
					when "00000011100001101" => rgb <= "000000";
					when "00000011100001110" => rgb <= "000000";
					when "00000011100001111" => rgb <= "000000";
					when "00000011100010000" => rgb <= "000000";
					when "00000011100010001" => rgb <= "000000";
					when "00000011100010010" => rgb <= "000000";
					when "00000011100010011" => rgb <= "000000";
					when "00000011100010100" => rgb <= "000000";
					when "00000011100010101" => rgb <= "000000";
					when "00000011100010110" => rgb <= "000000";
					when "00000011100010111" => rgb <= "000000";
					when "00000011100011000" => rgb <= "000000";
					when "00000011100011001" => rgb <= "000000";
					when "00000011100011010" => rgb <= "000000";
					when "00000011100011011" => rgb <= "000000";
					when "00000011100011100" => rgb <= "000000";
					when "00000011100011101" => rgb <= "000000";
					when "00000011100011110" => rgb <= "000000";
					when "00000011100011111" => rgb <= "000000";
					when "00000011100100000" => rgb <= "000000";
					when "00000011100100001" => rgb <= "000000";
					when "00000011100100010" => rgb <= "000000";
					when "00000011100100011" => rgb <= "000000";
					when "00000011100100100" => rgb <= "000000";
					when "00000011100100101" => rgb <= "000000";
					when "00000011100100110" => rgb <= "000000";
					when "00000011100100111" => rgb <= "000000";
					when "00000011100101000" => rgb <= "000000";
					when "00000011100101001" => rgb <= "000000";
					when "00000011100101010" => rgb <= "000000";
					when "00000011100101011" => rgb <= "000000";
					when "00000011100101100" => rgb <= "000000";
					when "00000011100101101" => rgb <= "000000";
					when "00000011100101110" => rgb <= "000000";
					when "00000011100101111" => rgb <= "000000";
					when "00000011100110000" => rgb <= "000000";
					when "00000011100110001" => rgb <= "000000";
					when "00000011100110010" => rgb <= "000000";
					when "00000011100110011" => rgb <= "000000";
					when "00000011100110100" => rgb <= "000000";
					when "00000011100110101" => rgb <= "000000";
					when "00000011100110110" => rgb <= "000000";
					when "00000011100110111" => rgb <= "000000";
					when "00000011100111000" => rgb <= "000000";
					when "00000011100111001" => rgb <= "000000";
					when "00000011100111010" => rgb <= "000000";
					when "00000011100111011" => rgb <= "000000";
					when "00000011100111100" => rgb <= "000000";
					when "00000011100111101" => rgb <= "000000";
					when "00000011100111110" => rgb <= "000000";
					when "00000011100111111" => rgb <= "000000";
					when "00000100000000000" => rgb <= "000000";
					when "00000100000000001" => rgb <= "000000";
					when "00000100000000010" => rgb <= "000000";
					when "00000100000000011" => rgb <= "000000";
					when "00000100000000100" => rgb <= "000000";
					when "00000100000000101" => rgb <= "000000";
					when "00000100000000110" => rgb <= "000000";
					when "00000100000000111" => rgb <= "000000";
					when "00000100000001000" => rgb <= "000000";
					when "00000100000001001" => rgb <= "000000";
					when "00000100000001010" => rgb <= "000000";
					when "00000100000001011" => rgb <= "000000";
					when "00000100000001100" => rgb <= "000000";
					when "00000100000001101" => rgb <= "000000";
					when "00000100000001110" => rgb <= "000000";
					when "00000100000001111" => rgb <= "000000";
					when "00000100000010000" => rgb <= "000000";
					when "00000100000010001" => rgb <= "000000";
					when "00000100000010010" => rgb <= "000000";
					when "00000100000010011" => rgb <= "000000";
					when "00000100000010100" => rgb <= "000000";
					when "00000100000010101" => rgb <= "000000";
					when "00000100000010110" => rgb <= "000000";
					when "00000100000010111" => rgb <= "000000";
					when "00000100000011000" => rgb <= "000000";
					when "00000100000011001" => rgb <= "000000";
					when "00000100000011010" => rgb <= "000000";
					when "00000100000011011" => rgb <= "000000";
					when "00000100000011100" => rgb <= "000000";
					when "00000100000011101" => rgb <= "000000";
					when "00000100000011110" => rgb <= "000000";
					when "00000100000011111" => rgb <= "000000";
					when "00000100000100000" => rgb <= "000000";
					when "00000100000100001" => rgb <= "000000";
					when "00000100000100010" => rgb <= "000000";
					when "00000100000100011" => rgb <= "000000";
					when "00000100000100100" => rgb <= "000000";
					when "00000100000100101" => rgb <= "000000";
					when "00000100000100110" => rgb <= "000000";
					when "00000100000100111" => rgb <= "000000";
					when "00000100000101000" => rgb <= "000000";
					when "00000100000101001" => rgb <= "000000";
					when "00000100000101010" => rgb <= "000000";
					when "00000100000101011" => rgb <= "000000";
					when "00000100000101100" => rgb <= "000000";
					when "00000100000101101" => rgb <= "000000";
					when "00000100000101110" => rgb <= "000000";
					when "00000100000101111" => rgb <= "000000";
					when "00000100000110000" => rgb <= "000000";
					when "00000100000110001" => rgb <= "000000";
					when "00000100000110010" => rgb <= "000000";
					when "00000100000110011" => rgb <= "000000";
					when "00000100000110100" => rgb <= "000000";
					when "00000100000110101" => rgb <= "000000";
					when "00000100000110110" => rgb <= "000000";
					when "00000100000110111" => rgb <= "000000";
					when "00000100000111000" => rgb <= "000000";
					when "00000100000111001" => rgb <= "000000";
					when "00000100000111010" => rgb <= "000000";
					when "00000100000111011" => rgb <= "000000";
					when "00000100000111100" => rgb <= "000000";
					when "00000100000111101" => rgb <= "000000";
					when "00000100000111110" => rgb <= "000000";
					when "00000100000111111" => rgb <= "000000";
					when "00000100001000000" => rgb <= "000000";
					when "00000100001000001" => rgb <= "000000";
					when "00000100001000010" => rgb <= "000000";
					when "00000100001000011" => rgb <= "000000";
					when "00000100001000100" => rgb <= "000000";
					when "00000100001000101" => rgb <= "000000";
					when "00000100001000110" => rgb <= "000000";
					when "00000100001000111" => rgb <= "000000";
					when "00000100001001000" => rgb <= "000000";
					when "00000100001001001" => rgb <= "000000";
					when "00000100001001010" => rgb <= "000000";
					when "00000100001001011" => rgb <= "000000";
					when "00000100001001100" => rgb <= "000000";
					when "00000100001001101" => rgb <= "000000";
					when "00000100001001110" => rgb <= "000000";
					when "00000100001001111" => rgb <= "000000";
					when "00000100001010000" => rgb <= "000000";
					when "00000100001010001" => rgb <= "000000";
					when "00000100001010010" => rgb <= "000000";
					when "00000100001010011" => rgb <= "000000";
					when "00000100001010100" => rgb <= "000000";
					when "00000100001010101" => rgb <= "000000";
					when "00000100001010110" => rgb <= "000000";
					when "00000100001010111" => rgb <= "000000";
					when "00000100001011000" => rgb <= "000000";
					when "00000100001011001" => rgb <= "000000";
					when "00000100001011010" => rgb <= "000000";
					when "00000100001011011" => rgb <= "000000";
					when "00000100001011100" => rgb <= "000000";
					when "00000100001011101" => rgb <= "000000";
					when "00000100001011110" => rgb <= "000000";
					when "00000100001011111" => rgb <= "000000";
					when "00000100001100000" => rgb <= "000000";
					when "00000100001100001" => rgb <= "000000";
					when "00000100001100010" => rgb <= "000000";
					when "00000100001100011" => rgb <= "000000";
					when "00000100001100100" => rgb <= "000000";
					when "00000100001100101" => rgb <= "000000";
					when "00000100001100110" => rgb <= "000000";
					when "00000100001100111" => rgb <= "000000";
					when "00000100001101000" => rgb <= "000000";
					when "00000100001101001" => rgb <= "000000";
					when "00000100001101010" => rgb <= "000000";
					when "00000100001101011" => rgb <= "000000";
					when "00000100001101100" => rgb <= "000000";
					when "00000100001101101" => rgb <= "000000";
					when "00000100001101110" => rgb <= "000000";
					when "00000100001101111" => rgb <= "000000";
					when "00000100001110000" => rgb <= "000000";
					when "00000100001110001" => rgb <= "000000";
					when "00000100001110010" => rgb <= "000000";
					when "00000100001110011" => rgb <= "000000";
					when "00000100001110100" => rgb <= "000000";
					when "00000100001110101" => rgb <= "000000";
					when "00000100001110110" => rgb <= "000000";
					when "00000100001110111" => rgb <= "000000";
					when "00000100001111000" => rgb <= "000000";
					when "00000100001111001" => rgb <= "000000";
					when "00000100001111010" => rgb <= "000000";
					when "00000100001111011" => rgb <= "000000";
					when "00000100001111100" => rgb <= "000000";
					when "00000100001111101" => rgb <= "000000";
					when "00000100001111110" => rgb <= "000000";
					when "00000100001111111" => rgb <= "000000";
					when "00000100010000000" => rgb <= "000000";
					when "00000100010000001" => rgb <= "000000";
					when "00000100010000010" => rgb <= "000000";
					when "00000100010000011" => rgb <= "000000";
					when "00000100010000100" => rgb <= "000000";
					when "00000100010000101" => rgb <= "000000";
					when "00000100010000110" => rgb <= "000000";
					when "00000100010000111" => rgb <= "000000";
					when "00000100010001000" => rgb <= "000000";
					when "00000100010001001" => rgb <= "000000";
					when "00000100010001010" => rgb <= "000000";
					when "00000100010001011" => rgb <= "000000";
					when "00000100010001100" => rgb <= "000000";
					when "00000100010001101" => rgb <= "000000";
					when "00000100010001110" => rgb <= "000000";
					when "00000100010001111" => rgb <= "000000";
					when "00000100010010000" => rgb <= "000000";
					when "00000100010010001" => rgb <= "000000";
					when "00000100010010010" => rgb <= "000000";
					when "00000100010010011" => rgb <= "000000";
					when "00000100010010100" => rgb <= "000000";
					when "00000100010010101" => rgb <= "000000";
					when "00000100010010110" => rgb <= "000000";
					when "00000100010010111" => rgb <= "000000";
					when "00000100010011000" => rgb <= "000000";
					when "00000100010011001" => rgb <= "000000";
					when "00000100010011010" => rgb <= "000000";
					when "00000100010011011" => rgb <= "000000";
					when "00000100010011100" => rgb <= "000000";
					when "00000100010011101" => rgb <= "000000";
					when "00000100010011110" => rgb <= "000000";
					when "00000100010011111" => rgb <= "000000";
					when "00000100010100000" => rgb <= "000000";
					when "00000100010100001" => rgb <= "000000";
					when "00000100010100010" => rgb <= "000000";
					when "00000100010100011" => rgb <= "000000";
					when "00000100010100100" => rgb <= "000000";
					when "00000100010100101" => rgb <= "000000";
					when "00000100010100110" => rgb <= "000000";
					when "00000100010100111" => rgb <= "000000";
					when "00000100010101000" => rgb <= "000000";
					when "00000100010101001" => rgb <= "000000";
					when "00000100010101010" => rgb <= "000000";
					when "00000100010101011" => rgb <= "000000";
					when "00000100010101100" => rgb <= "000000";
					when "00000100010101101" => rgb <= "000000";
					when "00000100010101110" => rgb <= "000000";
					when "00000100010101111" => rgb <= "000000";
					when "00000100010110000" => rgb <= "000000";
					when "00000100010110001" => rgb <= "000000";
					when "00000100010110010" => rgb <= "000000";
					when "00000100010110011" => rgb <= "000000";
					when "00000100010110100" => rgb <= "000000";
					when "00000100010110101" => rgb <= "000000";
					when "00000100010110110" => rgb <= "000000";
					when "00000100010110111" => rgb <= "000000";
					when "00000100010111000" => rgb <= "000000";
					when "00000100010111001" => rgb <= "000000";
					when "00000100010111010" => rgb <= "000000";
					when "00000100010111011" => rgb <= "000000";
					when "00000100010111100" => rgb <= "000000";
					when "00000100010111101" => rgb <= "000000";
					when "00000100010111110" => rgb <= "000000";
					when "00000100010111111" => rgb <= "000000";
					when "00000100011000000" => rgb <= "000000";
					when "00000100011000001" => rgb <= "000000";
					when "00000100011000010" => rgb <= "000000";
					when "00000100011000011" => rgb <= "000000";
					when "00000100011000100" => rgb <= "000000";
					when "00000100011000101" => rgb <= "000000";
					when "00000100011000110" => rgb <= "000000";
					when "00000100011000111" => rgb <= "000000";
					when "00000100011001000" => rgb <= "000000";
					when "00000100011001001" => rgb <= "000000";
					when "00000100011001010" => rgb <= "000000";
					when "00000100011001011" => rgb <= "000000";
					when "00000100011001100" => rgb <= "000000";
					when "00000100011001101" => rgb <= "000000";
					when "00000100011001110" => rgb <= "000000";
					when "00000100011001111" => rgb <= "000000";
					when "00000100011010000" => rgb <= "000000";
					when "00000100011010001" => rgb <= "000000";
					when "00000100011010010" => rgb <= "000000";
					when "00000100011010011" => rgb <= "000000";
					when "00000100011010100" => rgb <= "000000";
					when "00000100011010101" => rgb <= "000000";
					when "00000100011010110" => rgb <= "000000";
					when "00000100011010111" => rgb <= "000000";
					when "00000100011011000" => rgb <= "000000";
					when "00000100011011001" => rgb <= "000000";
					when "00000100011011010" => rgb <= "000000";
					when "00000100011011011" => rgb <= "000000";
					when "00000100011011100" => rgb <= "000000";
					when "00000100011011101" => rgb <= "000000";
					when "00000100011011110" => rgb <= "000000";
					when "00000100011011111" => rgb <= "000000";
					when "00000100011100000" => rgb <= "000000";
					when "00000100011100001" => rgb <= "000000";
					when "00000100011100010" => rgb <= "000000";
					when "00000100011100011" => rgb <= "000000";
					when "00000100011100100" => rgb <= "000000";
					when "00000100011100101" => rgb <= "000000";
					when "00000100011100110" => rgb <= "000000";
					when "00000100011100111" => rgb <= "000000";
					when "00000100011101000" => rgb <= "000000";
					when "00000100011101001" => rgb <= "000000";
					when "00000100011101010" => rgb <= "000000";
					when "00000100011101011" => rgb <= "000000";
					when "00000100011101100" => rgb <= "000000";
					when "00000100011101101" => rgb <= "000000";
					when "00000100011101110" => rgb <= "000000";
					when "00000100011101111" => rgb <= "000000";
					when "00000100011110000" => rgb <= "000000";
					when "00000100011110001" => rgb <= "000000";
					when "00000100011110010" => rgb <= "000000";
					when "00000100011110011" => rgb <= "000000";
					when "00000100011110100" => rgb <= "000000";
					when "00000100011110101" => rgb <= "000000";
					when "00000100011110110" => rgb <= "000000";
					when "00000100011110111" => rgb <= "000000";
					when "00000100011111000" => rgb <= "000000";
					when "00000100011111001" => rgb <= "000000";
					when "00000100011111010" => rgb <= "000000";
					when "00000100011111011" => rgb <= "000000";
					when "00000100011111100" => rgb <= "000000";
					when "00000100011111101" => rgb <= "000000";
					when "00000100011111110" => rgb <= "000000";
					when "00000100011111111" => rgb <= "000000";
					when "00000100100000000" => rgb <= "000000";
					when "00000100100000001" => rgb <= "000000";
					when "00000100100000010" => rgb <= "000000";
					when "00000100100000011" => rgb <= "000000";
					when "00000100100000100" => rgb <= "000000";
					when "00000100100000101" => rgb <= "000000";
					when "00000100100000110" => rgb <= "000000";
					when "00000100100000111" => rgb <= "000000";
					when "00000100100001000" => rgb <= "000000";
					when "00000100100001001" => rgb <= "000000";
					when "00000100100001010" => rgb <= "000000";
					when "00000100100001011" => rgb <= "000000";
					when "00000100100001100" => rgb <= "000000";
					when "00000100100001101" => rgb <= "000000";
					when "00000100100001110" => rgb <= "000000";
					when "00000100100001111" => rgb <= "000000";
					when "00000100100010000" => rgb <= "000000";
					when "00000100100010001" => rgb <= "000000";
					when "00000100100010010" => rgb <= "000000";
					when "00000100100010011" => rgb <= "000000";
					when "00000100100010100" => rgb <= "000000";
					when "00000100100010101" => rgb <= "000000";
					when "00000100100010110" => rgb <= "000000";
					when "00000100100010111" => rgb <= "000000";
					when "00000100100011000" => rgb <= "000000";
					when "00000100100011001" => rgb <= "000000";
					when "00000100100011010" => rgb <= "000000";
					when "00000100100011011" => rgb <= "000000";
					when "00000100100011100" => rgb <= "000000";
					when "00000100100011101" => rgb <= "000000";
					when "00000100100011110" => rgb <= "000000";
					when "00000100100011111" => rgb <= "000000";
					when "00000100100100000" => rgb <= "000000";
					when "00000100100100001" => rgb <= "000000";
					when "00000100100100010" => rgb <= "000000";
					when "00000100100100011" => rgb <= "000000";
					when "00000100100100100" => rgb <= "000000";
					when "00000100100100101" => rgb <= "000000";
					when "00000100100100110" => rgb <= "000000";
					when "00000100100100111" => rgb <= "000000";
					when "00000100100101000" => rgb <= "000000";
					when "00000100100101001" => rgb <= "000000";
					when "00000100100101010" => rgb <= "000000";
					when "00000100100101011" => rgb <= "000000";
					when "00000100100101100" => rgb <= "000000";
					when "00000100100101101" => rgb <= "000000";
					when "00000100100101110" => rgb <= "000000";
					when "00000100100101111" => rgb <= "000000";
					when "00000100100110000" => rgb <= "000000";
					when "00000100100110001" => rgb <= "000000";
					when "00000100100110010" => rgb <= "000000";
					when "00000100100110011" => rgb <= "000000";
					when "00000100100110100" => rgb <= "000000";
					when "00000100100110101" => rgb <= "000000";
					when "00000100100110110" => rgb <= "000000";
					when "00000100100110111" => rgb <= "000000";
					when "00000100100111000" => rgb <= "000000";
					when "00000100100111001" => rgb <= "000000";
					when "00000100100111010" => rgb <= "000000";
					when "00000100100111011" => rgb <= "000000";
					when "00000100100111100" => rgb <= "000000";
					when "00000100100111101" => rgb <= "000000";
					when "00000100100111110" => rgb <= "000000";
					when "00000100100111111" => rgb <= "000000";
					when "00000101000000000" => rgb <= "000000";
					when "00000101000000001" => rgb <= "000000";
					when "00000101000000010" => rgb <= "000000";
					when "00000101000000011" => rgb <= "000000";
					when "00000101000000100" => rgb <= "000000";
					when "00000101000000101" => rgb <= "000000";
					when "00000101000000110" => rgb <= "000000";
					when "00000101000000111" => rgb <= "000000";
					when "00000101000001000" => rgb <= "000000";
					when "00000101000001001" => rgb <= "000000";
					when "00000101000001010" => rgb <= "000000";
					when "00000101000001011" => rgb <= "000000";
					when "00000101000001100" => rgb <= "000000";
					when "00000101000001101" => rgb <= "000000";
					when "00000101000001110" => rgb <= "000000";
					when "00000101000001111" => rgb <= "000000";
					when "00000101000010000" => rgb <= "000000";
					when "00000101000010001" => rgb <= "000000";
					when "00000101000010010" => rgb <= "000000";
					when "00000101000010011" => rgb <= "000000";
					when "00000101000010100" => rgb <= "000000";
					when "00000101000010101" => rgb <= "000000";
					when "00000101000010110" => rgb <= "000000";
					when "00000101000010111" => rgb <= "000000";
					when "00000101000011000" => rgb <= "000000";
					when "00000101000011001" => rgb <= "000000";
					when "00000101000011010" => rgb <= "000000";
					when "00000101000011011" => rgb <= "000000";
					when "00000101000011100" => rgb <= "000000";
					when "00000101000011101" => rgb <= "000000";
					when "00000101000011110" => rgb <= "000000";
					when "00000101000011111" => rgb <= "000000";
					when "00000101000100000" => rgb <= "000000";
					when "00000101000100001" => rgb <= "000000";
					when "00000101000100010" => rgb <= "000000";
					when "00000101000100011" => rgb <= "000000";
					when "00000101000100100" => rgb <= "000000";
					when "00000101000100101" => rgb <= "000000";
					when "00000101000100110" => rgb <= "000000";
					when "00000101000100111" => rgb <= "000000";
					when "00000101000101000" => rgb <= "000000";
					when "00000101000101001" => rgb <= "000000";
					when "00000101000101010" => rgb <= "000000";
					when "00000101000101011" => rgb <= "000000";
					when "00000101000101100" => rgb <= "000000";
					when "00000101000101101" => rgb <= "000000";
					when "00000101000101110" => rgb <= "000000";
					when "00000101000101111" => rgb <= "000000";
					when "00000101000110000" => rgb <= "000000";
					when "00000101000110001" => rgb <= "000000";
					when "00000101000110010" => rgb <= "000000";
					when "00000101000110011" => rgb <= "000000";
					when "00000101000110100" => rgb <= "000000";
					when "00000101000110101" => rgb <= "000000";
					when "00000101000110110" => rgb <= "000000";
					when "00000101000110111" => rgb <= "000000";
					when "00000101000111000" => rgb <= "000000";
					when "00000101000111001" => rgb <= "000000";
					when "00000101000111010" => rgb <= "000000";
					when "00000101000111011" => rgb <= "000000";
					when "00000101000111100" => rgb <= "000000";
					when "00000101000111101" => rgb <= "000000";
					when "00000101000111110" => rgb <= "000000";
					when "00000101000111111" => rgb <= "000000";
					when "00000101001000000" => rgb <= "000000";
					when "00000101001000001" => rgb <= "000000";
					when "00000101001000010" => rgb <= "000000";
					when "00000101001000011" => rgb <= "000000";
					when "00000101001000100" => rgb <= "000000";
					when "00000101001000101" => rgb <= "000000";
					when "00000101001000110" => rgb <= "000000";
					when "00000101001000111" => rgb <= "000000";
					when "00000101001001000" => rgb <= "000000";
					when "00000101001001001" => rgb <= "000000";
					when "00000101001001010" => rgb <= "000000";
					when "00000101001001011" => rgb <= "000000";
					when "00000101001001100" => rgb <= "000000";
					when "00000101001001101" => rgb <= "000000";
					when "00000101001001110" => rgb <= "000000";
					when "00000101001001111" => rgb <= "000000";
					when "00000101001010000" => rgb <= "000000";
					when "00000101001010001" => rgb <= "000000";
					when "00000101001010010" => rgb <= "000000";
					when "00000101001010011" => rgb <= "000000";
					when "00000101001010100" => rgb <= "000000";
					when "00000101001010101" => rgb <= "000000";
					when "00000101001010110" => rgb <= "000000";
					when "00000101001010111" => rgb <= "000000";
					when "00000101001011000" => rgb <= "000000";
					when "00000101001011001" => rgb <= "000000";
					when "00000101001011010" => rgb <= "000000";
					when "00000101001011011" => rgb <= "000000";
					when "00000101001011100" => rgb <= "000000";
					when "00000101001011101" => rgb <= "000000";
					when "00000101001011110" => rgb <= "000000";
					when "00000101001011111" => rgb <= "000000";
					when "00000101001100000" => rgb <= "000000";
					when "00000101001100001" => rgb <= "000000";
					when "00000101001100010" => rgb <= "000000";
					when "00000101001100011" => rgb <= "000000";
					when "00000101001100100" => rgb <= "000000";
					when "00000101001100101" => rgb <= "000000";
					when "00000101001100110" => rgb <= "000000";
					when "00000101001100111" => rgb <= "000000";
					when "00000101001101000" => rgb <= "000000";
					when "00000101001101001" => rgb <= "000000";
					when "00000101001101010" => rgb <= "000000";
					when "00000101001101011" => rgb <= "000000";
					when "00000101001101100" => rgb <= "000000";
					when "00000101001101101" => rgb <= "000000";
					when "00000101001101110" => rgb <= "000000";
					when "00000101001101111" => rgb <= "000000";
					when "00000101001110000" => rgb <= "000000";
					when "00000101001110001" => rgb <= "000000";
					when "00000101001110010" => rgb <= "000000";
					when "00000101001110011" => rgb <= "000000";
					when "00000101001110100" => rgb <= "000000";
					when "00000101001110101" => rgb <= "000000";
					when "00000101001110110" => rgb <= "000000";
					when "00000101001110111" => rgb <= "000000";
					when "00000101001111000" => rgb <= "000000";
					when "00000101001111001" => rgb <= "000000";
					when "00000101001111010" => rgb <= "000000";
					when "00000101001111011" => rgb <= "000000";
					when "00000101001111100" => rgb <= "000000";
					when "00000101001111101" => rgb <= "000000";
					when "00000101001111110" => rgb <= "000000";
					when "00000101001111111" => rgb <= "000000";
					when "00000101010000000" => rgb <= "000000";
					when "00000101010000001" => rgb <= "000000";
					when "00000101010000010" => rgb <= "000000";
					when "00000101010000011" => rgb <= "000000";
					when "00000101010000100" => rgb <= "000000";
					when "00000101010000101" => rgb <= "000000";
					when "00000101010000110" => rgb <= "000000";
					when "00000101010000111" => rgb <= "000000";
					when "00000101010001000" => rgb <= "000000";
					when "00000101010001001" => rgb <= "000000";
					when "00000101010001010" => rgb <= "000000";
					when "00000101010001011" => rgb <= "000000";
					when "00000101010001100" => rgb <= "000000";
					when "00000101010001101" => rgb <= "000000";
					when "00000101010001110" => rgb <= "000000";
					when "00000101010001111" => rgb <= "000000";
					when "00000101010010000" => rgb <= "000000";
					when "00000101010010001" => rgb <= "000000";
					when "00000101010010010" => rgb <= "000000";
					when "00000101010010011" => rgb <= "000000";
					when "00000101010010100" => rgb <= "000000";
					when "00000101010010101" => rgb <= "000000";
					when "00000101010010110" => rgb <= "000000";
					when "00000101010010111" => rgb <= "000000";
					when "00000101010011000" => rgb <= "000000";
					when "00000101010011001" => rgb <= "000000";
					when "00000101010011010" => rgb <= "000000";
					when "00000101010011011" => rgb <= "000000";
					when "00000101010011100" => rgb <= "000000";
					when "00000101010011101" => rgb <= "000000";
					when "00000101010011110" => rgb <= "000000";
					when "00000101010011111" => rgb <= "000000";
					when "00000101010100000" => rgb <= "000000";
					when "00000101010100001" => rgb <= "000000";
					when "00000101010100010" => rgb <= "000000";
					when "00000101010100011" => rgb <= "000000";
					when "00000101010100100" => rgb <= "000000";
					when "00000101010100101" => rgb <= "000000";
					when "00000101010100110" => rgb <= "000000";
					when "00000101010100111" => rgb <= "000000";
					when "00000101010101000" => rgb <= "000000";
					when "00000101010101001" => rgb <= "000000";
					when "00000101010101010" => rgb <= "000000";
					when "00000101010101011" => rgb <= "000000";
					when "00000101010101100" => rgb <= "000000";
					when "00000101010101101" => rgb <= "000000";
					when "00000101010101110" => rgb <= "000000";
					when "00000101010101111" => rgb <= "000000";
					when "00000101010110000" => rgb <= "000000";
					when "00000101010110001" => rgb <= "000000";
					when "00000101010110010" => rgb <= "000000";
					when "00000101010110011" => rgb <= "000000";
					when "00000101010110100" => rgb <= "000000";
					when "00000101010110101" => rgb <= "000000";
					when "00000101010110110" => rgb <= "000000";
					when "00000101010110111" => rgb <= "000000";
					when "00000101010111000" => rgb <= "000000";
					when "00000101010111001" => rgb <= "000000";
					when "00000101010111010" => rgb <= "000000";
					when "00000101010111011" => rgb <= "000000";
					when "00000101010111100" => rgb <= "000000";
					when "00000101010111101" => rgb <= "000000";
					when "00000101010111110" => rgb <= "000000";
					when "00000101010111111" => rgb <= "000000";
					when "00000101011000000" => rgb <= "000000";
					when "00000101011000001" => rgb <= "000000";
					when "00000101011000010" => rgb <= "000000";
					when "00000101011000011" => rgb <= "000000";
					when "00000101011000100" => rgb <= "000000";
					when "00000101011000101" => rgb <= "000000";
					when "00000101011000110" => rgb <= "000000";
					when "00000101011000111" => rgb <= "000000";
					when "00000101011001000" => rgb <= "000000";
					when "00000101011001001" => rgb <= "000000";
					when "00000101011001010" => rgb <= "000000";
					when "00000101011001011" => rgb <= "000000";
					when "00000101011001100" => rgb <= "000000";
					when "00000101011001101" => rgb <= "000000";
					when "00000101011001110" => rgb <= "000000";
					when "00000101011001111" => rgb <= "000000";
					when "00000101011010000" => rgb <= "000000";
					when "00000101011010001" => rgb <= "000000";
					when "00000101011010010" => rgb <= "000000";
					when "00000101011010011" => rgb <= "000000";
					when "00000101011010100" => rgb <= "000000";
					when "00000101011010101" => rgb <= "000000";
					when "00000101011010110" => rgb <= "000000";
					when "00000101011010111" => rgb <= "000000";
					when "00000101011011000" => rgb <= "000000";
					when "00000101011011001" => rgb <= "000000";
					when "00000101011011010" => rgb <= "000000";
					when "00000101011011011" => rgb <= "000000";
					when "00000101011011100" => rgb <= "000000";
					when "00000101011011101" => rgb <= "000000";
					when "00000101011011110" => rgb <= "000000";
					when "00000101011011111" => rgb <= "000000";
					when "00000101011100000" => rgb <= "000000";
					when "00000101011100001" => rgb <= "000000";
					when "00000101011100010" => rgb <= "000000";
					when "00000101011100011" => rgb <= "000000";
					when "00000101011100100" => rgb <= "000000";
					when "00000101011100101" => rgb <= "000000";
					when "00000101011100110" => rgb <= "000000";
					when "00000101011100111" => rgb <= "000000";
					when "00000101011101000" => rgb <= "000000";
					when "00000101011101001" => rgb <= "000000";
					when "00000101011101010" => rgb <= "000000";
					when "00000101011101011" => rgb <= "000000";
					when "00000101011101100" => rgb <= "000000";
					when "00000101011101101" => rgb <= "000000";
					when "00000101011101110" => rgb <= "000000";
					when "00000101011101111" => rgb <= "000000";
					when "00000101011110000" => rgb <= "000000";
					when "00000101011110001" => rgb <= "000000";
					when "00000101011110010" => rgb <= "000000";
					when "00000101011110011" => rgb <= "000000";
					when "00000101011110100" => rgb <= "000000";
					when "00000101011110101" => rgb <= "000000";
					when "00000101011110110" => rgb <= "000000";
					when "00000101011110111" => rgb <= "000000";
					when "00000101011111000" => rgb <= "000000";
					when "00000101011111001" => rgb <= "000000";
					when "00000101011111010" => rgb <= "000000";
					when "00000101011111011" => rgb <= "000000";
					when "00000101011111100" => rgb <= "000000";
					when "00000101011111101" => rgb <= "000000";
					when "00000101011111110" => rgb <= "000000";
					when "00000101011111111" => rgb <= "000000";
					when "00000101100000000" => rgb <= "000000";
					when "00000101100000001" => rgb <= "000000";
					when "00000101100000010" => rgb <= "000000";
					when "00000101100000011" => rgb <= "000000";
					when "00000101100000100" => rgb <= "000000";
					when "00000101100000101" => rgb <= "000000";
					when "00000101100000110" => rgb <= "000000";
					when "00000101100000111" => rgb <= "000000";
					when "00000101100001000" => rgb <= "000000";
					when "00000101100001001" => rgb <= "000000";
					when "00000101100001010" => rgb <= "000000";
					when "00000101100001011" => rgb <= "000000";
					when "00000101100001100" => rgb <= "000000";
					when "00000101100001101" => rgb <= "000000";
					when "00000101100001110" => rgb <= "000000";
					when "00000101100001111" => rgb <= "000000";
					when "00000101100010000" => rgb <= "000000";
					when "00000101100010001" => rgb <= "000000";
					when "00000101100010010" => rgb <= "000000";
					when "00000101100010011" => rgb <= "000000";
					when "00000101100010100" => rgb <= "000000";
					when "00000101100010101" => rgb <= "000000";
					when "00000101100010110" => rgb <= "000000";
					when "00000101100010111" => rgb <= "000000";
					when "00000101100011000" => rgb <= "000000";
					when "00000101100011001" => rgb <= "000000";
					when "00000101100011010" => rgb <= "000000";
					when "00000101100011011" => rgb <= "000000";
					when "00000101100011100" => rgb <= "000000";
					when "00000101100011101" => rgb <= "000000";
					when "00000101100011110" => rgb <= "000000";
					when "00000101100011111" => rgb <= "000000";
					when "00000101100100000" => rgb <= "000000";
					when "00000101100100001" => rgb <= "000000";
					when "00000101100100010" => rgb <= "000000";
					when "00000101100100011" => rgb <= "000000";
					when "00000101100100100" => rgb <= "000000";
					when "00000101100100101" => rgb <= "000000";
					when "00000101100100110" => rgb <= "000000";
					when "00000101100100111" => rgb <= "000000";
					when "00000101100101000" => rgb <= "000000";
					when "00000101100101001" => rgb <= "000000";
					when "00000101100101010" => rgb <= "000000";
					when "00000101100101011" => rgb <= "000000";
					when "00000101100101100" => rgb <= "000000";
					when "00000101100101101" => rgb <= "000000";
					when "00000101100101110" => rgb <= "000000";
					when "00000101100101111" => rgb <= "000000";
					when "00000101100110000" => rgb <= "000000";
					when "00000101100110001" => rgb <= "000000";
					when "00000101100110010" => rgb <= "000000";
					when "00000101100110011" => rgb <= "000000";
					when "00000101100110100" => rgb <= "000000";
					when "00000101100110101" => rgb <= "000000";
					when "00000101100110110" => rgb <= "000000";
					when "00000101100110111" => rgb <= "000000";
					when "00000101100111000" => rgb <= "000000";
					when "00000101100111001" => rgb <= "000000";
					when "00000101100111010" => rgb <= "000000";
					when "00000101100111011" => rgb <= "000000";
					when "00000101100111100" => rgb <= "000000";
					when "00000101100111101" => rgb <= "000000";
					when "00000101100111110" => rgb <= "000000";
					when "00000101100111111" => rgb <= "000000";
					when "00000110000000000" => rgb <= "000000";
					when "00000110000000001" => rgb <= "000000";
					when "00000110000000010" => rgb <= "000000";
					when "00000110000000011" => rgb <= "000000";
					when "00000110000000100" => rgb <= "000000";
					when "00000110000000101" => rgb <= "000000";
					when "00000110000000110" => rgb <= "000000";
					when "00000110000000111" => rgb <= "000000";
					when "00000110000001000" => rgb <= "000000";
					when "00000110000001001" => rgb <= "000000";
					when "00000110000001010" => rgb <= "000000";
					when "00000110000001011" => rgb <= "000000";
					when "00000110000001100" => rgb <= "000000";
					when "00000110000001101" => rgb <= "000000";
					when "00000110000001110" => rgb <= "000000";
					when "00000110000001111" => rgb <= "000000";
					when "00000110000010000" => rgb <= "000000";
					when "00000110000010001" => rgb <= "000000";
					when "00000110000010010" => rgb <= "000000";
					when "00000110000010011" => rgb <= "000000";
					when "00000110000010100" => rgb <= "000000";
					when "00000110000010101" => rgb <= "000000";
					when "00000110000010110" => rgb <= "000000";
					when "00000110000010111" => rgb <= "000000";
					when "00000110000011000" => rgb <= "000000";
					when "00000110000011001" => rgb <= "000000";
					when "00000110000011010" => rgb <= "000000";
					when "00000110000011011" => rgb <= "000000";
					when "00000110000011100" => rgb <= "000000";
					when "00000110000011101" => rgb <= "000000";
					when "00000110000011110" => rgb <= "000000";
					when "00000110000011111" => rgb <= "000000";
					when "00000110000100000" => rgb <= "000000";
					when "00000110000100001" => rgb <= "000000";
					when "00000110000100010" => rgb <= "000000";
					when "00000110000100011" => rgb <= "000000";
					when "00000110000100100" => rgb <= "000000";
					when "00000110000100101" => rgb <= "000000";
					when "00000110000100110" => rgb <= "000000";
					when "00000110000100111" => rgb <= "000000";
					when "00000110000101000" => rgb <= "000000";
					when "00000110000101001" => rgb <= "000000";
					when "00000110000101010" => rgb <= "000000";
					when "00000110000101011" => rgb <= "000000";
					when "00000110000101100" => rgb <= "000000";
					when "00000110000101101" => rgb <= "000000";
					when "00000110000101110" => rgb <= "000000";
					when "00000110000101111" => rgb <= "000000";
					when "00000110000110000" => rgb <= "000000";
					when "00000110000110001" => rgb <= "000000";
					when "00000110000110010" => rgb <= "000000";
					when "00000110000110011" => rgb <= "000000";
					when "00000110000110100" => rgb <= "000000";
					when "00000110000110101" => rgb <= "000000";
					when "00000110000110110" => rgb <= "000000";
					when "00000110000110111" => rgb <= "000000";
					when "00000110000111000" => rgb <= "000000";
					when "00000110000111001" => rgb <= "000000";
					when "00000110000111010" => rgb <= "000000";
					when "00000110000111011" => rgb <= "000000";
					when "00000110000111100" => rgb <= "000000";
					when "00000110000111101" => rgb <= "000000";
					when "00000110000111110" => rgb <= "000000";
					when "00000110000111111" => rgb <= "000000";
					when "00000110001000000" => rgb <= "000000";
					when "00000110001000001" => rgb <= "000000";
					when "00000110001000010" => rgb <= "000000";
					when "00000110001000011" => rgb <= "000000";
					when "00000110001000100" => rgb <= "000000";
					when "00000110001000101" => rgb <= "000000";
					when "00000110001000110" => rgb <= "000000";
					when "00000110001000111" => rgb <= "000000";
					when "00000110001001000" => rgb <= "000000";
					when "00000110001001001" => rgb <= "000000";
					when "00000110001001010" => rgb <= "000000";
					when "00000110001001011" => rgb <= "000000";
					when "00000110001001100" => rgb <= "000000";
					when "00000110001001101" => rgb <= "000000";
					when "00000110001001110" => rgb <= "000000";
					when "00000110001001111" => rgb <= "000000";
					when "00000110001010000" => rgb <= "000000";
					when "00000110001010001" => rgb <= "000000";
					when "00000110001010010" => rgb <= "000000";
					when "00000110001010011" => rgb <= "000000";
					when "00000110001010100" => rgb <= "000000";
					when "00000110001010101" => rgb <= "000000";
					when "00000110001010110" => rgb <= "000000";
					when "00000110001010111" => rgb <= "000000";
					when "00000110001011000" => rgb <= "000000";
					when "00000110001011001" => rgb <= "000000";
					when "00000110001011010" => rgb <= "000000";
					when "00000110001011011" => rgb <= "000000";
					when "00000110001011100" => rgb <= "000000";
					when "00000110001011101" => rgb <= "000000";
					when "00000110001011110" => rgb <= "000000";
					when "00000110001011111" => rgb <= "000000";
					when "00000110001100000" => rgb <= "000000";
					when "00000110001100001" => rgb <= "000000";
					when "00000110001100010" => rgb <= "000000";
					when "00000110001100011" => rgb <= "000000";
					when "00000110001100100" => rgb <= "000000";
					when "00000110001100101" => rgb <= "000000";
					when "00000110001100110" => rgb <= "000000";
					when "00000110001100111" => rgb <= "000000";
					when "00000110001101000" => rgb <= "000000";
					when "00000110001101001" => rgb <= "000000";
					when "00000110001101010" => rgb <= "000000";
					when "00000110001101011" => rgb <= "000000";
					when "00000110001101100" => rgb <= "000000";
					when "00000110001101101" => rgb <= "000000";
					when "00000110001101110" => rgb <= "000000";
					when "00000110001101111" => rgb <= "000000";
					when "00000110001110000" => rgb <= "000000";
					when "00000110001110001" => rgb <= "000000";
					when "00000110001110010" => rgb <= "000000";
					when "00000110001110011" => rgb <= "000000";
					when "00000110001110100" => rgb <= "000000";
					when "00000110001110101" => rgb <= "000000";
					when "00000110001110110" => rgb <= "000000";
					when "00000110001110111" => rgb <= "000000";
					when "00000110001111000" => rgb <= "000000";
					when "00000110001111001" => rgb <= "000000";
					when "00000110001111010" => rgb <= "000000";
					when "00000110001111011" => rgb <= "000000";
					when "00000110001111100" => rgb <= "000000";
					when "00000110001111101" => rgb <= "000000";
					when "00000110001111110" => rgb <= "000000";
					when "00000110001111111" => rgb <= "000000";
					when "00000110010000000" => rgb <= "000000";
					when "00000110010000001" => rgb <= "000000";
					when "00000110010000010" => rgb <= "000000";
					when "00000110010000011" => rgb <= "000000";
					when "00000110010000100" => rgb <= "000000";
					when "00000110010000101" => rgb <= "000000";
					when "00000110010000110" => rgb <= "000000";
					when "00000110010000111" => rgb <= "000000";
					when "00000110010001000" => rgb <= "000000";
					when "00000110010001001" => rgb <= "000000";
					when "00000110010001010" => rgb <= "000000";
					when "00000110010001011" => rgb <= "000000";
					when "00000110010001100" => rgb <= "000000";
					when "00000110010001101" => rgb <= "000000";
					when "00000110010001110" => rgb <= "000000";
					when "00000110010001111" => rgb <= "000000";
					when "00000110010010000" => rgb <= "000000";
					when "00000110010010001" => rgb <= "000000";
					when "00000110010010010" => rgb <= "000000";
					when "00000110010010011" => rgb <= "000000";
					when "00000110010010100" => rgb <= "000000";
					when "00000110010010101" => rgb <= "000000";
					when "00000110010010110" => rgb <= "000000";
					when "00000110010010111" => rgb <= "000000";
					when "00000110010011000" => rgb <= "000000";
					when "00000110010011001" => rgb <= "000000";
					when "00000110010011010" => rgb <= "000000";
					when "00000110010011011" => rgb <= "000000";
					when "00000110010011100" => rgb <= "000000";
					when "00000110010011101" => rgb <= "000000";
					when "00000110010011110" => rgb <= "000000";
					when "00000110010011111" => rgb <= "000000";
					when "00000110010100000" => rgb <= "000000";
					when "00000110010100001" => rgb <= "000000";
					when "00000110010100010" => rgb <= "000000";
					when "00000110010100011" => rgb <= "000000";
					when "00000110010100100" => rgb <= "000000";
					when "00000110010100101" => rgb <= "000000";
					when "00000110010100110" => rgb <= "000000";
					when "00000110010100111" => rgb <= "000000";
					when "00000110010101000" => rgb <= "000000";
					when "00000110010101001" => rgb <= "000000";
					when "00000110010101010" => rgb <= "000000";
					when "00000110010101011" => rgb <= "000000";
					when "00000110010101100" => rgb <= "000000";
					when "00000110010101101" => rgb <= "000000";
					when "00000110010101110" => rgb <= "000000";
					when "00000110010101111" => rgb <= "000000";
					when "00000110010110000" => rgb <= "000000";
					when "00000110010110001" => rgb <= "000000";
					when "00000110010110010" => rgb <= "000000";
					when "00000110010110011" => rgb <= "000000";
					when "00000110010110100" => rgb <= "000000";
					when "00000110010110101" => rgb <= "000000";
					when "00000110010110110" => rgb <= "000000";
					when "00000110010110111" => rgb <= "000000";
					when "00000110010111000" => rgb <= "000000";
					when "00000110010111001" => rgb <= "000000";
					when "00000110010111010" => rgb <= "000000";
					when "00000110010111011" => rgb <= "000000";
					when "00000110010111100" => rgb <= "000000";
					when "00000110010111101" => rgb <= "000000";
					when "00000110010111110" => rgb <= "000000";
					when "00000110010111111" => rgb <= "000000";
					when "00000110011000000" => rgb <= "000000";
					when "00000110011000001" => rgb <= "000000";
					when "00000110011000010" => rgb <= "000000";
					when "00000110011000011" => rgb <= "000000";
					when "00000110011000100" => rgb <= "000000";
					when "00000110011000101" => rgb <= "000000";
					when "00000110011000110" => rgb <= "000000";
					when "00000110011000111" => rgb <= "000000";
					when "00000110011001000" => rgb <= "000000";
					when "00000110011001001" => rgb <= "000000";
					when "00000110011001010" => rgb <= "000000";
					when "00000110011001011" => rgb <= "000000";
					when "00000110011001100" => rgb <= "000000";
					when "00000110011001101" => rgb <= "000000";
					when "00000110011001110" => rgb <= "000000";
					when "00000110011001111" => rgb <= "000000";
					when "00000110011010000" => rgb <= "000000";
					when "00000110011010001" => rgb <= "000000";
					when "00000110011010010" => rgb <= "000000";
					when "00000110011010011" => rgb <= "000000";
					when "00000110011010100" => rgb <= "000000";
					when "00000110011010101" => rgb <= "000000";
					when "00000110011010110" => rgb <= "000000";
					when "00000110011010111" => rgb <= "000000";
					when "00000110011011000" => rgb <= "000000";
					when "00000110011011001" => rgb <= "000000";
					when "00000110011011010" => rgb <= "000000";
					when "00000110011011011" => rgb <= "000000";
					when "00000110011011100" => rgb <= "000000";
					when "00000110011011101" => rgb <= "000000";
					when "00000110011011110" => rgb <= "000000";
					when "00000110011011111" => rgb <= "000000";
					when "00000110011100000" => rgb <= "000000";
					when "00000110011100001" => rgb <= "000000";
					when "00000110011100010" => rgb <= "000000";
					when "00000110011100011" => rgb <= "000000";
					when "00000110011100100" => rgb <= "000000";
					when "00000110011100101" => rgb <= "000000";
					when "00000110011100110" => rgb <= "000000";
					when "00000110011100111" => rgb <= "000000";
					when "00000110011101000" => rgb <= "000000";
					when "00000110011101001" => rgb <= "000000";
					when "00000110011101010" => rgb <= "000000";
					when "00000110011101011" => rgb <= "000000";
					when "00000110011101100" => rgb <= "000000";
					when "00000110011101101" => rgb <= "000000";
					when "00000110011101110" => rgb <= "000000";
					when "00000110011101111" => rgb <= "000000";
					when "00000110011110000" => rgb <= "000000";
					when "00000110011110001" => rgb <= "000000";
					when "00000110011110010" => rgb <= "000000";
					when "00000110011110011" => rgb <= "000000";
					when "00000110011110100" => rgb <= "000000";
					when "00000110011110101" => rgb <= "000000";
					when "00000110011110110" => rgb <= "000000";
					when "00000110011110111" => rgb <= "000000";
					when "00000110011111000" => rgb <= "000000";
					when "00000110011111001" => rgb <= "000000";
					when "00000110011111010" => rgb <= "000000";
					when "00000110011111011" => rgb <= "000000";
					when "00000110011111100" => rgb <= "000000";
					when "00000110011111101" => rgb <= "000000";
					when "00000110011111110" => rgb <= "000000";
					when "00000110011111111" => rgb <= "000000";
					when "00000110100000000" => rgb <= "000000";
					when "00000110100000001" => rgb <= "000000";
					when "00000110100000010" => rgb <= "000000";
					when "00000110100000011" => rgb <= "000000";
					when "00000110100000100" => rgb <= "000000";
					when "00000110100000101" => rgb <= "000000";
					when "00000110100000110" => rgb <= "000000";
					when "00000110100000111" => rgb <= "000000";
					when "00000110100001000" => rgb <= "000000";
					when "00000110100001001" => rgb <= "000000";
					when "00000110100001010" => rgb <= "000000";
					when "00000110100001011" => rgb <= "000000";
					when "00000110100001100" => rgb <= "000000";
					when "00000110100001101" => rgb <= "000000";
					when "00000110100001110" => rgb <= "000000";
					when "00000110100001111" => rgb <= "000000";
					when "00000110100010000" => rgb <= "000000";
					when "00000110100010001" => rgb <= "000000";
					when "00000110100010010" => rgb <= "000000";
					when "00000110100010011" => rgb <= "000000";
					when "00000110100010100" => rgb <= "000000";
					when "00000110100010101" => rgb <= "000000";
					when "00000110100010110" => rgb <= "000000";
					when "00000110100010111" => rgb <= "000000";
					when "00000110100011000" => rgb <= "000000";
					when "00000110100011001" => rgb <= "000000";
					when "00000110100011010" => rgb <= "000000";
					when "00000110100011011" => rgb <= "000000";
					when "00000110100011100" => rgb <= "000000";
					when "00000110100011101" => rgb <= "000000";
					when "00000110100011110" => rgb <= "000000";
					when "00000110100011111" => rgb <= "000000";
					when "00000110100100000" => rgb <= "000000";
					when "00000110100100001" => rgb <= "000000";
					when "00000110100100010" => rgb <= "000000";
					when "00000110100100011" => rgb <= "000000";
					when "00000110100100100" => rgb <= "000000";
					when "00000110100100101" => rgb <= "000000";
					when "00000110100100110" => rgb <= "000000";
					when "00000110100100111" => rgb <= "000000";
					when "00000110100101000" => rgb <= "000000";
					when "00000110100101001" => rgb <= "000000";
					when "00000110100101010" => rgb <= "000000";
					when "00000110100101011" => rgb <= "000000";
					when "00000110100101100" => rgb <= "000000";
					when "00000110100101101" => rgb <= "000000";
					when "00000110100101110" => rgb <= "000000";
					when "00000110100101111" => rgb <= "000000";
					when "00000110100110000" => rgb <= "000000";
					when "00000110100110001" => rgb <= "000000";
					when "00000110100110010" => rgb <= "000000";
					when "00000110100110011" => rgb <= "000000";
					when "00000110100110100" => rgb <= "000000";
					when "00000110100110101" => rgb <= "000000";
					when "00000110100110110" => rgb <= "000000";
					when "00000110100110111" => rgb <= "000000";
					when "00000110100111000" => rgb <= "000000";
					when "00000110100111001" => rgb <= "000000";
					when "00000110100111010" => rgb <= "000000";
					when "00000110100111011" => rgb <= "000000";
					when "00000110100111100" => rgb <= "000000";
					when "00000110100111101" => rgb <= "000000";
					when "00000110100111110" => rgb <= "000000";
					when "00000110100111111" => rgb <= "000000";
					when "00000111000000000" => rgb <= "000000";
					when "00000111000000001" => rgb <= "000000";
					when "00000111000000010" => rgb <= "000000";
					when "00000111000000011" => rgb <= "000000";
					when "00000111000000100" => rgb <= "000000";
					when "00000111000000101" => rgb <= "000000";
					when "00000111000000110" => rgb <= "000000";
					when "00000111000000111" => rgb <= "000000";
					when "00000111000001000" => rgb <= "000000";
					when "00000111000001001" => rgb <= "000000";
					when "00000111000001010" => rgb <= "000000";
					when "00000111000001011" => rgb <= "000000";
					when "00000111000001100" => rgb <= "000000";
					when "00000111000001101" => rgb <= "000000";
					when "00000111000001110" => rgb <= "000000";
					when "00000111000001111" => rgb <= "000000";
					when "00000111000010000" => rgb <= "000000";
					when "00000111000010001" => rgb <= "000000";
					when "00000111000010010" => rgb <= "000000";
					when "00000111000010011" => rgb <= "000000";
					when "00000111000010100" => rgb <= "000000";
					when "00000111000010101" => rgb <= "000000";
					when "00000111000010110" => rgb <= "000000";
					when "00000111000010111" => rgb <= "000000";
					when "00000111000011000" => rgb <= "000000";
					when "00000111000011001" => rgb <= "000000";
					when "00000111000011010" => rgb <= "000000";
					when "00000111000011011" => rgb <= "000000";
					when "00000111000011100" => rgb <= "000000";
					when "00000111000011101" => rgb <= "000000";
					when "00000111000011110" => rgb <= "000000";
					when "00000111000011111" => rgb <= "000000";
					when "00000111000100000" => rgb <= "000000";
					when "00000111000100001" => rgb <= "000000";
					when "00000111000100010" => rgb <= "000000";
					when "00000111000100011" => rgb <= "000000";
					when "00000111000100100" => rgb <= "000000";
					when "00000111000100101" => rgb <= "000000";
					when "00000111000100110" => rgb <= "000000";
					when "00000111000100111" => rgb <= "000000";
					when "00000111000101000" => rgb <= "000000";
					when "00000111000101001" => rgb <= "000000";
					when "00000111000101010" => rgb <= "000000";
					when "00000111000101011" => rgb <= "000000";
					when "00000111000101100" => rgb <= "000000";
					when "00000111000101101" => rgb <= "000000";
					when "00000111000101110" => rgb <= "000000";
					when "00000111000101111" => rgb <= "000000";
					when "00000111000110000" => rgb <= "000000";
					when "00000111000110001" => rgb <= "000000";
					when "00000111000110010" => rgb <= "000000";
					when "00000111000110011" => rgb <= "000000";
					when "00000111000110100" => rgb <= "000000";
					when "00000111000110101" => rgb <= "000000";
					when "00000111000110110" => rgb <= "000000";
					when "00000111000110111" => rgb <= "000000";
					when "00000111000111000" => rgb <= "000000";
					when "00000111000111001" => rgb <= "000000";
					when "00000111000111010" => rgb <= "000000";
					when "00000111000111011" => rgb <= "000000";
					when "00000111000111100" => rgb <= "000000";
					when "00000111000111101" => rgb <= "000000";
					when "00000111000111110" => rgb <= "000000";
					when "00000111000111111" => rgb <= "000000";
					when "00000111001000000" => rgb <= "000000";
					when "00000111001000001" => rgb <= "000000";
					when "00000111001000010" => rgb <= "000000";
					when "00000111001000011" => rgb <= "000000";
					when "00000111001000100" => rgb <= "000000";
					when "00000111001000101" => rgb <= "000000";
					when "00000111001000110" => rgb <= "000000";
					when "00000111001000111" => rgb <= "000000";
					when "00000111001001000" => rgb <= "000000";
					when "00000111001001001" => rgb <= "000000";
					when "00000111001001010" => rgb <= "000000";
					when "00000111001001011" => rgb <= "000000";
					when "00000111001001100" => rgb <= "000000";
					when "00000111001001101" => rgb <= "000000";
					when "00000111001001110" => rgb <= "000000";
					when "00000111001001111" => rgb <= "000000";
					when "00000111001010000" => rgb <= "000000";
					when "00000111001010001" => rgb <= "000000";
					when "00000111001010010" => rgb <= "000000";
					when "00000111001010011" => rgb <= "000000";
					when "00000111001010100" => rgb <= "000000";
					when "00000111001010101" => rgb <= "000000";
					when "00000111001010110" => rgb <= "000000";
					when "00000111001010111" => rgb <= "000000";
					when "00000111001011000" => rgb <= "000000";
					when "00000111001011001" => rgb <= "000000";
					when "00000111001011010" => rgb <= "000000";
					when "00000111001011011" => rgb <= "000000";
					when "00000111001011100" => rgb <= "000000";
					when "00000111001011101" => rgb <= "000000";
					when "00000111001011110" => rgb <= "000000";
					when "00000111001011111" => rgb <= "000000";
					when "00000111001100000" => rgb <= "000000";
					when "00000111001100001" => rgb <= "000000";
					when "00000111001100010" => rgb <= "000000";
					when "00000111001100011" => rgb <= "000000";
					when "00000111001100100" => rgb <= "000000";
					when "00000111001100101" => rgb <= "000000";
					when "00000111001100110" => rgb <= "000000";
					when "00000111001100111" => rgb <= "000000";
					when "00000111001101000" => rgb <= "000000";
					when "00000111001101001" => rgb <= "000000";
					when "00000111001101010" => rgb <= "000000";
					when "00000111001101011" => rgb <= "000000";
					when "00000111001101100" => rgb <= "000000";
					when "00000111001101101" => rgb <= "000000";
					when "00000111001101110" => rgb <= "000000";
					when "00000111001101111" => rgb <= "000000";
					when "00000111001110000" => rgb <= "000000";
					when "00000111001110001" => rgb <= "000000";
					when "00000111001110010" => rgb <= "000000";
					when "00000111001110011" => rgb <= "000000";
					when "00000111001110100" => rgb <= "000000";
					when "00000111001110101" => rgb <= "000000";
					when "00000111001110110" => rgb <= "000000";
					when "00000111001110111" => rgb <= "000000";
					when "00000111001111000" => rgb <= "000000";
					when "00000111001111001" => rgb <= "000000";
					when "00000111001111010" => rgb <= "000000";
					when "00000111001111011" => rgb <= "000000";
					when "00000111001111100" => rgb <= "000000";
					when "00000111001111101" => rgb <= "000000";
					when "00000111001111110" => rgb <= "000000";
					when "00000111001111111" => rgb <= "000000";
					when "00000111010000000" => rgb <= "000000";
					when "00000111010000001" => rgb <= "000000";
					when "00000111010000010" => rgb <= "000000";
					when "00000111010000011" => rgb <= "000000";
					when "00000111010000100" => rgb <= "000000";
					when "00000111010000101" => rgb <= "000000";
					when "00000111010000110" => rgb <= "000000";
					when "00000111010000111" => rgb <= "000000";
					when "00000111010001000" => rgb <= "000000";
					when "00000111010001001" => rgb <= "000000";
					when "00000111010001010" => rgb <= "000000";
					when "00000111010001011" => rgb <= "000000";
					when "00000111010001100" => rgb <= "000000";
					when "00000111010001101" => rgb <= "000000";
					when "00000111010001110" => rgb <= "000000";
					when "00000111010001111" => rgb <= "000000";
					when "00000111010010000" => rgb <= "000000";
					when "00000111010010001" => rgb <= "000000";
					when "00000111010010010" => rgb <= "000000";
					when "00000111010010011" => rgb <= "000000";
					when "00000111010010100" => rgb <= "000000";
					when "00000111010010101" => rgb <= "000000";
					when "00000111010010110" => rgb <= "000000";
					when "00000111010010111" => rgb <= "000000";
					when "00000111010011000" => rgb <= "000000";
					when "00000111010011001" => rgb <= "000000";
					when "00000111010011010" => rgb <= "000000";
					when "00000111010011011" => rgb <= "000000";
					when "00000111010011100" => rgb <= "000000";
					when "00000111010011101" => rgb <= "000000";
					when "00000111010011110" => rgb <= "000000";
					when "00000111010011111" => rgb <= "000000";
					when "00000111010100000" => rgb <= "000000";
					when "00000111010100001" => rgb <= "000000";
					when "00000111010100010" => rgb <= "000000";
					when "00000111010100011" => rgb <= "000000";
					when "00000111010100100" => rgb <= "000000";
					when "00000111010100101" => rgb <= "000000";
					when "00000111010100110" => rgb <= "000000";
					when "00000111010100111" => rgb <= "000000";
					when "00000111010101000" => rgb <= "000000";
					when "00000111010101001" => rgb <= "000000";
					when "00000111010101010" => rgb <= "000000";
					when "00000111010101011" => rgb <= "000000";
					when "00000111010101100" => rgb <= "000000";
					when "00000111010101101" => rgb <= "000000";
					when "00000111010101110" => rgb <= "000000";
					when "00000111010101111" => rgb <= "000000";
					when "00000111010110000" => rgb <= "000000";
					when "00000111010110001" => rgb <= "000000";
					when "00000111010110010" => rgb <= "000000";
					when "00000111010110011" => rgb <= "000000";
					when "00000111010110100" => rgb <= "000000";
					when "00000111010110101" => rgb <= "000000";
					when "00000111010110110" => rgb <= "000000";
					when "00000111010110111" => rgb <= "000000";
					when "00000111010111000" => rgb <= "000000";
					when "00000111010111001" => rgb <= "000000";
					when "00000111010111010" => rgb <= "000000";
					when "00000111010111011" => rgb <= "000000";
					when "00000111010111100" => rgb <= "000000";
					when "00000111010111101" => rgb <= "000000";
					when "00000111010111110" => rgb <= "000000";
					when "00000111010111111" => rgb <= "000000";
					when "00000111011000000" => rgb <= "000000";
					when "00000111011000001" => rgb <= "000000";
					when "00000111011000010" => rgb <= "000000";
					when "00000111011000011" => rgb <= "000000";
					when "00000111011000100" => rgb <= "000000";
					when "00000111011000101" => rgb <= "000000";
					when "00000111011000110" => rgb <= "000000";
					when "00000111011000111" => rgb <= "000000";
					when "00000111011001000" => rgb <= "000000";
					when "00000111011001001" => rgb <= "000000";
					when "00000111011001010" => rgb <= "000000";
					when "00000111011001011" => rgb <= "000000";
					when "00000111011001100" => rgb <= "000000";
					when "00000111011001101" => rgb <= "000000";
					when "00000111011001110" => rgb <= "000000";
					when "00000111011001111" => rgb <= "000000";
					when "00000111011010000" => rgb <= "000000";
					when "00000111011010001" => rgb <= "000000";
					when "00000111011010010" => rgb <= "000000";
					when "00000111011010011" => rgb <= "000000";
					when "00000111011010100" => rgb <= "000000";
					when "00000111011010101" => rgb <= "000000";
					when "00000111011010110" => rgb <= "000000";
					when "00000111011010111" => rgb <= "000000";
					when "00000111011011000" => rgb <= "000000";
					when "00000111011011001" => rgb <= "000000";
					when "00000111011011010" => rgb <= "000000";
					when "00000111011011011" => rgb <= "000000";
					when "00000111011011100" => rgb <= "000000";
					when "00000111011011101" => rgb <= "000000";
					when "00000111011011110" => rgb <= "000000";
					when "00000111011011111" => rgb <= "000000";
					when "00000111011100000" => rgb <= "000000";
					when "00000111011100001" => rgb <= "000000";
					when "00000111011100010" => rgb <= "000000";
					when "00000111011100011" => rgb <= "000000";
					when "00000111011100100" => rgb <= "000000";
					when "00000111011100101" => rgb <= "000000";
					when "00000111011100110" => rgb <= "000000";
					when "00000111011100111" => rgb <= "000000";
					when "00000111011101000" => rgb <= "000000";
					when "00000111011101001" => rgb <= "000000";
					when "00000111011101010" => rgb <= "000000";
					when "00000111011101011" => rgb <= "000000";
					when "00000111011101100" => rgb <= "000000";
					when "00000111011101101" => rgb <= "000000";
					when "00000111011101110" => rgb <= "000000";
					when "00000111011101111" => rgb <= "000000";
					when "00000111011110000" => rgb <= "000000";
					when "00000111011110001" => rgb <= "000000";
					when "00000111011110010" => rgb <= "000000";
					when "00000111011110011" => rgb <= "000000";
					when "00000111011110100" => rgb <= "000000";
					when "00000111011110101" => rgb <= "000000";
					when "00000111011110110" => rgb <= "000000";
					when "00000111011110111" => rgb <= "000000";
					when "00000111011111000" => rgb <= "000000";
					when "00000111011111001" => rgb <= "000000";
					when "00000111011111010" => rgb <= "000000";
					when "00000111011111011" => rgb <= "000000";
					when "00000111011111100" => rgb <= "000000";
					when "00000111011111101" => rgb <= "000000";
					when "00000111011111110" => rgb <= "000000";
					when "00000111011111111" => rgb <= "000000";
					when "00000111100000000" => rgb <= "000000";
					when "00000111100000001" => rgb <= "000000";
					when "00000111100000010" => rgb <= "000000";
					when "00000111100000011" => rgb <= "000000";
					when "00000111100000100" => rgb <= "000000";
					when "00000111100000101" => rgb <= "000000";
					when "00000111100000110" => rgb <= "000000";
					when "00000111100000111" => rgb <= "000000";
					when "00000111100001000" => rgb <= "000000";
					when "00000111100001001" => rgb <= "000000";
					when "00000111100001010" => rgb <= "000000";
					when "00000111100001011" => rgb <= "000000";
					when "00000111100001100" => rgb <= "000000";
					when "00000111100001101" => rgb <= "000000";
					when "00000111100001110" => rgb <= "000000";
					when "00000111100001111" => rgb <= "000000";
					when "00000111100010000" => rgb <= "000000";
					when "00000111100010001" => rgb <= "000000";
					when "00000111100010010" => rgb <= "000000";
					when "00000111100010011" => rgb <= "000000";
					when "00000111100010100" => rgb <= "000000";
					when "00000111100010101" => rgb <= "000000";
					when "00000111100010110" => rgb <= "000000";
					when "00000111100010111" => rgb <= "000000";
					when "00000111100011000" => rgb <= "000000";
					when "00000111100011001" => rgb <= "000000";
					when "00000111100011010" => rgb <= "000000";
					when "00000111100011011" => rgb <= "000000";
					when "00000111100011100" => rgb <= "000000";
					when "00000111100011101" => rgb <= "000000";
					when "00000111100011110" => rgb <= "000000";
					when "00000111100011111" => rgb <= "000000";
					when "00000111100100000" => rgb <= "000000";
					when "00000111100100001" => rgb <= "000000";
					when "00000111100100010" => rgb <= "000000";
					when "00000111100100011" => rgb <= "000000";
					when "00000111100100100" => rgb <= "000000";
					when "00000111100100101" => rgb <= "000000";
					when "00000111100100110" => rgb <= "000000";
					when "00000111100100111" => rgb <= "000000";
					when "00000111100101000" => rgb <= "000000";
					when "00000111100101001" => rgb <= "000000";
					when "00000111100101010" => rgb <= "000000";
					when "00000111100101011" => rgb <= "000000";
					when "00000111100101100" => rgb <= "000000";
					when "00000111100101101" => rgb <= "000000";
					when "00000111100101110" => rgb <= "000000";
					when "00000111100101111" => rgb <= "000000";
					when "00000111100110000" => rgb <= "000000";
					when "00000111100110001" => rgb <= "000000";
					when "00000111100110010" => rgb <= "000000";
					when "00000111100110011" => rgb <= "000000";
					when "00000111100110100" => rgb <= "000000";
					when "00000111100110101" => rgb <= "000000";
					when "00000111100110110" => rgb <= "000000";
					when "00000111100110111" => rgb <= "000000";
					when "00000111100111000" => rgb <= "000000";
					when "00000111100111001" => rgb <= "000000";
					when "00000111100111010" => rgb <= "000000";
					when "00000111100111011" => rgb <= "000000";
					when "00000111100111100" => rgb <= "000000";
					when "00000111100111101" => rgb <= "000000";
					when "00000111100111110" => rgb <= "000000";
					when "00000111100111111" => rgb <= "000000";
					when "00001000000000000" => rgb <= "000000";
					when "00001000000000001" => rgb <= "000000";
					when "00001000000000010" => rgb <= "000000";
					when "00001000000000011" => rgb <= "000000";
					when "00001000000000100" => rgb <= "000000";
					when "00001000000000101" => rgb <= "000000";
					when "00001000000000110" => rgb <= "000000";
					when "00001000000000111" => rgb <= "000000";
					when "00001000000001000" => rgb <= "000000";
					when "00001000000001001" => rgb <= "000000";
					when "00001000000001010" => rgb <= "000000";
					when "00001000000001011" => rgb <= "000000";
					when "00001000000001100" => rgb <= "000000";
					when "00001000000001101" => rgb <= "000000";
					when "00001000000001110" => rgb <= "000000";
					when "00001000000001111" => rgb <= "000000";
					when "00001000000010000" => rgb <= "000000";
					when "00001000000010001" => rgb <= "000000";
					when "00001000000010010" => rgb <= "000000";
					when "00001000000010011" => rgb <= "000000";
					when "00001000000010100" => rgb <= "000000";
					when "00001000000010101" => rgb <= "000000";
					when "00001000000010110" => rgb <= "000000";
					when "00001000000010111" => rgb <= "000000";
					when "00001000000011000" => rgb <= "000000";
					when "00001000000011001" => rgb <= "000000";
					when "00001000000011010" => rgb <= "000000";
					when "00001000000011011" => rgb <= "000000";
					when "00001000000011100" => rgb <= "000000";
					when "00001000000011101" => rgb <= "000000";
					when "00001000000011110" => rgb <= "000000";
					when "00001000000011111" => rgb <= "000000";
					when "00001000000100000" => rgb <= "000000";
					when "00001000000100001" => rgb <= "000000";
					when "00001000000100010" => rgb <= "000000";
					when "00001000000100011" => rgb <= "000000";
					when "00001000000100100" => rgb <= "000000";
					when "00001000000100101" => rgb <= "000000";
					when "00001000000100110" => rgb <= "000000";
					when "00001000000100111" => rgb <= "000000";
					when "00001000000101000" => rgb <= "000000";
					when "00001000000101001" => rgb <= "000000";
					when "00001000000101010" => rgb <= "000000";
					when "00001000000101011" => rgb <= "000000";
					when "00001000000101100" => rgb <= "000000";
					when "00001000000101101" => rgb <= "000000";
					when "00001000000101110" => rgb <= "000000";
					when "00001000000101111" => rgb <= "000000";
					when "00001000000110000" => rgb <= "000000";
					when "00001000000110001" => rgb <= "000000";
					when "00001000000110010" => rgb <= "000000";
					when "00001000000110011" => rgb <= "000000";
					when "00001000000110100" => rgb <= "000000";
					when "00001000000110101" => rgb <= "000000";
					when "00001000000110110" => rgb <= "000000";
					when "00001000000110111" => rgb <= "000000";
					when "00001000000111000" => rgb <= "000000";
					when "00001000000111001" => rgb <= "000000";
					when "00001000000111010" => rgb <= "000000";
					when "00001000000111011" => rgb <= "000000";
					when "00001000000111100" => rgb <= "000000";
					when "00001000000111101" => rgb <= "000000";
					when "00001000000111110" => rgb <= "000000";
					when "00001000000111111" => rgb <= "000000";
					when "00001000001000000" => rgb <= "000000";
					when "00001000001000001" => rgb <= "000000";
					when "00001000001000010" => rgb <= "000000";
					when "00001000001000011" => rgb <= "000000";
					when "00001000001000100" => rgb <= "000000";
					when "00001000001000101" => rgb <= "000000";
					when "00001000001000110" => rgb <= "000000";
					when "00001000001000111" => rgb <= "000000";
					when "00001000001001000" => rgb <= "000000";
					when "00001000001001001" => rgb <= "000000";
					when "00001000001001010" => rgb <= "000000";
					when "00001000001001011" => rgb <= "000000";
					when "00001000001001100" => rgb <= "000000";
					when "00001000001001101" => rgb <= "000000";
					when "00001000001001110" => rgb <= "000000";
					when "00001000001001111" => rgb <= "000000";
					when "00001000001010000" => rgb <= "000000";
					when "00001000001010001" => rgb <= "000000";
					when "00001000001010010" => rgb <= "000000";
					when "00001000001010011" => rgb <= "000000";
					when "00001000001010100" => rgb <= "000000";
					when "00001000001010101" => rgb <= "000000";
					when "00001000001010110" => rgb <= "000000";
					when "00001000001010111" => rgb <= "000000";
					when "00001000001011000" => rgb <= "000000";
					when "00001000001011001" => rgb <= "000000";
					when "00001000001011010" => rgb <= "000000";
					when "00001000001011011" => rgb <= "000000";
					when "00001000001011100" => rgb <= "000000";
					when "00001000001011101" => rgb <= "000000";
					when "00001000001011110" => rgb <= "000000";
					when "00001000001011111" => rgb <= "000000";
					when "00001000001100000" => rgb <= "000000";
					when "00001000001100001" => rgb <= "000000";
					when "00001000001100010" => rgb <= "000000";
					when "00001000001100011" => rgb <= "000000";
					when "00001000001100100" => rgb <= "000000";
					when "00001000001100101" => rgb <= "000000";
					when "00001000001100110" => rgb <= "000000";
					when "00001000001100111" => rgb <= "000000";
					when "00001000001101000" => rgb <= "000000";
					when "00001000001101001" => rgb <= "000000";
					when "00001000001101010" => rgb <= "000000";
					when "00001000001101011" => rgb <= "000000";
					when "00001000001101100" => rgb <= "000000";
					when "00001000001101101" => rgb <= "000000";
					when "00001000001101110" => rgb <= "000000";
					when "00001000001101111" => rgb <= "000000";
					when "00001000001110000" => rgb <= "000000";
					when "00001000001110001" => rgb <= "000000";
					when "00001000001110010" => rgb <= "000000";
					when "00001000001110011" => rgb <= "000000";
					when "00001000001110100" => rgb <= "000000";
					when "00001000001110101" => rgb <= "000000";
					when "00001000001110110" => rgb <= "000000";
					when "00001000001110111" => rgb <= "000000";
					when "00001000001111000" => rgb <= "000000";
					when "00001000001111001" => rgb <= "000000";
					when "00001000001111010" => rgb <= "000000";
					when "00001000001111011" => rgb <= "000000";
					when "00001000001111100" => rgb <= "000000";
					when "00001000001111101" => rgb <= "000000";
					when "00001000001111110" => rgb <= "000000";
					when "00001000001111111" => rgb <= "000000";
					when "00001000010000000" => rgb <= "000000";
					when "00001000010000001" => rgb <= "000000";
					when "00001000010000010" => rgb <= "000000";
					when "00001000010000011" => rgb <= "000000";
					when "00001000010000100" => rgb <= "000000";
					when "00001000010000101" => rgb <= "000000";
					when "00001000010000110" => rgb <= "000000";
					when "00001000010000111" => rgb <= "000000";
					when "00001000010001000" => rgb <= "000000";
					when "00001000010001001" => rgb <= "000000";
					when "00001000010001010" => rgb <= "000000";
					when "00001000010001011" => rgb <= "000000";
					when "00001000010001100" => rgb <= "000000";
					when "00001000010001101" => rgb <= "000000";
					when "00001000010001110" => rgb <= "000000";
					when "00001000010001111" => rgb <= "000000";
					when "00001000010010000" => rgb <= "000000";
					when "00001000010010001" => rgb <= "000000";
					when "00001000010010010" => rgb <= "000000";
					when "00001000010010011" => rgb <= "000000";
					when "00001000010010100" => rgb <= "000000";
					when "00001000010010101" => rgb <= "000000";
					when "00001000010010110" => rgb <= "000000";
					when "00001000010010111" => rgb <= "000000";
					when "00001000010011000" => rgb <= "000000";
					when "00001000010011001" => rgb <= "000000";
					when "00001000010011010" => rgb <= "000000";
					when "00001000010011011" => rgb <= "000000";
					when "00001000010011100" => rgb <= "000000";
					when "00001000010011101" => rgb <= "000000";
					when "00001000010011110" => rgb <= "000000";
					when "00001000010011111" => rgb <= "000000";
					when "00001000010100000" => rgb <= "000000";
					when "00001000010100001" => rgb <= "000000";
					when "00001000010100010" => rgb <= "000000";
					when "00001000010100011" => rgb <= "000000";
					when "00001000010100100" => rgb <= "000000";
					when "00001000010100101" => rgb <= "000000";
					when "00001000010100110" => rgb <= "000000";
					when "00001000010100111" => rgb <= "000000";
					when "00001000010101000" => rgb <= "000000";
					when "00001000010101001" => rgb <= "000000";
					when "00001000010101010" => rgb <= "000000";
					when "00001000010101011" => rgb <= "000000";
					when "00001000010101100" => rgb <= "000000";
					when "00001000010101101" => rgb <= "000000";
					when "00001000010101110" => rgb <= "000000";
					when "00001000010101111" => rgb <= "000000";
					when "00001000010110000" => rgb <= "000000";
					when "00001000010110001" => rgb <= "000000";
					when "00001000010110010" => rgb <= "000000";
					when "00001000010110011" => rgb <= "000000";
					when "00001000010110100" => rgb <= "000000";
					when "00001000010110101" => rgb <= "000000";
					when "00001000010110110" => rgb <= "000000";
					when "00001000010110111" => rgb <= "000000";
					when "00001000010111000" => rgb <= "000000";
					when "00001000010111001" => rgb <= "000000";
					when "00001000010111010" => rgb <= "000000";
					when "00001000010111011" => rgb <= "000000";
					when "00001000010111100" => rgb <= "000000";
					when "00001000010111101" => rgb <= "000000";
					when "00001000010111110" => rgb <= "000000";
					when "00001000010111111" => rgb <= "000000";
					when "00001000011000000" => rgb <= "000000";
					when "00001000011000001" => rgb <= "000000";
					when "00001000011000010" => rgb <= "000000";
					when "00001000011000011" => rgb <= "000000";
					when "00001000011000100" => rgb <= "000000";
					when "00001000011000101" => rgb <= "000000";
					when "00001000011000110" => rgb <= "000000";
					when "00001000011000111" => rgb <= "000000";
					when "00001000011001000" => rgb <= "000000";
					when "00001000011001001" => rgb <= "000000";
					when "00001000011001010" => rgb <= "000000";
					when "00001000011001011" => rgb <= "000000";
					when "00001000011001100" => rgb <= "000000";
					when "00001000011001101" => rgb <= "000000";
					when "00001000011001110" => rgb <= "000000";
					when "00001000011001111" => rgb <= "000000";
					when "00001000011010000" => rgb <= "000000";
					when "00001000011010001" => rgb <= "000000";
					when "00001000011010010" => rgb <= "000000";
					when "00001000011010011" => rgb <= "000000";
					when "00001000011010100" => rgb <= "000000";
					when "00001000011010101" => rgb <= "000000";
					when "00001000011010110" => rgb <= "000000";
					when "00001000011010111" => rgb <= "000000";
					when "00001000011011000" => rgb <= "000000";
					when "00001000011011001" => rgb <= "000000";
					when "00001000011011010" => rgb <= "000000";
					when "00001000011011011" => rgb <= "000000";
					when "00001000011011100" => rgb <= "000000";
					when "00001000011011101" => rgb <= "000000";
					when "00001000011011110" => rgb <= "000000";
					when "00001000011011111" => rgb <= "000000";
					when "00001000011100000" => rgb <= "000000";
					when "00001000011100001" => rgb <= "000000";
					when "00001000011100010" => rgb <= "000000";
					when "00001000011100011" => rgb <= "000000";
					when "00001000011100100" => rgb <= "000000";
					when "00001000011100101" => rgb <= "000000";
					when "00001000011100110" => rgb <= "000000";
					when "00001000011100111" => rgb <= "000000";
					when "00001000011101000" => rgb <= "000000";
					when "00001000011101001" => rgb <= "000000";
					when "00001000011101010" => rgb <= "000000";
					when "00001000011101011" => rgb <= "000000";
					when "00001000011101100" => rgb <= "000000";
					when "00001000011101101" => rgb <= "000000";
					when "00001000011101110" => rgb <= "000000";
					when "00001000011101111" => rgb <= "000000";
					when "00001000011110000" => rgb <= "000000";
					when "00001000011110001" => rgb <= "000000";
					when "00001000011110010" => rgb <= "000000";
					when "00001000011110011" => rgb <= "000000";
					when "00001000011110100" => rgb <= "000000";
					when "00001000011110101" => rgb <= "000000";
					when "00001000011110110" => rgb <= "000000";
					when "00001000011110111" => rgb <= "000000";
					when "00001000011111000" => rgb <= "000000";
					when "00001000011111001" => rgb <= "000000";
					when "00001000011111010" => rgb <= "000000";
					when "00001000011111011" => rgb <= "000000";
					when "00001000011111100" => rgb <= "000000";
					when "00001000011111101" => rgb <= "000000";
					when "00001000011111110" => rgb <= "000000";
					when "00001000011111111" => rgb <= "000000";
					when "00001000100000000" => rgb <= "000000";
					when "00001000100000001" => rgb <= "000000";
					when "00001000100000010" => rgb <= "000000";
					when "00001000100000011" => rgb <= "000000";
					when "00001000100000100" => rgb <= "000000";
					when "00001000100000101" => rgb <= "000000";
					when "00001000100000110" => rgb <= "000000";
					when "00001000100000111" => rgb <= "000000";
					when "00001000100001000" => rgb <= "000000";
					when "00001000100001001" => rgb <= "000000";
					when "00001000100001010" => rgb <= "000000";
					when "00001000100001011" => rgb <= "000000";
					when "00001000100001100" => rgb <= "000000";
					when "00001000100001101" => rgb <= "000000";
					when "00001000100001110" => rgb <= "000000";
					when "00001000100001111" => rgb <= "000000";
					when "00001000100010000" => rgb <= "000000";
					when "00001000100010001" => rgb <= "000000";
					when "00001000100010010" => rgb <= "000000";
					when "00001000100010011" => rgb <= "000000";
					when "00001000100010100" => rgb <= "000000";
					when "00001000100010101" => rgb <= "000000";
					when "00001000100010110" => rgb <= "000000";
					when "00001000100010111" => rgb <= "000000";
					when "00001000100011000" => rgb <= "000000";
					when "00001000100011001" => rgb <= "000000";
					when "00001000100011010" => rgb <= "000000";
					when "00001000100011011" => rgb <= "000000";
					when "00001000100011100" => rgb <= "000000";
					when "00001000100011101" => rgb <= "000000";
					when "00001000100011110" => rgb <= "000000";
					when "00001000100011111" => rgb <= "000000";
					when "00001000100100000" => rgb <= "000000";
					when "00001000100100001" => rgb <= "000000";
					when "00001000100100010" => rgb <= "000000";
					when "00001000100100011" => rgb <= "000000";
					when "00001000100100100" => rgb <= "000000";
					when "00001000100100101" => rgb <= "000000";
					when "00001000100100110" => rgb <= "000000";
					when "00001000100100111" => rgb <= "000000";
					when "00001000100101000" => rgb <= "000000";
					when "00001000100101001" => rgb <= "000000";
					when "00001000100101010" => rgb <= "000000";
					when "00001000100101011" => rgb <= "000000";
					when "00001000100101100" => rgb <= "000000";
					when "00001000100101101" => rgb <= "000000";
					when "00001000100101110" => rgb <= "000000";
					when "00001000100101111" => rgb <= "000000";
					when "00001000100110000" => rgb <= "000000";
					when "00001000100110001" => rgb <= "000000";
					when "00001000100110010" => rgb <= "000000";
					when "00001000100110011" => rgb <= "000000";
					when "00001000100110100" => rgb <= "000000";
					when "00001000100110101" => rgb <= "000000";
					when "00001000100110110" => rgb <= "000000";
					when "00001000100110111" => rgb <= "000000";
					when "00001000100111000" => rgb <= "000000";
					when "00001000100111001" => rgb <= "000000";
					when "00001000100111010" => rgb <= "000000";
					when "00001000100111011" => rgb <= "000000";
					when "00001000100111100" => rgb <= "000000";
					when "00001000100111101" => rgb <= "000000";
					when "00001000100111110" => rgb <= "000000";
					when "00001000100111111" => rgb <= "000000";
					when "00001001000000000" => rgb <= "000000";
					when "00001001000000001" => rgb <= "000000";
					when "00001001000000010" => rgb <= "000000";
					when "00001001000000011" => rgb <= "000000";
					when "00001001000000100" => rgb <= "000000";
					when "00001001000000101" => rgb <= "000000";
					when "00001001000000110" => rgb <= "000000";
					when "00001001000000111" => rgb <= "000000";
					when "00001001000001000" => rgb <= "000000";
					when "00001001000001001" => rgb <= "000000";
					when "00001001000001010" => rgb <= "000000";
					when "00001001000001011" => rgb <= "000000";
					when "00001001000001100" => rgb <= "000000";
					when "00001001000001101" => rgb <= "000000";
					when "00001001000001110" => rgb <= "000000";
					when "00001001000001111" => rgb <= "000000";
					when "00001001000010000" => rgb <= "000000";
					when "00001001000010001" => rgb <= "000000";
					when "00001001000010010" => rgb <= "000000";
					when "00001001000010011" => rgb <= "000000";
					when "00001001000010100" => rgb <= "000000";
					when "00001001000010101" => rgb <= "000000";
					when "00001001000010110" => rgb <= "000000";
					when "00001001000010111" => rgb <= "000000";
					when "00001001000011000" => rgb <= "000000";
					when "00001001000011001" => rgb <= "000000";
					when "00001001000011010" => rgb <= "000000";
					when "00001001000011011" => rgb <= "000000";
					when "00001001000011100" => rgb <= "000000";
					when "00001001000011101" => rgb <= "000000";
					when "00001001000011110" => rgb <= "000000";
					when "00001001000011111" => rgb <= "000000";
					when "00001001000100000" => rgb <= "000000";
					when "00001001000100001" => rgb <= "000000";
					when "00001001000100010" => rgb <= "000000";
					when "00001001000100011" => rgb <= "000000";
					when "00001001000100100" => rgb <= "000000";
					when "00001001000100101" => rgb <= "000000";
					when "00001001000100110" => rgb <= "000000";
					when "00001001000100111" => rgb <= "000000";
					when "00001001000101000" => rgb <= "000000";
					when "00001001000101001" => rgb <= "000000";
					when "00001001000101010" => rgb <= "000000";
					when "00001001000101011" => rgb <= "000000";
					when "00001001000101100" => rgb <= "000000";
					when "00001001000101101" => rgb <= "000000";
					when "00001001000101110" => rgb <= "000000";
					when "00001001000101111" => rgb <= "000000";
					when "00001001000110000" => rgb <= "000000";
					when "00001001000110001" => rgb <= "000000";
					when "00001001000110010" => rgb <= "000000";
					when "00001001000110011" => rgb <= "000000";
					when "00001001000110100" => rgb <= "000000";
					when "00001001000110101" => rgb <= "000000";
					when "00001001000110110" => rgb <= "000000";
					when "00001001000110111" => rgb <= "000000";
					when "00001001000111000" => rgb <= "000000";
					when "00001001000111001" => rgb <= "000000";
					when "00001001000111010" => rgb <= "000000";
					when "00001001000111011" => rgb <= "000000";
					when "00001001000111100" => rgb <= "000000";
					when "00001001000111101" => rgb <= "000000";
					when "00001001000111110" => rgb <= "000000";
					when "00001001000111111" => rgb <= "000000";
					when "00001001001000000" => rgb <= "000000";
					when "00001001001000001" => rgb <= "000000";
					when "00001001001000010" => rgb <= "000000";
					when "00001001001000011" => rgb <= "000000";
					when "00001001001000100" => rgb <= "000000";
					when "00001001001000101" => rgb <= "000000";
					when "00001001001000110" => rgb <= "000000";
					when "00001001001000111" => rgb <= "000000";
					when "00001001001001000" => rgb <= "000000";
					when "00001001001001001" => rgb <= "000000";
					when "00001001001001010" => rgb <= "000000";
					when "00001001001001011" => rgb <= "000000";
					when "00001001001001100" => rgb <= "000000";
					when "00001001001001101" => rgb <= "000000";
					when "00001001001001110" => rgb <= "000000";
					when "00001001001001111" => rgb <= "000000";
					when "00001001001010000" => rgb <= "000000";
					when "00001001001010001" => rgb <= "000000";
					when "00001001001010010" => rgb <= "000000";
					when "00001001001010011" => rgb <= "000000";
					when "00001001001010100" => rgb <= "000000";
					when "00001001001010101" => rgb <= "000000";
					when "00001001001010110" => rgb <= "000000";
					when "00001001001010111" => rgb <= "000000";
					when "00001001001011000" => rgb <= "000000";
					when "00001001001011001" => rgb <= "000000";
					when "00001001001011010" => rgb <= "000000";
					when "00001001001011011" => rgb <= "000000";
					when "00001001001011100" => rgb <= "000000";
					when "00001001001011101" => rgb <= "000000";
					when "00001001001011110" => rgb <= "000000";
					when "00001001001011111" => rgb <= "000000";
					when "00001001001100000" => rgb <= "000000";
					when "00001001001100001" => rgb <= "000000";
					when "00001001001100010" => rgb <= "000000";
					when "00001001001100011" => rgb <= "000000";
					when "00001001001100100" => rgb <= "000000";
					when "00001001001100101" => rgb <= "000000";
					when "00001001001100110" => rgb <= "000000";
					when "00001001001100111" => rgb <= "000000";
					when "00001001001101000" => rgb <= "000000";
					when "00001001001101001" => rgb <= "000000";
					when "00001001001101010" => rgb <= "000000";
					when "00001001001101011" => rgb <= "000000";
					when "00001001001101100" => rgb <= "000000";
					when "00001001001101101" => rgb <= "000000";
					when "00001001001101110" => rgb <= "000000";
					when "00001001001101111" => rgb <= "000000";
					when "00001001001110000" => rgb <= "000000";
					when "00001001001110001" => rgb <= "000000";
					when "00001001001110010" => rgb <= "000000";
					when "00001001001110011" => rgb <= "000000";
					when "00001001001110100" => rgb <= "000000";
					when "00001001001110101" => rgb <= "000000";
					when "00001001001110110" => rgb <= "000000";
					when "00001001001110111" => rgb <= "000000";
					when "00001001001111000" => rgb <= "000000";
					when "00001001001111001" => rgb <= "000000";
					when "00001001001111010" => rgb <= "000000";
					when "00001001001111011" => rgb <= "000000";
					when "00001001001111100" => rgb <= "000000";
					when "00001001001111101" => rgb <= "000000";
					when "00001001001111110" => rgb <= "000000";
					when "00001001001111111" => rgb <= "000000";
					when "00001001010000000" => rgb <= "000000";
					when "00001001010000001" => rgb <= "000000";
					when "00001001010000010" => rgb <= "000000";
					when "00001001010000011" => rgb <= "000000";
					when "00001001010000100" => rgb <= "000000";
					when "00001001010000101" => rgb <= "000000";
					when "00001001010000110" => rgb <= "000000";
					when "00001001010000111" => rgb <= "000000";
					when "00001001010001000" => rgb <= "000000";
					when "00001001010001001" => rgb <= "000000";
					when "00001001010001010" => rgb <= "000000";
					when "00001001010001011" => rgb <= "000000";
					when "00001001010001100" => rgb <= "000000";
					when "00001001010001101" => rgb <= "000000";
					when "00001001010001110" => rgb <= "000000";
					when "00001001010001111" => rgb <= "000000";
					when "00001001010010000" => rgb <= "000000";
					when "00001001010010001" => rgb <= "000000";
					when "00001001010010010" => rgb <= "000000";
					when "00001001010010011" => rgb <= "000000";
					when "00001001010010100" => rgb <= "000000";
					when "00001001010010101" => rgb <= "000000";
					when "00001001010010110" => rgb <= "000000";
					when "00001001010010111" => rgb <= "000000";
					when "00001001010011000" => rgb <= "000000";
					when "00001001010011001" => rgb <= "000000";
					when "00001001010011010" => rgb <= "000000";
					when "00001001010011011" => rgb <= "000000";
					when "00001001010011100" => rgb <= "000000";
					when "00001001010011101" => rgb <= "000000";
					when "00001001010011110" => rgb <= "000000";
					when "00001001010011111" => rgb <= "000000";
					when "00001001010100000" => rgb <= "000000";
					when "00001001010100001" => rgb <= "000000";
					when "00001001010100010" => rgb <= "000000";
					when "00001001010100011" => rgb <= "000000";
					when "00001001010100100" => rgb <= "000000";
					when "00001001010100101" => rgb <= "000000";
					when "00001001010100110" => rgb <= "000000";
					when "00001001010100111" => rgb <= "000000";
					when "00001001010101000" => rgb <= "000000";
					when "00001001010101001" => rgb <= "000000";
					when "00001001010101010" => rgb <= "000000";
					when "00001001010101011" => rgb <= "000000";
					when "00001001010101100" => rgb <= "000000";
					when "00001001010101101" => rgb <= "000000";
					when "00001001010101110" => rgb <= "000000";
					when "00001001010101111" => rgb <= "000000";
					when "00001001010110000" => rgb <= "000000";
					when "00001001010110001" => rgb <= "000000";
					when "00001001010110010" => rgb <= "000000";
					when "00001001010110011" => rgb <= "000000";
					when "00001001010110100" => rgb <= "000000";
					when "00001001010110101" => rgb <= "000000";
					when "00001001010110110" => rgb <= "000000";
					when "00001001010110111" => rgb <= "000000";
					when "00001001010111000" => rgb <= "000000";
					when "00001001010111001" => rgb <= "000000";
					when "00001001010111010" => rgb <= "000000";
					when "00001001010111011" => rgb <= "000000";
					when "00001001010111100" => rgb <= "000000";
					when "00001001010111101" => rgb <= "000000";
					when "00001001010111110" => rgb <= "000000";
					when "00001001010111111" => rgb <= "000000";
					when "00001001011000000" => rgb <= "000000";
					when "00001001011000001" => rgb <= "000000";
					when "00001001011000010" => rgb <= "000000";
					when "00001001011000011" => rgb <= "000000";
					when "00001001011000100" => rgb <= "000000";
					when "00001001011000101" => rgb <= "000000";
					when "00001001011000110" => rgb <= "000000";
					when "00001001011000111" => rgb <= "000000";
					when "00001001011001000" => rgb <= "000000";
					when "00001001011001001" => rgb <= "000000";
					when "00001001011001010" => rgb <= "000000";
					when "00001001011001011" => rgb <= "000000";
					when "00001001011001100" => rgb <= "000000";
					when "00001001011001101" => rgb <= "000000";
					when "00001001011001110" => rgb <= "000000";
					when "00001001011001111" => rgb <= "000000";
					when "00001001011010000" => rgb <= "000000";
					when "00001001011010001" => rgb <= "000000";
					when "00001001011010010" => rgb <= "000000";
					when "00001001011010011" => rgb <= "000000";
					when "00001001011010100" => rgb <= "000000";
					when "00001001011010101" => rgb <= "000000";
					when "00001001011010110" => rgb <= "000000";
					when "00001001011010111" => rgb <= "000000";
					when "00001001011011000" => rgb <= "000000";
					when "00001001011011001" => rgb <= "000000";
					when "00001001011011010" => rgb <= "000000";
					when "00001001011011011" => rgb <= "000000";
					when "00001001011011100" => rgb <= "000000";
					when "00001001011011101" => rgb <= "000000";
					when "00001001011011110" => rgb <= "000000";
					when "00001001011011111" => rgb <= "000000";
					when "00001001011100000" => rgb <= "000000";
					when "00001001011100001" => rgb <= "000000";
					when "00001001011100010" => rgb <= "000000";
					when "00001001011100011" => rgb <= "000000";
					when "00001001011100100" => rgb <= "000000";
					when "00001001011100101" => rgb <= "000000";
					when "00001001011100110" => rgb <= "000000";
					when "00001001011100111" => rgb <= "000000";
					when "00001001011101000" => rgb <= "000000";
					when "00001001011101001" => rgb <= "000000";
					when "00001001011101010" => rgb <= "000000";
					when "00001001011101011" => rgb <= "000000";
					when "00001001011101100" => rgb <= "000000";
					when "00001001011101101" => rgb <= "000000";
					when "00001001011101110" => rgb <= "000000";
					when "00001001011101111" => rgb <= "000000";
					when "00001001011110000" => rgb <= "000000";
					when "00001001011110001" => rgb <= "000000";
					when "00001001011110010" => rgb <= "000000";
					when "00001001011110011" => rgb <= "000000";
					when "00001001011110100" => rgb <= "000000";
					when "00001001011110101" => rgb <= "000000";
					when "00001001011110110" => rgb <= "000000";
					when "00001001011110111" => rgb <= "000000";
					when "00001001011111000" => rgb <= "000000";
					when "00001001011111001" => rgb <= "000000";
					when "00001001011111010" => rgb <= "000000";
					when "00001001011111011" => rgb <= "000000";
					when "00001001011111100" => rgb <= "000000";
					when "00001001011111101" => rgb <= "000000";
					when "00001001011111110" => rgb <= "000000";
					when "00001001011111111" => rgb <= "000000";
					when "00001001100000000" => rgb <= "000000";
					when "00001001100000001" => rgb <= "000000";
					when "00001001100000010" => rgb <= "000000";
					when "00001001100000011" => rgb <= "000000";
					when "00001001100000100" => rgb <= "000000";
					when "00001001100000101" => rgb <= "000000";
					when "00001001100000110" => rgb <= "000000";
					when "00001001100000111" => rgb <= "000000";
					when "00001001100001000" => rgb <= "000000";
					when "00001001100001001" => rgb <= "000000";
					when "00001001100001010" => rgb <= "000000";
					when "00001001100001011" => rgb <= "000000";
					when "00001001100001100" => rgb <= "000000";
					when "00001001100001101" => rgb <= "000000";
					when "00001001100001110" => rgb <= "000000";
					when "00001001100001111" => rgb <= "000000";
					when "00001001100010000" => rgb <= "000000";
					when "00001001100010001" => rgb <= "000000";
					when "00001001100010010" => rgb <= "000000";
					when "00001001100010011" => rgb <= "000000";
					when "00001001100010100" => rgb <= "000000";
					when "00001001100010101" => rgb <= "000000";
					when "00001001100010110" => rgb <= "000000";
					when "00001001100010111" => rgb <= "000000";
					when "00001001100011000" => rgb <= "000000";
					when "00001001100011001" => rgb <= "000000";
					when "00001001100011010" => rgb <= "000000";
					when "00001001100011011" => rgb <= "000000";
					when "00001001100011100" => rgb <= "000000";
					when "00001001100011101" => rgb <= "000000";
					when "00001001100011110" => rgb <= "000000";
					when "00001001100011111" => rgb <= "000000";
					when "00001001100100000" => rgb <= "000000";
					when "00001001100100001" => rgb <= "000000";
					when "00001001100100010" => rgb <= "000000";
					when "00001001100100011" => rgb <= "000000";
					when "00001001100100100" => rgb <= "000000";
					when "00001001100100101" => rgb <= "000000";
					when "00001001100100110" => rgb <= "000000";
					when "00001001100100111" => rgb <= "000000";
					when "00001001100101000" => rgb <= "000000";
					when "00001001100101001" => rgb <= "000000";
					when "00001001100101010" => rgb <= "000000";
					when "00001001100101011" => rgb <= "000000";
					when "00001001100101100" => rgb <= "000000";
					when "00001001100101101" => rgb <= "000000";
					when "00001001100101110" => rgb <= "000000";
					when "00001001100101111" => rgb <= "000000";
					when "00001001100110000" => rgb <= "000000";
					when "00001001100110001" => rgb <= "000000";
					when "00001001100110010" => rgb <= "000000";
					when "00001001100110011" => rgb <= "000000";
					when "00001001100110100" => rgb <= "000000";
					when "00001001100110101" => rgb <= "000000";
					when "00001001100110110" => rgb <= "000000";
					when "00001001100110111" => rgb <= "000000";
					when "00001001100111000" => rgb <= "000000";
					when "00001001100111001" => rgb <= "000000";
					when "00001001100111010" => rgb <= "000000";
					when "00001001100111011" => rgb <= "000000";
					when "00001001100111100" => rgb <= "000000";
					when "00001001100111101" => rgb <= "000000";
					when "00001001100111110" => rgb <= "000000";
					when "00001001100111111" => rgb <= "000000";
					when "00001010000000000" => rgb <= "000000";
					when "00001010000000001" => rgb <= "000000";
					when "00001010000000010" => rgb <= "000000";
					when "00001010000000011" => rgb <= "000000";
					when "00001010000000100" => rgb <= "000000";
					when "00001010000000101" => rgb <= "000000";
					when "00001010000000110" => rgb <= "000000";
					when "00001010000000111" => rgb <= "000000";
					when "00001010000001000" => rgb <= "000000";
					when "00001010000001001" => rgb <= "000000";
					when "00001010000001010" => rgb <= "000000";
					when "00001010000001011" => rgb <= "000000";
					when "00001010000001100" => rgb <= "000000";
					when "00001010000001101" => rgb <= "000000";
					when "00001010000001110" => rgb <= "000000";
					when "00001010000001111" => rgb <= "000000";
					when "00001010000010000" => rgb <= "000000";
					when "00001010000010001" => rgb <= "000000";
					when "00001010000010010" => rgb <= "000000";
					when "00001010000010011" => rgb <= "000000";
					when "00001010000010100" => rgb <= "000000";
					when "00001010000010101" => rgb <= "000000";
					when "00001010000010110" => rgb <= "000000";
					when "00001010000010111" => rgb <= "000000";
					when "00001010000011000" => rgb <= "000000";
					when "00001010000011001" => rgb <= "000000";
					when "00001010000011010" => rgb <= "000000";
					when "00001010000011011" => rgb <= "000000";
					when "00001010000011100" => rgb <= "000000";
					when "00001010000011101" => rgb <= "000000";
					when "00001010000011110" => rgb <= "000000";
					when "00001010000011111" => rgb <= "000000";
					when "00001010000100000" => rgb <= "000000";
					when "00001010000100001" => rgb <= "000000";
					when "00001010000100010" => rgb <= "000000";
					when "00001010000100011" => rgb <= "000000";
					when "00001010000100100" => rgb <= "000000";
					when "00001010000100101" => rgb <= "000000";
					when "00001010000100110" => rgb <= "000000";
					when "00001010000100111" => rgb <= "000000";
					when "00001010000101000" => rgb <= "000000";
					when "00001010000101001" => rgb <= "000000";
					when "00001010000101010" => rgb <= "000000";
					when "00001010000101011" => rgb <= "000000";
					when "00001010000101100" => rgb <= "000000";
					when "00001010000101101" => rgb <= "000000";
					when "00001010000101110" => rgb <= "000000";
					when "00001010000101111" => rgb <= "000000";
					when "00001010000110000" => rgb <= "000000";
					when "00001010000110001" => rgb <= "000000";
					when "00001010000110010" => rgb <= "000000";
					when "00001010000110011" => rgb <= "000000";
					when "00001010000110100" => rgb <= "000000";
					when "00001010000110101" => rgb <= "000000";
					when "00001010000110110" => rgb <= "000000";
					when "00001010000110111" => rgb <= "000000";
					when "00001010000111000" => rgb <= "000000";
					when "00001010000111001" => rgb <= "000000";
					when "00001010000111010" => rgb <= "000000";
					when "00001010000111011" => rgb <= "000000";
					when "00001010000111100" => rgb <= "000000";
					when "00001010000111101" => rgb <= "000000";
					when "00001010000111110" => rgb <= "000000";
					when "00001010000111111" => rgb <= "000000";
					when "00001010001000000" => rgb <= "000000";
					when "00001010001000001" => rgb <= "000000";
					when "00001010001000010" => rgb <= "000000";
					when "00001010001000011" => rgb <= "000000";
					when "00001010001000100" => rgb <= "000000";
					when "00001010001000101" => rgb <= "000000";
					when "00001010001000110" => rgb <= "000000";
					when "00001010001000111" => rgb <= "000000";
					when "00001010001001000" => rgb <= "000000";
					when "00001010001001001" => rgb <= "000000";
					when "00001010001001010" => rgb <= "000000";
					when "00001010001001011" => rgb <= "000000";
					when "00001010001001100" => rgb <= "000000";
					when "00001010001001101" => rgb <= "000000";
					when "00001010001001110" => rgb <= "000000";
					when "00001010001001111" => rgb <= "000000";
					when "00001010001010000" => rgb <= "000000";
					when "00001010001010001" => rgb <= "000000";
					when "00001010001010010" => rgb <= "000000";
					when "00001010001010011" => rgb <= "000000";
					when "00001010001010100" => rgb <= "000000";
					when "00001010001010101" => rgb <= "000000";
					when "00001010001010110" => rgb <= "000000";
					when "00001010001010111" => rgb <= "000000";
					when "00001010001011000" => rgb <= "000000";
					when "00001010001011001" => rgb <= "000000";
					when "00001010001011010" => rgb <= "000000";
					when "00001010001011011" => rgb <= "000000";
					when "00001010001011100" => rgb <= "000000";
					when "00001010001011101" => rgb <= "000000";
					when "00001010001011110" => rgb <= "000000";
					when "00001010001011111" => rgb <= "000000";
					when "00001010001100000" => rgb <= "000000";
					when "00001010001100001" => rgb <= "000000";
					when "00001010001100010" => rgb <= "000000";
					when "00001010001100011" => rgb <= "000000";
					when "00001010001100100" => rgb <= "000000";
					when "00001010001100101" => rgb <= "000000";
					when "00001010001100110" => rgb <= "000000";
					when "00001010001100111" => rgb <= "000000";
					when "00001010001101000" => rgb <= "000000";
					when "00001010001101001" => rgb <= "000000";
					when "00001010001101010" => rgb <= "000000";
					when "00001010001101011" => rgb <= "000000";
					when "00001010001101100" => rgb <= "000000";
					when "00001010001101101" => rgb <= "000000";
					when "00001010001101110" => rgb <= "000000";
					when "00001010001101111" => rgb <= "000000";
					when "00001010001110000" => rgb <= "000000";
					when "00001010001110001" => rgb <= "000000";
					when "00001010001110010" => rgb <= "000000";
					when "00001010001110011" => rgb <= "000000";
					when "00001010001110100" => rgb <= "000000";
					when "00001010001110101" => rgb <= "000000";
					when "00001010001110110" => rgb <= "000000";
					when "00001010001110111" => rgb <= "000000";
					when "00001010001111000" => rgb <= "000000";
					when "00001010001111001" => rgb <= "000000";
					when "00001010001111010" => rgb <= "000000";
					when "00001010001111011" => rgb <= "000000";
					when "00001010001111100" => rgb <= "000000";
					when "00001010001111101" => rgb <= "000000";
					when "00001010001111110" => rgb <= "000000";
					when "00001010001111111" => rgb <= "000000";
					when "00001010010000000" => rgb <= "000000";
					when "00001010010000001" => rgb <= "000000";
					when "00001010010000010" => rgb <= "000000";
					when "00001010010000011" => rgb <= "000000";
					when "00001010010000100" => rgb <= "000000";
					when "00001010010000101" => rgb <= "000000";
					when "00001010010000110" => rgb <= "000000";
					when "00001010010000111" => rgb <= "000000";
					when "00001010010001000" => rgb <= "000000";
					when "00001010010001001" => rgb <= "000000";
					when "00001010010001010" => rgb <= "000000";
					when "00001010010001011" => rgb <= "000000";
					when "00001010010001100" => rgb <= "000000";
					when "00001010010001101" => rgb <= "000000";
					when "00001010010001110" => rgb <= "000000";
					when "00001010010001111" => rgb <= "000000";
					when "00001010010010000" => rgb <= "000000";
					when "00001010010010001" => rgb <= "000000";
					when "00001010010010010" => rgb <= "000000";
					when "00001010010010011" => rgb <= "000000";
					when "00001010010010100" => rgb <= "000000";
					when "00001010010010101" => rgb <= "000000";
					when "00001010010010110" => rgb <= "000000";
					when "00001010010010111" => rgb <= "000000";
					when "00001010010011000" => rgb <= "000000";
					when "00001010010011001" => rgb <= "000000";
					when "00001010010011010" => rgb <= "000000";
					when "00001010010011011" => rgb <= "000000";
					when "00001010010011100" => rgb <= "000000";
					when "00001010010011101" => rgb <= "000000";
					when "00001010010011110" => rgb <= "000000";
					when "00001010010011111" => rgb <= "000000";
					when "00001010010100000" => rgb <= "000000";
					when "00001010010100001" => rgb <= "000000";
					when "00001010010100010" => rgb <= "000000";
					when "00001010010100011" => rgb <= "000000";
					when "00001010010100100" => rgb <= "000000";
					when "00001010010100101" => rgb <= "000000";
					when "00001010010100110" => rgb <= "000000";
					when "00001010010100111" => rgb <= "000000";
					when "00001010010101000" => rgb <= "000000";
					when "00001010010101001" => rgb <= "000000";
					when "00001010010101010" => rgb <= "000000";
					when "00001010010101011" => rgb <= "000000";
					when "00001010010101100" => rgb <= "000000";
					when "00001010010101101" => rgb <= "000000";
					when "00001010010101110" => rgb <= "000000";
					when "00001010010101111" => rgb <= "000000";
					when "00001010010110000" => rgb <= "000000";
					when "00001010010110001" => rgb <= "000000";
					when "00001010010110010" => rgb <= "000000";
					when "00001010010110011" => rgb <= "000000";
					when "00001010010110100" => rgb <= "000000";
					when "00001010010110101" => rgb <= "000000";
					when "00001010010110110" => rgb <= "000000";
					when "00001010010110111" => rgb <= "000000";
					when "00001010010111000" => rgb <= "000000";
					when "00001010010111001" => rgb <= "000000";
					when "00001010010111010" => rgb <= "000000";
					when "00001010010111011" => rgb <= "000000";
					when "00001010010111100" => rgb <= "000000";
					when "00001010010111101" => rgb <= "000000";
					when "00001010010111110" => rgb <= "000000";
					when "00001010010111111" => rgb <= "000000";
					when "00001010011000000" => rgb <= "000000";
					when "00001010011000001" => rgb <= "000000";
					when "00001010011000010" => rgb <= "000000";
					when "00001010011000011" => rgb <= "000000";
					when "00001010011000100" => rgb <= "000000";
					when "00001010011000101" => rgb <= "000000";
					when "00001010011000110" => rgb <= "000000";
					when "00001010011000111" => rgb <= "000000";
					when "00001010011001000" => rgb <= "000000";
					when "00001010011001001" => rgb <= "000000";
					when "00001010011001010" => rgb <= "000000";
					when "00001010011001011" => rgb <= "000000";
					when "00001010011001100" => rgb <= "000000";
					when "00001010011001101" => rgb <= "000000";
					when "00001010011001110" => rgb <= "000000";
					when "00001010011001111" => rgb <= "000000";
					when "00001010011010000" => rgb <= "000000";
					when "00001010011010001" => rgb <= "000000";
					when "00001010011010010" => rgb <= "000000";
					when "00001010011010011" => rgb <= "000000";
					when "00001010011010100" => rgb <= "000000";
					when "00001010011010101" => rgb <= "000000";
					when "00001010011010110" => rgb <= "000000";
					when "00001010011010111" => rgb <= "000000";
					when "00001010011011000" => rgb <= "000000";
					when "00001010011011001" => rgb <= "000000";
					when "00001010011011010" => rgb <= "000000";
					when "00001010011011011" => rgb <= "000000";
					when "00001010011011100" => rgb <= "000000";
					when "00001010011011101" => rgb <= "000000";
					when "00001010011011110" => rgb <= "000000";
					when "00001010011011111" => rgb <= "000000";
					when "00001010011100000" => rgb <= "000000";
					when "00001010011100001" => rgb <= "000000";
					when "00001010011100010" => rgb <= "000000";
					when "00001010011100011" => rgb <= "000000";
					when "00001010011100100" => rgb <= "000000";
					when "00001010011100101" => rgb <= "000000";
					when "00001010011100110" => rgb <= "000000";
					when "00001010011100111" => rgb <= "000000";
					when "00001010011101000" => rgb <= "000000";
					when "00001010011101001" => rgb <= "000000";
					when "00001010011101010" => rgb <= "000000";
					when "00001010011101011" => rgb <= "000000";
					when "00001010011101100" => rgb <= "000000";
					when "00001010011101101" => rgb <= "000000";
					when "00001010011101110" => rgb <= "000000";
					when "00001010011101111" => rgb <= "000000";
					when "00001010011110000" => rgb <= "000000";
					when "00001010011110001" => rgb <= "000000";
					when "00001010011110010" => rgb <= "000000";
					when "00001010011110011" => rgb <= "000000";
					when "00001010011110100" => rgb <= "000000";
					when "00001010011110101" => rgb <= "000000";
					when "00001010011110110" => rgb <= "000000";
					when "00001010011110111" => rgb <= "000000";
					when "00001010011111000" => rgb <= "000000";
					when "00001010011111001" => rgb <= "000000";
					when "00001010011111010" => rgb <= "000000";
					when "00001010011111011" => rgb <= "000000";
					when "00001010011111100" => rgb <= "000000";
					when "00001010011111101" => rgb <= "000000";
					when "00001010011111110" => rgb <= "000000";
					when "00001010011111111" => rgb <= "000000";
					when "00001010100000000" => rgb <= "000000";
					when "00001010100000001" => rgb <= "000000";
					when "00001010100000010" => rgb <= "000000";
					when "00001010100000011" => rgb <= "000000";
					when "00001010100000100" => rgb <= "000000";
					when "00001010100000101" => rgb <= "000000";
					when "00001010100000110" => rgb <= "000000";
					when "00001010100000111" => rgb <= "000000";
					when "00001010100001000" => rgb <= "000000";
					when "00001010100001001" => rgb <= "000000";
					when "00001010100001010" => rgb <= "000000";
					when "00001010100001011" => rgb <= "000000";
					when "00001010100001100" => rgb <= "000000";
					when "00001010100001101" => rgb <= "000000";
					when "00001010100001110" => rgb <= "000000";
					when "00001010100001111" => rgb <= "000000";
					when "00001010100010000" => rgb <= "000000";
					when "00001010100010001" => rgb <= "000000";
					when "00001010100010010" => rgb <= "000000";
					when "00001010100010011" => rgb <= "000000";
					when "00001010100010100" => rgb <= "000000";
					when "00001010100010101" => rgb <= "000000";
					when "00001010100010110" => rgb <= "000000";
					when "00001010100010111" => rgb <= "000000";
					when "00001010100011000" => rgb <= "000000";
					when "00001010100011001" => rgb <= "000000";
					when "00001010100011010" => rgb <= "000000";
					when "00001010100011011" => rgb <= "000000";
					when "00001010100011100" => rgb <= "000000";
					when "00001010100011101" => rgb <= "000000";
					when "00001010100011110" => rgb <= "000000";
					when "00001010100011111" => rgb <= "000000";
					when "00001010100100000" => rgb <= "000000";
					when "00001010100100001" => rgb <= "000000";
					when "00001010100100010" => rgb <= "000000";
					when "00001010100100011" => rgb <= "000000";
					when "00001010100100100" => rgb <= "000000";
					when "00001010100100101" => rgb <= "000000";
					when "00001010100100110" => rgb <= "000000";
					when "00001010100100111" => rgb <= "000000";
					when "00001010100101000" => rgb <= "000000";
					when "00001010100101001" => rgb <= "000000";
					when "00001010100101010" => rgb <= "000000";
					when "00001010100101011" => rgb <= "000000";
					when "00001010100101100" => rgb <= "000000";
					when "00001010100101101" => rgb <= "000000";
					when "00001010100101110" => rgb <= "000000";
					when "00001010100101111" => rgb <= "000000";
					when "00001010100110000" => rgb <= "000000";
					when "00001010100110001" => rgb <= "000000";
					when "00001010100110010" => rgb <= "000000";
					when "00001010100110011" => rgb <= "000000";
					when "00001010100110100" => rgb <= "000000";
					when "00001010100110101" => rgb <= "000000";
					when "00001010100110110" => rgb <= "000000";
					when "00001010100110111" => rgb <= "000000";
					when "00001010100111000" => rgb <= "000000";
					when "00001010100111001" => rgb <= "000000";
					when "00001010100111010" => rgb <= "000000";
					when "00001010100111011" => rgb <= "000000";
					when "00001010100111100" => rgb <= "000000";
					when "00001010100111101" => rgb <= "000000";
					when "00001010100111110" => rgb <= "000000";
					when "00001010100111111" => rgb <= "000000";
					when "00001011000000000" => rgb <= "000000";
					when "00001011000000001" => rgb <= "000000";
					when "00001011000000010" => rgb <= "000000";
					when "00001011000000011" => rgb <= "000000";
					when "00001011000000100" => rgb <= "000000";
					when "00001011000000101" => rgb <= "000000";
					when "00001011000000110" => rgb <= "000000";
					when "00001011000000111" => rgb <= "000000";
					when "00001011000001000" => rgb <= "000000";
					when "00001011000001001" => rgb <= "000000";
					when "00001011000001010" => rgb <= "000000";
					when "00001011000001011" => rgb <= "000000";
					when "00001011000001100" => rgb <= "000000";
					when "00001011000001101" => rgb <= "000000";
					when "00001011000001110" => rgb <= "000000";
					when "00001011000001111" => rgb <= "000000";
					when "00001011000010000" => rgb <= "000000";
					when "00001011000010001" => rgb <= "000000";
					when "00001011000010010" => rgb <= "000000";
					when "00001011000010011" => rgb <= "000000";
					when "00001011000010100" => rgb <= "000000";
					when "00001011000010101" => rgb <= "000000";
					when "00001011000010110" => rgb <= "000000";
					when "00001011000010111" => rgb <= "000000";
					when "00001011000011000" => rgb <= "000000";
					when "00001011000011001" => rgb <= "000000";
					when "00001011000011010" => rgb <= "000000";
					when "00001011000011011" => rgb <= "000000";
					when "00001011000011100" => rgb <= "000000";
					when "00001011000011101" => rgb <= "000000";
					when "00001011000011110" => rgb <= "000000";
					when "00001011000011111" => rgb <= "000000";
					when "00001011000100000" => rgb <= "000000";
					when "00001011000100001" => rgb <= "000000";
					when "00001011000100010" => rgb <= "000000";
					when "00001011000100011" => rgb <= "000000";
					when "00001011000100100" => rgb <= "000000";
					when "00001011000100101" => rgb <= "000000";
					when "00001011000100110" => rgb <= "000000";
					when "00001011000100111" => rgb <= "000000";
					when "00001011000101000" => rgb <= "000000";
					when "00001011000101001" => rgb <= "000000";
					when "00001011000101010" => rgb <= "000000";
					when "00001011000101011" => rgb <= "000000";
					when "00001011000101100" => rgb <= "000000";
					when "00001011000101101" => rgb <= "000000";
					when "00001011000101110" => rgb <= "000000";
					when "00001011000101111" => rgb <= "000000";
					when "00001011000110000" => rgb <= "000000";
					when "00001011000110001" => rgb <= "000000";
					when "00001011000110010" => rgb <= "000000";
					when "00001011000110011" => rgb <= "000000";
					when "00001011000110100" => rgb <= "000000";
					when "00001011000110101" => rgb <= "000000";
					when "00001011000110110" => rgb <= "000000";
					when "00001011000110111" => rgb <= "000000";
					when "00001011000111000" => rgb <= "000000";
					when "00001011000111001" => rgb <= "000000";
					when "00001011000111010" => rgb <= "000000";
					when "00001011000111011" => rgb <= "000000";
					when "00001011000111100" => rgb <= "000000";
					when "00001011000111101" => rgb <= "000000";
					when "00001011000111110" => rgb <= "000000";
					when "00001011000111111" => rgb <= "000000";
					when "00001011001000000" => rgb <= "000000";
					when "00001011001000001" => rgb <= "000000";
					when "00001011001000010" => rgb <= "000000";
					when "00001011001000011" => rgb <= "000000";
					when "00001011001000100" => rgb <= "000000";
					when "00001011001000101" => rgb <= "000000";
					when "00001011001000110" => rgb <= "000000";
					when "00001011001000111" => rgb <= "000000";
					when "00001011001001000" => rgb <= "000000";
					when "00001011001001001" => rgb <= "000000";
					when "00001011001001010" => rgb <= "000000";
					when "00001011001001011" => rgb <= "000000";
					when "00001011001001100" => rgb <= "000000";
					when "00001011001001101" => rgb <= "000000";
					when "00001011001001110" => rgb <= "000000";
					when "00001011001001111" => rgb <= "000000";
					when "00001011001010000" => rgb <= "000000";
					when "00001011001010001" => rgb <= "000000";
					when "00001011001010010" => rgb <= "000000";
					when "00001011001010011" => rgb <= "000000";
					when "00001011001010100" => rgb <= "000000";
					when "00001011001010101" => rgb <= "000000";
					when "00001011001010110" => rgb <= "000000";
					when "00001011001010111" => rgb <= "000000";
					when "00001011001011000" => rgb <= "000000";
					when "00001011001011001" => rgb <= "000000";
					when "00001011001011010" => rgb <= "000000";
					when "00001011001011011" => rgb <= "000000";
					when "00001011001011100" => rgb <= "000000";
					when "00001011001011101" => rgb <= "000000";
					when "00001011001011110" => rgb <= "000000";
					when "00001011001011111" => rgb <= "000000";
					when "00001011001100000" => rgb <= "000000";
					when "00001011001100001" => rgb <= "000000";
					when "00001011001100010" => rgb <= "000000";
					when "00001011001100011" => rgb <= "000000";
					when "00001011001100100" => rgb <= "000000";
					when "00001011001100101" => rgb <= "000000";
					when "00001011001100110" => rgb <= "000000";
					when "00001011001100111" => rgb <= "000000";
					when "00001011001101000" => rgb <= "000000";
					when "00001011001101001" => rgb <= "000000";
					when "00001011001101010" => rgb <= "000000";
					when "00001011001101011" => rgb <= "000000";
					when "00001011001101100" => rgb <= "000000";
					when "00001011001101101" => rgb <= "000000";
					when "00001011001101110" => rgb <= "000000";
					when "00001011001101111" => rgb <= "000000";
					when "00001011001110000" => rgb <= "000000";
					when "00001011001110001" => rgb <= "000000";
					when "00001011001110010" => rgb <= "000000";
					when "00001011001110011" => rgb <= "000000";
					when "00001011001110100" => rgb <= "000000";
					when "00001011001110101" => rgb <= "000000";
					when "00001011001110110" => rgb <= "000000";
					when "00001011001110111" => rgb <= "000000";
					when "00001011001111000" => rgb <= "000000";
					when "00001011001111001" => rgb <= "000000";
					when "00001011001111010" => rgb <= "000000";
					when "00001011001111011" => rgb <= "000000";
					when "00001011001111100" => rgb <= "000000";
					when "00001011001111101" => rgb <= "000000";
					when "00001011001111110" => rgb <= "000000";
					when "00001011001111111" => rgb <= "000000";
					when "00001011010000000" => rgb <= "000000";
					when "00001011010000001" => rgb <= "000000";
					when "00001011010000010" => rgb <= "000000";
					when "00001011010000011" => rgb <= "000000";
					when "00001011010000100" => rgb <= "000000";
					when "00001011010000101" => rgb <= "000000";
					when "00001011010000110" => rgb <= "000000";
					when "00001011010000111" => rgb <= "000000";
					when "00001011010001000" => rgb <= "000000";
					when "00001011010001001" => rgb <= "000000";
					when "00001011010001010" => rgb <= "000000";
					when "00001011010001011" => rgb <= "000000";
					when "00001011010001100" => rgb <= "000000";
					when "00001011010001101" => rgb <= "000000";
					when "00001011010001110" => rgb <= "000000";
					when "00001011010001111" => rgb <= "000000";
					when "00001011010010000" => rgb <= "000000";
					when "00001011010010001" => rgb <= "000000";
					when "00001011010010010" => rgb <= "000000";
					when "00001011010010011" => rgb <= "000000";
					when "00001011010010100" => rgb <= "000000";
					when "00001011010010101" => rgb <= "000000";
					when "00001011010010110" => rgb <= "000000";
					when "00001011010010111" => rgb <= "000000";
					when "00001011010011000" => rgb <= "000000";
					when "00001011010011001" => rgb <= "000000";
					when "00001011010011010" => rgb <= "000000";
					when "00001011010011011" => rgb <= "000000";
					when "00001011010011100" => rgb <= "000000";
					when "00001011010011101" => rgb <= "000000";
					when "00001011010011110" => rgb <= "000000";
					when "00001011010011111" => rgb <= "000000";
					when "00001011010100000" => rgb <= "000000";
					when "00001011010100001" => rgb <= "000000";
					when "00001011010100010" => rgb <= "000000";
					when "00001011010100011" => rgb <= "000000";
					when "00001011010100100" => rgb <= "000000";
					when "00001011010100101" => rgb <= "000000";
					when "00001011010100110" => rgb <= "000000";
					when "00001011010100111" => rgb <= "000000";
					when "00001011010101000" => rgb <= "000000";
					when "00001011010101001" => rgb <= "000000";
					when "00001011010101010" => rgb <= "000000";
					when "00001011010101011" => rgb <= "000000";
					when "00001011010101100" => rgb <= "000000";
					when "00001011010101101" => rgb <= "000000";
					when "00001011010101110" => rgb <= "000000";
					when "00001011010101111" => rgb <= "000000";
					when "00001011010110000" => rgb <= "000000";
					when "00001011010110001" => rgb <= "000000";
					when "00001011010110010" => rgb <= "000000";
					when "00001011010110011" => rgb <= "000000";
					when "00001011010110100" => rgb <= "000000";
					when "00001011010110101" => rgb <= "000000";
					when "00001011010110110" => rgb <= "000000";
					when "00001011010110111" => rgb <= "000000";
					when "00001011010111000" => rgb <= "000000";
					when "00001011010111001" => rgb <= "000000";
					when "00001011010111010" => rgb <= "000000";
					when "00001011010111011" => rgb <= "000000";
					when "00001011010111100" => rgb <= "000000";
					when "00001011010111101" => rgb <= "000000";
					when "00001011010111110" => rgb <= "000000";
					when "00001011010111111" => rgb <= "000000";
					when "00001011011000000" => rgb <= "000000";
					when "00001011011000001" => rgb <= "000000";
					when "00001011011000010" => rgb <= "000000";
					when "00001011011000011" => rgb <= "000000";
					when "00001011011000100" => rgb <= "000000";
					when "00001011011000101" => rgb <= "000000";
					when "00001011011000110" => rgb <= "000000";
					when "00001011011000111" => rgb <= "000000";
					when "00001011011001000" => rgb <= "000000";
					when "00001011011001001" => rgb <= "000000";
					when "00001011011001010" => rgb <= "000000";
					when "00001011011001011" => rgb <= "000000";
					when "00001011011001100" => rgb <= "000000";
					when "00001011011001101" => rgb <= "000000";
					when "00001011011001110" => rgb <= "000000";
					when "00001011011001111" => rgb <= "000000";
					when "00001011011010000" => rgb <= "000000";
					when "00001011011010001" => rgb <= "000000";
					when "00001011011010010" => rgb <= "000000";
					when "00001011011010011" => rgb <= "000000";
					when "00001011011010100" => rgb <= "000000";
					when "00001011011010101" => rgb <= "000000";
					when "00001011011010110" => rgb <= "000000";
					when "00001011011010111" => rgb <= "000000";
					when "00001011011011000" => rgb <= "000000";
					when "00001011011011001" => rgb <= "000000";
					when "00001011011011010" => rgb <= "000000";
					when "00001011011011011" => rgb <= "000000";
					when "00001011011011100" => rgb <= "000000";
					when "00001011011011101" => rgb <= "000000";
					when "00001011011011110" => rgb <= "000000";
					when "00001011011011111" => rgb <= "000000";
					when "00001011011100000" => rgb <= "000000";
					when "00001011011100001" => rgb <= "000000";
					when "00001011011100010" => rgb <= "000000";
					when "00001011011100011" => rgb <= "000000";
					when "00001011011100100" => rgb <= "000000";
					when "00001011011100101" => rgb <= "000000";
					when "00001011011100110" => rgb <= "000000";
					when "00001011011100111" => rgb <= "000000";
					when "00001011011101000" => rgb <= "000000";
					when "00001011011101001" => rgb <= "000000";
					when "00001011011101010" => rgb <= "000000";
					when "00001011011101011" => rgb <= "000000";
					when "00001011011101100" => rgb <= "000000";
					when "00001011011101101" => rgb <= "000000";
					when "00001011011101110" => rgb <= "000000";
					when "00001011011101111" => rgb <= "000000";
					when "00001011011110000" => rgb <= "000000";
					when "00001011011110001" => rgb <= "000000";
					when "00001011011110010" => rgb <= "000000";
					when "00001011011110011" => rgb <= "000000";
					when "00001011011110100" => rgb <= "000000";
					when "00001011011110101" => rgb <= "000000";
					when "00001011011110110" => rgb <= "000000";
					when "00001011011110111" => rgb <= "000000";
					when "00001011011111000" => rgb <= "000000";
					when "00001011011111001" => rgb <= "000000";
					when "00001011011111010" => rgb <= "000000";
					when "00001011011111011" => rgb <= "000000";
					when "00001011011111100" => rgb <= "000000";
					when "00001011011111101" => rgb <= "000000";
					when "00001011011111110" => rgb <= "000000";
					when "00001011011111111" => rgb <= "000000";
					when "00001011100000000" => rgb <= "000000";
					when "00001011100000001" => rgb <= "000000";
					when "00001011100000010" => rgb <= "000000";
					when "00001011100000011" => rgb <= "000000";
					when "00001011100000100" => rgb <= "000000";
					when "00001011100000101" => rgb <= "000000";
					when "00001011100000110" => rgb <= "000000";
					when "00001011100000111" => rgb <= "000000";
					when "00001011100001000" => rgb <= "000000";
					when "00001011100001001" => rgb <= "000000";
					when "00001011100001010" => rgb <= "000000";
					when "00001011100001011" => rgb <= "000000";
					when "00001011100001100" => rgb <= "000000";
					when "00001011100001101" => rgb <= "000000";
					when "00001011100001110" => rgb <= "000000";
					when "00001011100001111" => rgb <= "000000";
					when "00001011100010000" => rgb <= "000000";
					when "00001011100010001" => rgb <= "000000";
					when "00001011100010010" => rgb <= "000000";
					when "00001011100010011" => rgb <= "000000";
					when "00001011100010100" => rgb <= "000000";
					when "00001011100010101" => rgb <= "000000";
					when "00001011100010110" => rgb <= "000000";
					when "00001011100010111" => rgb <= "000000";
					when "00001011100011000" => rgb <= "000000";
					when "00001011100011001" => rgb <= "000000";
					when "00001011100011010" => rgb <= "000000";
					when "00001011100011011" => rgb <= "000000";
					when "00001011100011100" => rgb <= "000000";
					when "00001011100011101" => rgb <= "000000";
					when "00001011100011110" => rgb <= "000000";
					when "00001011100011111" => rgb <= "000000";
					when "00001011100100000" => rgb <= "000000";
					when "00001011100100001" => rgb <= "000000";
					when "00001011100100010" => rgb <= "000000";
					when "00001011100100011" => rgb <= "000000";
					when "00001011100100100" => rgb <= "000000";
					when "00001011100100101" => rgb <= "000000";
					when "00001011100100110" => rgb <= "000000";
					when "00001011100100111" => rgb <= "000000";
					when "00001011100101000" => rgb <= "000000";
					when "00001011100101001" => rgb <= "000000";
					when "00001011100101010" => rgb <= "000000";
					when "00001011100101011" => rgb <= "000000";
					when "00001011100101100" => rgb <= "000000";
					when "00001011100101101" => rgb <= "000000";
					when "00001011100101110" => rgb <= "000000";
					when "00001011100101111" => rgb <= "000000";
					when "00001011100110000" => rgb <= "000000";
					when "00001011100110001" => rgb <= "000000";
					when "00001011100110010" => rgb <= "000000";
					when "00001011100110011" => rgb <= "000000";
					when "00001011100110100" => rgb <= "000000";
					when "00001011100110101" => rgb <= "000000";
					when "00001011100110110" => rgb <= "000000";
					when "00001011100110111" => rgb <= "000000";
					when "00001011100111000" => rgb <= "000000";
					when "00001011100111001" => rgb <= "000000";
					when "00001011100111010" => rgb <= "000000";
					when "00001011100111011" => rgb <= "000000";
					when "00001011100111100" => rgb <= "000000";
					when "00001011100111101" => rgb <= "000000";
					when "00001011100111110" => rgb <= "000000";
					when "00001011100111111" => rgb <= "000000";
					when "00001100000000000" => rgb <= "000000";
					when "00001100000000001" => rgb <= "000000";
					when "00001100000000010" => rgb <= "000000";
					when "00001100000000011" => rgb <= "000000";
					when "00001100000000100" => rgb <= "000000";
					when "00001100000000101" => rgb <= "000000";
					when "00001100000000110" => rgb <= "000000";
					when "00001100000000111" => rgb <= "000000";
					when "00001100000001000" => rgb <= "000000";
					when "00001100000001001" => rgb <= "000000";
					when "00001100000001010" => rgb <= "000000";
					when "00001100000001011" => rgb <= "000000";
					when "00001100000001100" => rgb <= "000000";
					when "00001100000001101" => rgb <= "000000";
					when "00001100000001110" => rgb <= "000000";
					when "00001100000001111" => rgb <= "000000";
					when "00001100000010000" => rgb <= "000000";
					when "00001100000010001" => rgb <= "000000";
					when "00001100000010010" => rgb <= "000000";
					when "00001100000010011" => rgb <= "000000";
					when "00001100000010100" => rgb <= "000000";
					when "00001100000010101" => rgb <= "000000";
					when "00001100000010110" => rgb <= "000000";
					when "00001100000010111" => rgb <= "000000";
					when "00001100000011000" => rgb <= "000000";
					when "00001100000011001" => rgb <= "000000";
					when "00001100000011010" => rgb <= "000000";
					when "00001100000011011" => rgb <= "000000";
					when "00001100000011100" => rgb <= "000000";
					when "00001100000011101" => rgb <= "000000";
					when "00001100000011110" => rgb <= "000000";
					when "00001100000011111" => rgb <= "000000";
					when "00001100000100000" => rgb <= "000000";
					when "00001100000100001" => rgb <= "000000";
					when "00001100000100010" => rgb <= "000000";
					when "00001100000100011" => rgb <= "000000";
					when "00001100000100100" => rgb <= "000000";
					when "00001100000100101" => rgb <= "000000";
					when "00001100000100110" => rgb <= "000000";
					when "00001100000100111" => rgb <= "000000";
					when "00001100000101000" => rgb <= "000000";
					when "00001100000101001" => rgb <= "000000";
					when "00001100000101010" => rgb <= "000000";
					when "00001100000101011" => rgb <= "000000";
					when "00001100000101100" => rgb <= "000000";
					when "00001100000101101" => rgb <= "000000";
					when "00001100000101110" => rgb <= "000000";
					when "00001100000101111" => rgb <= "000000";
					when "00001100000110000" => rgb <= "000000";
					when "00001100000110001" => rgb <= "000000";
					when "00001100000110010" => rgb <= "000000";
					when "00001100000110011" => rgb <= "000000";
					when "00001100000110100" => rgb <= "000000";
					when "00001100000110101" => rgb <= "000000";
					when "00001100000110110" => rgb <= "000000";
					when "00001100000110111" => rgb <= "000000";
					when "00001100000111000" => rgb <= "000000";
					when "00001100000111001" => rgb <= "000000";
					when "00001100000111010" => rgb <= "000000";
					when "00001100000111011" => rgb <= "000000";
					when "00001100000111100" => rgb <= "000000";
					when "00001100000111101" => rgb <= "000000";
					when "00001100000111110" => rgb <= "000000";
					when "00001100000111111" => rgb <= "000000";
					when "00001100001000000" => rgb <= "000000";
					when "00001100001000001" => rgb <= "000000";
					when "00001100001000010" => rgb <= "000000";
					when "00001100001000011" => rgb <= "000000";
					when "00001100001000100" => rgb <= "000000";
					when "00001100001000101" => rgb <= "000000";
					when "00001100001000110" => rgb <= "000000";
					when "00001100001000111" => rgb <= "000000";
					when "00001100001001000" => rgb <= "000000";
					when "00001100001001001" => rgb <= "000000";
					when "00001100001001010" => rgb <= "000000";
					when "00001100001001011" => rgb <= "000000";
					when "00001100001001100" => rgb <= "000000";
					when "00001100001001101" => rgb <= "000000";
					when "00001100001001110" => rgb <= "000000";
					when "00001100001001111" => rgb <= "000000";
					when "00001100001010000" => rgb <= "000000";
					when "00001100001010001" => rgb <= "000000";
					when "00001100001010010" => rgb <= "000000";
					when "00001100001010011" => rgb <= "000000";
					when "00001100001010100" => rgb <= "000000";
					when "00001100001010101" => rgb <= "000000";
					when "00001100001010110" => rgb <= "000000";
					when "00001100001010111" => rgb <= "000000";
					when "00001100001011000" => rgb <= "000000";
					when "00001100001011001" => rgb <= "000000";
					when "00001100001011010" => rgb <= "000000";
					when "00001100001011011" => rgb <= "000000";
					when "00001100001011100" => rgb <= "000000";
					when "00001100001011101" => rgb <= "000000";
					when "00001100001011110" => rgb <= "000000";
					when "00001100001011111" => rgb <= "000000";
					when "00001100001100000" => rgb <= "000000";
					when "00001100001100001" => rgb <= "000000";
					when "00001100001100010" => rgb <= "000000";
					when "00001100001100011" => rgb <= "000000";
					when "00001100001100100" => rgb <= "000000";
					when "00001100001100101" => rgb <= "000000";
					when "00001100001100110" => rgb <= "000000";
					when "00001100001100111" => rgb <= "000000";
					when "00001100001101000" => rgb <= "000000";
					when "00001100001101001" => rgb <= "000000";
					when "00001100001101010" => rgb <= "000000";
					when "00001100001101011" => rgb <= "000000";
					when "00001100001101100" => rgb <= "000000";
					when "00001100001101101" => rgb <= "000000";
					when "00001100001101110" => rgb <= "000000";
					when "00001100001101111" => rgb <= "000000";
					when "00001100001110000" => rgb <= "000000";
					when "00001100001110001" => rgb <= "000000";
					when "00001100001110010" => rgb <= "000000";
					when "00001100001110011" => rgb <= "000000";
					when "00001100001110100" => rgb <= "000000";
					when "00001100001110101" => rgb <= "000000";
					when "00001100001110110" => rgb <= "000000";
					when "00001100001110111" => rgb <= "000000";
					when "00001100001111000" => rgb <= "000000";
					when "00001100001111001" => rgb <= "000000";
					when "00001100001111010" => rgb <= "000000";
					when "00001100001111011" => rgb <= "000000";
					when "00001100001111100" => rgb <= "000000";
					when "00001100001111101" => rgb <= "000000";
					when "00001100001111110" => rgb <= "000000";
					when "00001100001111111" => rgb <= "000000";
					when "00001100010000000" => rgb <= "000000";
					when "00001100010000001" => rgb <= "000000";
					when "00001100010000010" => rgb <= "000000";
					when "00001100010000011" => rgb <= "000000";
					when "00001100010000100" => rgb <= "000000";
					when "00001100010000101" => rgb <= "000000";
					when "00001100010000110" => rgb <= "000000";
					when "00001100010000111" => rgb <= "000000";
					when "00001100010001000" => rgb <= "000000";
					when "00001100010001001" => rgb <= "000000";
					when "00001100010001010" => rgb <= "000000";
					when "00001100010001011" => rgb <= "000000";
					when "00001100010001100" => rgb <= "000000";
					when "00001100010001101" => rgb <= "000000";
					when "00001100010001110" => rgb <= "000000";
					when "00001100010001111" => rgb <= "000000";
					when "00001100010010000" => rgb <= "000000";
					when "00001100010010001" => rgb <= "000000";
					when "00001100010010010" => rgb <= "000000";
					when "00001100010010011" => rgb <= "000000";
					when "00001100010010100" => rgb <= "000000";
					when "00001100010010101" => rgb <= "000000";
					when "00001100010010110" => rgb <= "000000";
					when "00001100010010111" => rgb <= "000000";
					when "00001100010011000" => rgb <= "000000";
					when "00001100010011001" => rgb <= "000000";
					when "00001100010011010" => rgb <= "000000";
					when "00001100010011011" => rgb <= "000000";
					when "00001100010011100" => rgb <= "000000";
					when "00001100010011101" => rgb <= "000000";
					when "00001100010011110" => rgb <= "000000";
					when "00001100010011111" => rgb <= "000000";
					when "00001100010100000" => rgb <= "000000";
					when "00001100010100001" => rgb <= "000000";
					when "00001100010100010" => rgb <= "000000";
					when "00001100010100011" => rgb <= "000000";
					when "00001100010100100" => rgb <= "000000";
					when "00001100010100101" => rgb <= "000000";
					when "00001100010100110" => rgb <= "000000";
					when "00001100010100111" => rgb <= "000000";
					when "00001100010101000" => rgb <= "000000";
					when "00001100010101001" => rgb <= "000000";
					when "00001100010101010" => rgb <= "000000";
					when "00001100010101011" => rgb <= "000000";
					when "00001100010101100" => rgb <= "000000";
					when "00001100010101101" => rgb <= "000000";
					when "00001100010101110" => rgb <= "000000";
					when "00001100010101111" => rgb <= "000000";
					when "00001100010110000" => rgb <= "000000";
					when "00001100010110001" => rgb <= "000000";
					when "00001100010110010" => rgb <= "000000";
					when "00001100010110011" => rgb <= "000000";
					when "00001100010110100" => rgb <= "000000";
					when "00001100010110101" => rgb <= "000000";
					when "00001100010110110" => rgb <= "000000";
					when "00001100010110111" => rgb <= "000000";
					when "00001100010111000" => rgb <= "000000";
					when "00001100010111001" => rgb <= "000000";
					when "00001100010111010" => rgb <= "000000";
					when "00001100010111011" => rgb <= "000000";
					when "00001100010111100" => rgb <= "000000";
					when "00001100010111101" => rgb <= "000000";
					when "00001100010111110" => rgb <= "000000";
					when "00001100010111111" => rgb <= "000000";
					when "00001100011000000" => rgb <= "000000";
					when "00001100011000001" => rgb <= "000000";
					when "00001100011000010" => rgb <= "000000";
					when "00001100011000011" => rgb <= "000000";
					when "00001100011000100" => rgb <= "000000";
					when "00001100011000101" => rgb <= "000000";
					when "00001100011000110" => rgb <= "000000";
					when "00001100011000111" => rgb <= "000000";
					when "00001100011001000" => rgb <= "000000";
					when "00001100011001001" => rgb <= "000000";
					when "00001100011001010" => rgb <= "000000";
					when "00001100011001011" => rgb <= "000000";
					when "00001100011001100" => rgb <= "000000";
					when "00001100011001101" => rgb <= "000000";
					when "00001100011001110" => rgb <= "000000";
					when "00001100011001111" => rgb <= "000000";
					when "00001100011010000" => rgb <= "000000";
					when "00001100011010001" => rgb <= "000000";
					when "00001100011010010" => rgb <= "000000";
					when "00001100011010011" => rgb <= "000000";
					when "00001100011010100" => rgb <= "000000";
					when "00001100011010101" => rgb <= "000000";
					when "00001100011010110" => rgb <= "000000";
					when "00001100011010111" => rgb <= "000000";
					when "00001100011011000" => rgb <= "000000";
					when "00001100011011001" => rgb <= "000000";
					when "00001100011011010" => rgb <= "000000";
					when "00001100011011011" => rgb <= "000000";
					when "00001100011011100" => rgb <= "000000";
					when "00001100011011101" => rgb <= "000000";
					when "00001100011011110" => rgb <= "000000";
					when "00001100011011111" => rgb <= "000000";
					when "00001100011100000" => rgb <= "000000";
					when "00001100011100001" => rgb <= "000000";
					when "00001100011100010" => rgb <= "000000";
					when "00001100011100011" => rgb <= "000000";
					when "00001100011100100" => rgb <= "000000";
					when "00001100011100101" => rgb <= "000000";
					when "00001100011100110" => rgb <= "000000";
					when "00001100011100111" => rgb <= "000000";
					when "00001100011101000" => rgb <= "000000";
					when "00001100011101001" => rgb <= "000000";
					when "00001100011101010" => rgb <= "000000";
					when "00001100011101011" => rgb <= "000000";
					when "00001100011101100" => rgb <= "000000";
					when "00001100011101101" => rgb <= "000000";
					when "00001100011101110" => rgb <= "000000";
					when "00001100011101111" => rgb <= "000000";
					when "00001100011110000" => rgb <= "000000";
					when "00001100011110001" => rgb <= "000000";
					when "00001100011110010" => rgb <= "000000";
					when "00001100011110011" => rgb <= "000000";
					when "00001100011110100" => rgb <= "000000";
					when "00001100011110101" => rgb <= "000000";
					when "00001100011110110" => rgb <= "000000";
					when "00001100011110111" => rgb <= "000000";
					when "00001100011111000" => rgb <= "000000";
					when "00001100011111001" => rgb <= "000000";
					when "00001100011111010" => rgb <= "000000";
					when "00001100011111011" => rgb <= "000000";
					when "00001100011111100" => rgb <= "000000";
					when "00001100011111101" => rgb <= "000000";
					when "00001100011111110" => rgb <= "000000";
					when "00001100011111111" => rgb <= "000000";
					when "00001100100000000" => rgb <= "000000";
					when "00001100100000001" => rgb <= "000000";
					when "00001100100000010" => rgb <= "000000";
					when "00001100100000011" => rgb <= "000000";
					when "00001100100000100" => rgb <= "000000";
					when "00001100100000101" => rgb <= "000000";
					when "00001100100000110" => rgb <= "000000";
					when "00001100100000111" => rgb <= "000000";
					when "00001100100001000" => rgb <= "000000";
					when "00001100100001001" => rgb <= "000000";
					when "00001100100001010" => rgb <= "000000";
					when "00001100100001011" => rgb <= "000000";
					when "00001100100001100" => rgb <= "000000";
					when "00001100100001101" => rgb <= "000000";
					when "00001100100001110" => rgb <= "000000";
					when "00001100100001111" => rgb <= "000000";
					when "00001100100010000" => rgb <= "000000";
					when "00001100100010001" => rgb <= "000000";
					when "00001100100010010" => rgb <= "000000";
					when "00001100100010011" => rgb <= "000000";
					when "00001100100010100" => rgb <= "000000";
					when "00001100100010101" => rgb <= "000000";
					when "00001100100010110" => rgb <= "000000";
					when "00001100100010111" => rgb <= "000000";
					when "00001100100011000" => rgb <= "000000";
					when "00001100100011001" => rgb <= "000000";
					when "00001100100011010" => rgb <= "000000";
					when "00001100100011011" => rgb <= "000000";
					when "00001100100011100" => rgb <= "000000";
					when "00001100100011101" => rgb <= "000000";
					when "00001100100011110" => rgb <= "000000";
					when "00001100100011111" => rgb <= "000000";
					when "00001100100100000" => rgb <= "000000";
					when "00001100100100001" => rgb <= "000000";
					when "00001100100100010" => rgb <= "000000";
					when "00001100100100011" => rgb <= "000000";
					when "00001100100100100" => rgb <= "000000";
					when "00001100100100101" => rgb <= "000000";
					when "00001100100100110" => rgb <= "000000";
					when "00001100100100111" => rgb <= "000000";
					when "00001100100101000" => rgb <= "000000";
					when "00001100100101001" => rgb <= "000000";
					when "00001100100101010" => rgb <= "000000";
					when "00001100100101011" => rgb <= "000000";
					when "00001100100101100" => rgb <= "000000";
					when "00001100100101101" => rgb <= "000000";
					when "00001100100101110" => rgb <= "000000";
					when "00001100100101111" => rgb <= "000000";
					when "00001100100110000" => rgb <= "000000";
					when "00001100100110001" => rgb <= "000000";
					when "00001100100110010" => rgb <= "000000";
					when "00001100100110011" => rgb <= "000000";
					when "00001100100110100" => rgb <= "000000";
					when "00001100100110101" => rgb <= "000000";
					when "00001100100110110" => rgb <= "000000";
					when "00001100100110111" => rgb <= "000000";
					when "00001100100111000" => rgb <= "000000";
					when "00001100100111001" => rgb <= "000000";
					when "00001100100111010" => rgb <= "000000";
					when "00001100100111011" => rgb <= "000000";
					when "00001100100111100" => rgb <= "000000";
					when "00001100100111101" => rgb <= "000000";
					when "00001100100111110" => rgb <= "000000";
					when "00001100100111111" => rgb <= "000000";
					when "00001101000000000" => rgb <= "000000";
					when "00001101000000001" => rgb <= "000000";
					when "00001101000000010" => rgb <= "000000";
					when "00001101000000011" => rgb <= "000000";
					when "00001101000000100" => rgb <= "000000";
					when "00001101000000101" => rgb <= "000000";
					when "00001101000000110" => rgb <= "000000";
					when "00001101000000111" => rgb <= "000000";
					when "00001101000001000" => rgb <= "000000";
					when "00001101000001001" => rgb <= "000000";
					when "00001101000001010" => rgb <= "000000";
					when "00001101000001011" => rgb <= "000000";
					when "00001101000001100" => rgb <= "000000";
					when "00001101000001101" => rgb <= "000000";
					when "00001101000001110" => rgb <= "000000";
					when "00001101000001111" => rgb <= "000000";
					when "00001101000010000" => rgb <= "000000";
					when "00001101000010001" => rgb <= "000000";
					when "00001101000010010" => rgb <= "000000";
					when "00001101000010011" => rgb <= "000000";
					when "00001101000010100" => rgb <= "000000";
					when "00001101000010101" => rgb <= "000000";
					when "00001101000010110" => rgb <= "000000";
					when "00001101000010111" => rgb <= "000000";
					when "00001101000011000" => rgb <= "000000";
					when "00001101000011001" => rgb <= "000000";
					when "00001101000011010" => rgb <= "000000";
					when "00001101000011011" => rgb <= "000000";
					when "00001101000011100" => rgb <= "000000";
					when "00001101000011101" => rgb <= "000000";
					when "00001101000011110" => rgb <= "000000";
					when "00001101000011111" => rgb <= "000000";
					when "00001101000100000" => rgb <= "000000";
					when "00001101000100001" => rgb <= "000000";
					when "00001101000100010" => rgb <= "000000";
					when "00001101000100011" => rgb <= "000000";
					when "00001101000100100" => rgb <= "000000";
					when "00001101000100101" => rgb <= "000000";
					when "00001101000100110" => rgb <= "000000";
					when "00001101000100111" => rgb <= "000000";
					when "00001101000101000" => rgb <= "000000";
					when "00001101000101001" => rgb <= "000000";
					when "00001101000101010" => rgb <= "000000";
					when "00001101000101011" => rgb <= "000000";
					when "00001101000101100" => rgb <= "000000";
					when "00001101000101101" => rgb <= "000000";
					when "00001101000101110" => rgb <= "000000";
					when "00001101000101111" => rgb <= "000000";
					when "00001101000110000" => rgb <= "000000";
					when "00001101000110001" => rgb <= "000000";
					when "00001101000110010" => rgb <= "000000";
					when "00001101000110011" => rgb <= "000000";
					when "00001101000110100" => rgb <= "000000";
					when "00001101000110101" => rgb <= "000000";
					when "00001101000110110" => rgb <= "000000";
					when "00001101000110111" => rgb <= "000000";
					when "00001101000111000" => rgb <= "000000";
					when "00001101000111001" => rgb <= "000000";
					when "00001101000111010" => rgb <= "000000";
					when "00001101000111011" => rgb <= "000000";
					when "00001101000111100" => rgb <= "000000";
					when "00001101000111101" => rgb <= "000000";
					when "00001101000111110" => rgb <= "000000";
					when "00001101000111111" => rgb <= "000000";
					when "00001101001000000" => rgb <= "000000";
					when "00001101001000001" => rgb <= "000000";
					when "00001101001000010" => rgb <= "000000";
					when "00001101001000011" => rgb <= "000000";
					when "00001101001000100" => rgb <= "000000";
					when "00001101001000101" => rgb <= "000000";
					when "00001101001000110" => rgb <= "000000";
					when "00001101001000111" => rgb <= "000000";
					when "00001101001001000" => rgb <= "000000";
					when "00001101001001001" => rgb <= "000000";
					when "00001101001001010" => rgb <= "000000";
					when "00001101001001011" => rgb <= "000000";
					when "00001101001001100" => rgb <= "000000";
					when "00001101001001101" => rgb <= "000000";
					when "00001101001001110" => rgb <= "000000";
					when "00001101001001111" => rgb <= "000000";
					when "00001101001010000" => rgb <= "000000";
					when "00001101001010001" => rgb <= "000000";
					when "00001101001010010" => rgb <= "000000";
					when "00001101001010011" => rgb <= "000000";
					when "00001101001010100" => rgb <= "000000";
					when "00001101001010101" => rgb <= "000000";
					when "00001101001010110" => rgb <= "000000";
					when "00001101001010111" => rgb <= "000000";
					when "00001101001011000" => rgb <= "000000";
					when "00001101001011001" => rgb <= "000000";
					when "00001101001011010" => rgb <= "000000";
					when "00001101001011011" => rgb <= "000000";
					when "00001101001011100" => rgb <= "000000";
					when "00001101001011101" => rgb <= "000000";
					when "00001101001011110" => rgb <= "000000";
					when "00001101001011111" => rgb <= "000000";
					when "00001101001100000" => rgb <= "000000";
					when "00001101001100001" => rgb <= "000000";
					when "00001101001100010" => rgb <= "000000";
					when "00001101001100011" => rgb <= "000000";
					when "00001101001100100" => rgb <= "000000";
					when "00001101001100101" => rgb <= "000000";
					when "00001101001100110" => rgb <= "000000";
					when "00001101001100111" => rgb <= "000000";
					when "00001101001101000" => rgb <= "000000";
					when "00001101001101001" => rgb <= "000000";
					when "00001101001101010" => rgb <= "000000";
					when "00001101001101011" => rgb <= "000000";
					when "00001101001101100" => rgb <= "000000";
					when "00001101001101101" => rgb <= "000000";
					when "00001101001101110" => rgb <= "000000";
					when "00001101001101111" => rgb <= "000000";
					when "00001101001110000" => rgb <= "000000";
					when "00001101001110001" => rgb <= "000000";
					when "00001101001110010" => rgb <= "000000";
					when "00001101001110011" => rgb <= "000000";
					when "00001101001110100" => rgb <= "000000";
					when "00001101001110101" => rgb <= "000000";
					when "00001101001110110" => rgb <= "000000";
					when "00001101001110111" => rgb <= "000000";
					when "00001101001111000" => rgb <= "000000";
					when "00001101001111001" => rgb <= "000000";
					when "00001101001111010" => rgb <= "000000";
					when "00001101001111011" => rgb <= "000000";
					when "00001101001111100" => rgb <= "000000";
					when "00001101001111101" => rgb <= "000000";
					when "00001101001111110" => rgb <= "000000";
					when "00001101001111111" => rgb <= "000000";
					when "00001101010000000" => rgb <= "000000";
					when "00001101010000001" => rgb <= "000000";
					when "00001101010000010" => rgb <= "000000";
					when "00001101010000011" => rgb <= "000000";
					when "00001101010000100" => rgb <= "000000";
					when "00001101010000101" => rgb <= "000000";
					when "00001101010000110" => rgb <= "000000";
					when "00001101010000111" => rgb <= "000000";
					when "00001101010001000" => rgb <= "000000";
					when "00001101010001001" => rgb <= "000000";
					when "00001101010001010" => rgb <= "000000";
					when "00001101010001011" => rgb <= "000000";
					when "00001101010001100" => rgb <= "000000";
					when "00001101010001101" => rgb <= "000000";
					when "00001101010001110" => rgb <= "000000";
					when "00001101010001111" => rgb <= "000000";
					when "00001101010010000" => rgb <= "000000";
					when "00001101010010001" => rgb <= "000000";
					when "00001101010010010" => rgb <= "000000";
					when "00001101010010011" => rgb <= "000000";
					when "00001101010010100" => rgb <= "000000";
					when "00001101010010101" => rgb <= "000000";
					when "00001101010010110" => rgb <= "000000";
					when "00001101010010111" => rgb <= "000000";
					when "00001101010011000" => rgb <= "000000";
					when "00001101010011001" => rgb <= "000000";
					when "00001101010011010" => rgb <= "000000";
					when "00001101010011011" => rgb <= "000000";
					when "00001101010011100" => rgb <= "000000";
					when "00001101010011101" => rgb <= "000000";
					when "00001101010011110" => rgb <= "000000";
					when "00001101010011111" => rgb <= "000000";
					when "00001101010100000" => rgb <= "000000";
					when "00001101010100001" => rgb <= "000000";
					when "00001101010100010" => rgb <= "000000";
					when "00001101010100011" => rgb <= "000000";
					when "00001101010100100" => rgb <= "000000";
					when "00001101010100101" => rgb <= "000000";
					when "00001101010100110" => rgb <= "000000";
					when "00001101010100111" => rgb <= "000000";
					when "00001101010101000" => rgb <= "000000";
					when "00001101010101001" => rgb <= "000000";
					when "00001101010101010" => rgb <= "000000";
					when "00001101010101011" => rgb <= "000000";
					when "00001101010101100" => rgb <= "000000";
					when "00001101010101101" => rgb <= "000000";
					when "00001101010101110" => rgb <= "000000";
					when "00001101010101111" => rgb <= "000000";
					when "00001101010110000" => rgb <= "000000";
					when "00001101010110001" => rgb <= "000000";
					when "00001101010110010" => rgb <= "000000";
					when "00001101010110011" => rgb <= "000000";
					when "00001101010110100" => rgb <= "000000";
					when "00001101010110101" => rgb <= "000000";
					when "00001101010110110" => rgb <= "000000";
					when "00001101010110111" => rgb <= "000000";
					when "00001101010111000" => rgb <= "000000";
					when "00001101010111001" => rgb <= "000000";
					when "00001101010111010" => rgb <= "000000";
					when "00001101010111011" => rgb <= "000000";
					when "00001101010111100" => rgb <= "000000";
					when "00001101010111101" => rgb <= "000000";
					when "00001101010111110" => rgb <= "000000";
					when "00001101010111111" => rgb <= "000000";
					when "00001101011000000" => rgb <= "000000";
					when "00001101011000001" => rgb <= "000000";
					when "00001101011000010" => rgb <= "000000";
					when "00001101011000011" => rgb <= "000000";
					when "00001101011000100" => rgb <= "000000";
					when "00001101011000101" => rgb <= "000000";
					when "00001101011000110" => rgb <= "000000";
					when "00001101011000111" => rgb <= "000000";
					when "00001101011001000" => rgb <= "000000";
					when "00001101011001001" => rgb <= "000000";
					when "00001101011001010" => rgb <= "000000";
					when "00001101011001011" => rgb <= "000000";
					when "00001101011001100" => rgb <= "000000";
					when "00001101011001101" => rgb <= "000000";
					when "00001101011001110" => rgb <= "000000";
					when "00001101011001111" => rgb <= "000000";
					when "00001101011010000" => rgb <= "000000";
					when "00001101011010001" => rgb <= "000000";
					when "00001101011010010" => rgb <= "000000";
					when "00001101011010011" => rgb <= "000000";
					when "00001101011010100" => rgb <= "000000";
					when "00001101011010101" => rgb <= "000000";
					when "00001101011010110" => rgb <= "000000";
					when "00001101011010111" => rgb <= "000000";
					when "00001101011011000" => rgb <= "000000";
					when "00001101011011001" => rgb <= "000000";
					when "00001101011011010" => rgb <= "000000";
					when "00001101011011011" => rgb <= "000000";
					when "00001101011011100" => rgb <= "000000";
					when "00001101011011101" => rgb <= "000000";
					when "00001101011011110" => rgb <= "000000";
					when "00001101011011111" => rgb <= "000000";
					when "00001101011100000" => rgb <= "000000";
					when "00001101011100001" => rgb <= "000000";
					when "00001101011100010" => rgb <= "000000";
					when "00001101011100011" => rgb <= "000000";
					when "00001101011100100" => rgb <= "000000";
					when "00001101011100101" => rgb <= "000000";
					when "00001101011100110" => rgb <= "000000";
					when "00001101011100111" => rgb <= "000000";
					when "00001101011101000" => rgb <= "000000";
					when "00001101011101001" => rgb <= "000000";
					when "00001101011101010" => rgb <= "000000";
					when "00001101011101011" => rgb <= "000000";
					when "00001101011101100" => rgb <= "000000";
					when "00001101011101101" => rgb <= "000000";
					when "00001101011101110" => rgb <= "000000";
					when "00001101011101111" => rgb <= "000000";
					when "00001101011110000" => rgb <= "000000";
					when "00001101011110001" => rgb <= "000000";
					when "00001101011110010" => rgb <= "000000";
					when "00001101011110011" => rgb <= "000000";
					when "00001101011110100" => rgb <= "000000";
					when "00001101011110101" => rgb <= "000000";
					when "00001101011110110" => rgb <= "000000";
					when "00001101011110111" => rgb <= "000000";
					when "00001101011111000" => rgb <= "000000";
					when "00001101011111001" => rgb <= "000000";
					when "00001101011111010" => rgb <= "000000";
					when "00001101011111011" => rgb <= "000000";
					when "00001101011111100" => rgb <= "000000";
					when "00001101011111101" => rgb <= "000000";
					when "00001101011111110" => rgb <= "000000";
					when "00001101011111111" => rgb <= "000000";
					when "00001101100000000" => rgb <= "000000";
					when "00001101100000001" => rgb <= "000000";
					when "00001101100000010" => rgb <= "000000";
					when "00001101100000011" => rgb <= "000000";
					when "00001101100000100" => rgb <= "000000";
					when "00001101100000101" => rgb <= "000000";
					when "00001101100000110" => rgb <= "000000";
					when "00001101100000111" => rgb <= "000000";
					when "00001101100001000" => rgb <= "000000";
					when "00001101100001001" => rgb <= "000000";
					when "00001101100001010" => rgb <= "000000";
					when "00001101100001011" => rgb <= "000000";
					when "00001101100001100" => rgb <= "000000";
					when "00001101100001101" => rgb <= "000000";
					when "00001101100001110" => rgb <= "000000";
					when "00001101100001111" => rgb <= "000000";
					when "00001101100010000" => rgb <= "000000";
					when "00001101100010001" => rgb <= "000000";
					when "00001101100010010" => rgb <= "000000";
					when "00001101100010011" => rgb <= "000000";
					when "00001101100010100" => rgb <= "000000";
					when "00001101100010101" => rgb <= "000000";
					when "00001101100010110" => rgb <= "000000";
					when "00001101100010111" => rgb <= "000000";
					when "00001101100011000" => rgb <= "000000";
					when "00001101100011001" => rgb <= "000000";
					when "00001101100011010" => rgb <= "000000";
					when "00001101100011011" => rgb <= "000000";
					when "00001101100011100" => rgb <= "000000";
					when "00001101100011101" => rgb <= "000000";
					when "00001101100011110" => rgb <= "000000";
					when "00001101100011111" => rgb <= "000000";
					when "00001101100100000" => rgb <= "000000";
					when "00001101100100001" => rgb <= "000000";
					when "00001101100100010" => rgb <= "000000";
					when "00001101100100011" => rgb <= "000000";
					when "00001101100100100" => rgb <= "000000";
					when "00001101100100101" => rgb <= "000000";
					when "00001101100100110" => rgb <= "000000";
					when "00001101100100111" => rgb <= "000000";
					when "00001101100101000" => rgb <= "000000";
					when "00001101100101001" => rgb <= "000000";
					when "00001101100101010" => rgb <= "000000";
					when "00001101100101011" => rgb <= "000000";
					when "00001101100101100" => rgb <= "000000";
					when "00001101100101101" => rgb <= "000000";
					when "00001101100101110" => rgb <= "000000";
					when "00001101100101111" => rgb <= "000000";
					when "00001101100110000" => rgb <= "000000";
					when "00001101100110001" => rgb <= "000000";
					when "00001101100110010" => rgb <= "000000";
					when "00001101100110011" => rgb <= "000000";
					when "00001101100110100" => rgb <= "000000";
					when "00001101100110101" => rgb <= "000000";
					when "00001101100110110" => rgb <= "000000";
					when "00001101100110111" => rgb <= "000000";
					when "00001101100111000" => rgb <= "000000";
					when "00001101100111001" => rgb <= "000000";
					when "00001101100111010" => rgb <= "000000";
					when "00001101100111011" => rgb <= "000000";
					when "00001101100111100" => rgb <= "000000";
					when "00001101100111101" => rgb <= "000000";
					when "00001101100111110" => rgb <= "000000";
					when "00001101100111111" => rgb <= "000000";
					when "00001110000000000" => rgb <= "000000";
					when "00001110000000001" => rgb <= "000000";
					when "00001110000000010" => rgb <= "000000";
					when "00001110000000011" => rgb <= "000000";
					when "00001110000000100" => rgb <= "000000";
					when "00001110000000101" => rgb <= "000000";
					when "00001110000000110" => rgb <= "000000";
					when "00001110000000111" => rgb <= "000000";
					when "00001110000001000" => rgb <= "000000";
					when "00001110000001001" => rgb <= "000000";
					when "00001110000001010" => rgb <= "000000";
					when "00001110000001011" => rgb <= "000000";
					when "00001110000001100" => rgb <= "000000";
					when "00001110000001101" => rgb <= "000000";
					when "00001110000001110" => rgb <= "000000";
					when "00001110000001111" => rgb <= "000000";
					when "00001110000010000" => rgb <= "000000";
					when "00001110000010001" => rgb <= "000000";
					when "00001110000010010" => rgb <= "000000";
					when "00001110000010011" => rgb <= "000000";
					when "00001110000010100" => rgb <= "000000";
					when "00001110000010101" => rgb <= "000000";
					when "00001110000010110" => rgb <= "000000";
					when "00001110000010111" => rgb <= "000000";
					when "00001110000011000" => rgb <= "000000";
					when "00001110000011001" => rgb <= "000000";
					when "00001110000011010" => rgb <= "000000";
					when "00001110000011011" => rgb <= "000000";
					when "00001110000011100" => rgb <= "000000";
					when "00001110000011101" => rgb <= "000000";
					when "00001110000011110" => rgb <= "000000";
					when "00001110000011111" => rgb <= "000000";
					when "00001110000100000" => rgb <= "000000";
					when "00001110000100001" => rgb <= "000000";
					when "00001110000100010" => rgb <= "000000";
					when "00001110000100011" => rgb <= "000000";
					when "00001110000100100" => rgb <= "000000";
					when "00001110000100101" => rgb <= "000000";
					when "00001110000100110" => rgb <= "000000";
					when "00001110000100111" => rgb <= "000000";
					when "00001110000101000" => rgb <= "000000";
					when "00001110000101001" => rgb <= "000000";
					when "00001110000101010" => rgb <= "000000";
					when "00001110000101011" => rgb <= "000000";
					when "00001110000101100" => rgb <= "000000";
					when "00001110000101101" => rgb <= "000000";
					when "00001110000101110" => rgb <= "000000";
					when "00001110000101111" => rgb <= "000000";
					when "00001110000110000" => rgb <= "000000";
					when "00001110000110001" => rgb <= "000000";
					when "00001110000110010" => rgb <= "000000";
					when "00001110000110011" => rgb <= "000000";
					when "00001110000110100" => rgb <= "000000";
					when "00001110000110101" => rgb <= "000000";
					when "00001110000110110" => rgb <= "000000";
					when "00001110000110111" => rgb <= "000000";
					when "00001110000111000" => rgb <= "000000";
					when "00001110000111001" => rgb <= "000000";
					when "00001110000111010" => rgb <= "000000";
					when "00001110000111011" => rgb <= "000000";
					when "00001110000111100" => rgb <= "000000";
					when "00001110000111101" => rgb <= "000000";
					when "00001110000111110" => rgb <= "000000";
					when "00001110000111111" => rgb <= "000000";
					when "00001110001000000" => rgb <= "000000";
					when "00001110001000001" => rgb <= "000000";
					when "00001110001000010" => rgb <= "000000";
					when "00001110001000011" => rgb <= "000000";
					when "00001110001000100" => rgb <= "000000";
					when "00001110001000101" => rgb <= "000000";
					when "00001110001000110" => rgb <= "000000";
					when "00001110001000111" => rgb <= "000000";
					when "00001110001001000" => rgb <= "000000";
					when "00001110001001001" => rgb <= "000000";
					when "00001110001001010" => rgb <= "000000";
					when "00001110001001011" => rgb <= "000000";
					when "00001110001001100" => rgb <= "000000";
					when "00001110001001101" => rgb <= "000000";
					when "00001110001001110" => rgb <= "000000";
					when "00001110001001111" => rgb <= "000000";
					when "00001110001010000" => rgb <= "000000";
					when "00001110001010001" => rgb <= "000000";
					when "00001110001010010" => rgb <= "000000";
					when "00001110001010011" => rgb <= "000000";
					when "00001110001010100" => rgb <= "000000";
					when "00001110001010101" => rgb <= "000000";
					when "00001110001010110" => rgb <= "000000";
					when "00001110001010111" => rgb <= "000000";
					when "00001110001011000" => rgb <= "000000";
					when "00001110001011001" => rgb <= "000000";
					when "00001110001011010" => rgb <= "000000";
					when "00001110001011011" => rgb <= "000000";
					when "00001110001011100" => rgb <= "000000";
					when "00001110001011101" => rgb <= "000000";
					when "00001110001011110" => rgb <= "000000";
					when "00001110001011111" => rgb <= "000000";
					when "00001110001100000" => rgb <= "000000";
					when "00001110001100001" => rgb <= "000000";
					when "00001110001100010" => rgb <= "000000";
					when "00001110001100011" => rgb <= "000000";
					when "00001110001100100" => rgb <= "000000";
					when "00001110001100101" => rgb <= "000000";
					when "00001110001100110" => rgb <= "000000";
					when "00001110001100111" => rgb <= "000000";
					when "00001110001101000" => rgb <= "000000";
					when "00001110001101001" => rgb <= "000000";
					when "00001110001101010" => rgb <= "000000";
					when "00001110001101011" => rgb <= "000000";
					when "00001110001101100" => rgb <= "000000";
					when "00001110001101101" => rgb <= "000000";
					when "00001110001101110" => rgb <= "000000";
					when "00001110001101111" => rgb <= "000000";
					when "00001110001110000" => rgb <= "000000";
					when "00001110001110001" => rgb <= "000000";
					when "00001110001110010" => rgb <= "000000";
					when "00001110001110011" => rgb <= "000000";
					when "00001110001110100" => rgb <= "000000";
					when "00001110001110101" => rgb <= "000000";
					when "00001110001110110" => rgb <= "000000";
					when "00001110001110111" => rgb <= "000000";
					when "00001110001111000" => rgb <= "000000";
					when "00001110001111001" => rgb <= "000000";
					when "00001110001111010" => rgb <= "000000";
					when "00001110001111011" => rgb <= "000000";
					when "00001110001111100" => rgb <= "000000";
					when "00001110001111101" => rgb <= "000000";
					when "00001110001111110" => rgb <= "000000";
					when "00001110001111111" => rgb <= "000000";
					when "00001110010000000" => rgb <= "000000";
					when "00001110010000001" => rgb <= "000000";
					when "00001110010000010" => rgb <= "000000";
					when "00001110010000011" => rgb <= "000000";
					when "00001110010000100" => rgb <= "000000";
					when "00001110010000101" => rgb <= "000000";
					when "00001110010000110" => rgb <= "000000";
					when "00001110010000111" => rgb <= "000000";
					when "00001110010001000" => rgb <= "000000";
					when "00001110010001001" => rgb <= "000000";
					when "00001110010001010" => rgb <= "000000";
					when "00001110010001011" => rgb <= "000000";
					when "00001110010001100" => rgb <= "000000";
					when "00001110010001101" => rgb <= "000000";
					when "00001110010001110" => rgb <= "000000";
					when "00001110010001111" => rgb <= "000000";
					when "00001110010010000" => rgb <= "000000";
					when "00001110010010001" => rgb <= "000000";
					when "00001110010010010" => rgb <= "000000";
					when "00001110010010011" => rgb <= "000000";
					when "00001110010010100" => rgb <= "000000";
					when "00001110010010101" => rgb <= "000000";
					when "00001110010010110" => rgb <= "000000";
					when "00001110010010111" => rgb <= "000000";
					when "00001110010011000" => rgb <= "000000";
					when "00001110010011001" => rgb <= "000000";
					when "00001110010011010" => rgb <= "000000";
					when "00001110010011011" => rgb <= "000000";
					when "00001110010011100" => rgb <= "000000";
					when "00001110010011101" => rgb <= "000000";
					when "00001110010011110" => rgb <= "000000";
					when "00001110010011111" => rgb <= "000000";
					when "00001110010100000" => rgb <= "000000";
					when "00001110010100001" => rgb <= "000000";
					when "00001110010100010" => rgb <= "000000";
					when "00001110010100011" => rgb <= "000000";
					when "00001110010100100" => rgb <= "000000";
					when "00001110010100101" => rgb <= "000000";
					when "00001110010100110" => rgb <= "000000";
					when "00001110010100111" => rgb <= "000000";
					when "00001110010101000" => rgb <= "000000";
					when "00001110010101001" => rgb <= "000000";
					when "00001110010101010" => rgb <= "000000";
					when "00001110010101011" => rgb <= "000000";
					when "00001110010101100" => rgb <= "000000";
					when "00001110010101101" => rgb <= "000000";
					when "00001110010101110" => rgb <= "000000";
					when "00001110010101111" => rgb <= "000000";
					when "00001110010110000" => rgb <= "000000";
					when "00001110010110001" => rgb <= "000000";
					when "00001110010110010" => rgb <= "000000";
					when "00001110010110011" => rgb <= "000000";
					when "00001110010110100" => rgb <= "000000";
					when "00001110010110101" => rgb <= "000000";
					when "00001110010110110" => rgb <= "000000";
					when "00001110010110111" => rgb <= "000000";
					when "00001110010111000" => rgb <= "000000";
					when "00001110010111001" => rgb <= "000000";
					when "00001110010111010" => rgb <= "000000";
					when "00001110010111011" => rgb <= "000000";
					when "00001110010111100" => rgb <= "000000";
					when "00001110010111101" => rgb <= "000000";
					when "00001110010111110" => rgb <= "000000";
					when "00001110010111111" => rgb <= "000000";
					when "00001110011000000" => rgb <= "000000";
					when "00001110011000001" => rgb <= "000000";
					when "00001110011000010" => rgb <= "000000";
					when "00001110011000011" => rgb <= "000000";
					when "00001110011000100" => rgb <= "000000";
					when "00001110011000101" => rgb <= "000000";
					when "00001110011000110" => rgb <= "000000";
					when "00001110011000111" => rgb <= "000000";
					when "00001110011001000" => rgb <= "000000";
					when "00001110011001001" => rgb <= "000000";
					when "00001110011001010" => rgb <= "000000";
					when "00001110011001011" => rgb <= "000000";
					when "00001110011001100" => rgb <= "000000";
					when "00001110011001101" => rgb <= "000000";
					when "00001110011001110" => rgb <= "000000";
					when "00001110011001111" => rgb <= "000000";
					when "00001110011010000" => rgb <= "000000";
					when "00001110011010001" => rgb <= "000000";
					when "00001110011010010" => rgb <= "000000";
					when "00001110011010011" => rgb <= "000000";
					when "00001110011010100" => rgb <= "000000";
					when "00001110011010101" => rgb <= "000000";
					when "00001110011010110" => rgb <= "000000";
					when "00001110011010111" => rgb <= "000000";
					when "00001110011011000" => rgb <= "000000";
					when "00001110011011001" => rgb <= "000000";
					when "00001110011011010" => rgb <= "000000";
					when "00001110011011011" => rgb <= "000000";
					when "00001110011011100" => rgb <= "000000";
					when "00001110011011101" => rgb <= "000000";
					when "00001110011011110" => rgb <= "000000";
					when "00001110011011111" => rgb <= "000000";
					when "00001110011100000" => rgb <= "000000";
					when "00001110011100001" => rgb <= "000000";
					when "00001110011100010" => rgb <= "000000";
					when "00001110011100011" => rgb <= "000000";
					when "00001110011100100" => rgb <= "000000";
					when "00001110011100101" => rgb <= "000000";
					when "00001110011100110" => rgb <= "000000";
					when "00001110011100111" => rgb <= "000000";
					when "00001110011101000" => rgb <= "000000";
					when "00001110011101001" => rgb <= "000000";
					when "00001110011101010" => rgb <= "000000";
					when "00001110011101011" => rgb <= "000000";
					when "00001110011101100" => rgb <= "000000";
					when "00001110011101101" => rgb <= "000000";
					when "00001110011101110" => rgb <= "000000";
					when "00001110011101111" => rgb <= "000000";
					when "00001110011110000" => rgb <= "000000";
					when "00001110011110001" => rgb <= "000000";
					when "00001110011110010" => rgb <= "000000";
					when "00001110011110011" => rgb <= "000000";
					when "00001110011110100" => rgb <= "000000";
					when "00001110011110101" => rgb <= "000000";
					when "00001110011110110" => rgb <= "000000";
					when "00001110011110111" => rgb <= "000000";
					when "00001110011111000" => rgb <= "000000";
					when "00001110011111001" => rgb <= "000000";
					when "00001110011111010" => rgb <= "000000";
					when "00001110011111011" => rgb <= "000000";
					when "00001110011111100" => rgb <= "000000";
					when "00001110011111101" => rgb <= "000000";
					when "00001110011111110" => rgb <= "000000";
					when "00001110011111111" => rgb <= "000000";
					when "00001110100000000" => rgb <= "000000";
					when "00001110100000001" => rgb <= "000000";
					when "00001110100000010" => rgb <= "000000";
					when "00001110100000011" => rgb <= "000000";
					when "00001110100000100" => rgb <= "000000";
					when "00001110100000101" => rgb <= "000000";
					when "00001110100000110" => rgb <= "000000";
					when "00001110100000111" => rgb <= "000000";
					when "00001110100001000" => rgb <= "000000";
					when "00001110100001001" => rgb <= "000000";
					when "00001110100001010" => rgb <= "000000";
					when "00001110100001011" => rgb <= "000000";
					when "00001110100001100" => rgb <= "000000";
					when "00001110100001101" => rgb <= "000000";
					when "00001110100001110" => rgb <= "000000";
					when "00001110100001111" => rgb <= "000000";
					when "00001110100010000" => rgb <= "000000";
					when "00001110100010001" => rgb <= "000000";
					when "00001110100010010" => rgb <= "000000";
					when "00001110100010011" => rgb <= "000000";
					when "00001110100010100" => rgb <= "000000";
					when "00001110100010101" => rgb <= "000000";
					when "00001110100010110" => rgb <= "000000";
					when "00001110100010111" => rgb <= "000000";
					when "00001110100011000" => rgb <= "000000";
					when "00001110100011001" => rgb <= "000000";
					when "00001110100011010" => rgb <= "000000";
					when "00001110100011011" => rgb <= "000000";
					when "00001110100011100" => rgb <= "000000";
					when "00001110100011101" => rgb <= "000000";
					when "00001110100011110" => rgb <= "000000";
					when "00001110100011111" => rgb <= "000000";
					when "00001110100100000" => rgb <= "000000";
					when "00001110100100001" => rgb <= "000000";
					when "00001110100100010" => rgb <= "000000";
					when "00001110100100011" => rgb <= "000000";
					when "00001110100100100" => rgb <= "000000";
					when "00001110100100101" => rgb <= "000000";
					when "00001110100100110" => rgb <= "000000";
					when "00001110100100111" => rgb <= "000000";
					when "00001110100101000" => rgb <= "000000";
					when "00001110100101001" => rgb <= "000000";
					when "00001110100101010" => rgb <= "000000";
					when "00001110100101011" => rgb <= "000000";
					when "00001110100101100" => rgb <= "000000";
					when "00001110100101101" => rgb <= "000000";
					when "00001110100101110" => rgb <= "000000";
					when "00001110100101111" => rgb <= "000000";
					when "00001110100110000" => rgb <= "000000";
					when "00001110100110001" => rgb <= "000000";
					when "00001110100110010" => rgb <= "000000";
					when "00001110100110011" => rgb <= "000000";
					when "00001110100110100" => rgb <= "000000";
					when "00001110100110101" => rgb <= "000000";
					when "00001110100110110" => rgb <= "000000";
					when "00001110100110111" => rgb <= "000000";
					when "00001110100111000" => rgb <= "000000";
					when "00001110100111001" => rgb <= "000000";
					when "00001110100111010" => rgb <= "000000";
					when "00001110100111011" => rgb <= "000000";
					when "00001110100111100" => rgb <= "000000";
					when "00001110100111101" => rgb <= "000000";
					when "00001110100111110" => rgb <= "000000";
					when "00001110100111111" => rgb <= "000000";
					when "00001111000000000" => rgb <= "000000";
					when "00001111000000001" => rgb <= "000000";
					when "00001111000000010" => rgb <= "000000";
					when "00001111000000011" => rgb <= "000000";
					when "00001111000000100" => rgb <= "000000";
					when "00001111000000101" => rgb <= "000000";
					when "00001111000000110" => rgb <= "000000";
					when "00001111000000111" => rgb <= "000000";
					when "00001111000001000" => rgb <= "000000";
					when "00001111000001001" => rgb <= "000000";
					when "00001111000001010" => rgb <= "000000";
					when "00001111000001011" => rgb <= "000000";
					when "00001111000001100" => rgb <= "000000";
					when "00001111000001101" => rgb <= "000000";
					when "00001111000001110" => rgb <= "000000";
					when "00001111000001111" => rgb <= "000000";
					when "00001111000010000" => rgb <= "000000";
					when "00001111000010001" => rgb <= "000000";
					when "00001111000010010" => rgb <= "000000";
					when "00001111000010011" => rgb <= "000000";
					when "00001111000010100" => rgb <= "000000";
					when "00001111000010101" => rgb <= "000000";
					when "00001111000010110" => rgb <= "000000";
					when "00001111000010111" => rgb <= "000000";
					when "00001111000011000" => rgb <= "000000";
					when "00001111000011001" => rgb <= "000000";
					when "00001111000011010" => rgb <= "000000";
					when "00001111000011011" => rgb <= "000000";
					when "00001111000011100" => rgb <= "000000";
					when "00001111000011101" => rgb <= "000000";
					when "00001111000011110" => rgb <= "000000";
					when "00001111000011111" => rgb <= "000000";
					when "00001111000100000" => rgb <= "000000";
					when "00001111000100001" => rgb <= "000000";
					when "00001111000100010" => rgb <= "000000";
					when "00001111000100011" => rgb <= "000000";
					when "00001111000100100" => rgb <= "000000";
					when "00001111000100101" => rgb <= "000000";
					when "00001111000100110" => rgb <= "000000";
					when "00001111000100111" => rgb <= "000000";
					when "00001111000101000" => rgb <= "000000";
					when "00001111000101001" => rgb <= "000000";
					when "00001111000101010" => rgb <= "000000";
					when "00001111000101011" => rgb <= "000000";
					when "00001111000101100" => rgb <= "000000";
					when "00001111000101101" => rgb <= "000000";
					when "00001111000101110" => rgb <= "000000";
					when "00001111000101111" => rgb <= "000000";
					when "00001111000110000" => rgb <= "000000";
					when "00001111000110001" => rgb <= "000000";
					when "00001111000110010" => rgb <= "000000";
					when "00001111000110011" => rgb <= "000000";
					when "00001111000110100" => rgb <= "000000";
					when "00001111000110101" => rgb <= "000000";
					when "00001111000110110" => rgb <= "000000";
					when "00001111000110111" => rgb <= "000000";
					when "00001111000111000" => rgb <= "000000";
					when "00001111000111001" => rgb <= "000000";
					when "00001111000111010" => rgb <= "000000";
					when "00001111000111011" => rgb <= "000000";
					when "00001111000111100" => rgb <= "000000";
					when "00001111000111101" => rgb <= "000000";
					when "00001111000111110" => rgb <= "000000";
					when "00001111000111111" => rgb <= "000000";
					when "00001111001000000" => rgb <= "000000";
					when "00001111001000001" => rgb <= "000000";
					when "00001111001000010" => rgb <= "000000";
					when "00001111001000011" => rgb <= "000000";
					when "00001111001000100" => rgb <= "000000";
					when "00001111001000101" => rgb <= "000000";
					when "00001111001000110" => rgb <= "000000";
					when "00001111001000111" => rgb <= "000000";
					when "00001111001001000" => rgb <= "000000";
					when "00001111001001001" => rgb <= "000000";
					when "00001111001001010" => rgb <= "000000";
					when "00001111001001011" => rgb <= "000000";
					when "00001111001001100" => rgb <= "000000";
					when "00001111001001101" => rgb <= "000000";
					when "00001111001001110" => rgb <= "000000";
					when "00001111001001111" => rgb <= "000000";
					when "00001111001010000" => rgb <= "000000";
					when "00001111001010001" => rgb <= "000000";
					when "00001111001010010" => rgb <= "000000";
					when "00001111001010011" => rgb <= "000000";
					when "00001111001010100" => rgb <= "000000";
					when "00001111001010101" => rgb <= "000000";
					when "00001111001010110" => rgb <= "000000";
					when "00001111001010111" => rgb <= "000000";
					when "00001111001011000" => rgb <= "000000";
					when "00001111001011001" => rgb <= "000000";
					when "00001111001011010" => rgb <= "000000";
					when "00001111001011011" => rgb <= "000000";
					when "00001111001011100" => rgb <= "000000";
					when "00001111001011101" => rgb <= "000000";
					when "00001111001011110" => rgb <= "000000";
					when "00001111001011111" => rgb <= "000000";
					when "00001111001100000" => rgb <= "000000";
					when "00001111001100001" => rgb <= "000000";
					when "00001111001100010" => rgb <= "000000";
					when "00001111001100011" => rgb <= "000000";
					when "00001111001100100" => rgb <= "000000";
					when "00001111001100101" => rgb <= "000000";
					when "00001111001100110" => rgb <= "000000";
					when "00001111001100111" => rgb <= "000000";
					when "00001111001101000" => rgb <= "000000";
					when "00001111001101001" => rgb <= "000000";
					when "00001111001101010" => rgb <= "000000";
					when "00001111001101011" => rgb <= "000000";
					when "00001111001101100" => rgb <= "000000";
					when "00001111001101101" => rgb <= "000000";
					when "00001111001101110" => rgb <= "000000";
					when "00001111001101111" => rgb <= "000000";
					when "00001111001110000" => rgb <= "000000";
					when "00001111001110001" => rgb <= "000000";
					when "00001111001110010" => rgb <= "000000";
					when "00001111001110011" => rgb <= "000000";
					when "00001111001110100" => rgb <= "000000";
					when "00001111001110101" => rgb <= "000000";
					when "00001111001110110" => rgb <= "000000";
					when "00001111001110111" => rgb <= "000000";
					when "00001111001111000" => rgb <= "000000";
					when "00001111001111001" => rgb <= "000000";
					when "00001111001111010" => rgb <= "000000";
					when "00001111001111011" => rgb <= "000000";
					when "00001111001111100" => rgb <= "000000";
					when "00001111001111101" => rgb <= "000000";
					when "00001111001111110" => rgb <= "000000";
					when "00001111001111111" => rgb <= "000000";
					when "00001111010000000" => rgb <= "000000";
					when "00001111010000001" => rgb <= "000000";
					when "00001111010000010" => rgb <= "000000";
					when "00001111010000011" => rgb <= "000000";
					when "00001111010000100" => rgb <= "000000";
					when "00001111010000101" => rgb <= "000000";
					when "00001111010000110" => rgb <= "000000";
					when "00001111010000111" => rgb <= "000000";
					when "00001111010001000" => rgb <= "000000";
					when "00001111010001001" => rgb <= "000000";
					when "00001111010001010" => rgb <= "000000";
					when "00001111010001011" => rgb <= "000000";
					when "00001111010001100" => rgb <= "000000";
					when "00001111010001101" => rgb <= "000000";
					when "00001111010001110" => rgb <= "000000";
					when "00001111010001111" => rgb <= "000000";
					when "00001111010010000" => rgb <= "000000";
					when "00001111010010001" => rgb <= "000000";
					when "00001111010010010" => rgb <= "000000";
					when "00001111010010011" => rgb <= "000000";
					when "00001111010010100" => rgb <= "000000";
					when "00001111010010101" => rgb <= "000000";
					when "00001111010010110" => rgb <= "000000";
					when "00001111010010111" => rgb <= "000000";
					when "00001111010011000" => rgb <= "000000";
					when "00001111010011001" => rgb <= "000000";
					when "00001111010011010" => rgb <= "000000";
					when "00001111010011011" => rgb <= "000000";
					when "00001111010011100" => rgb <= "000000";
					when "00001111010011101" => rgb <= "000000";
					when "00001111010011110" => rgb <= "000000";
					when "00001111010011111" => rgb <= "000000";
					when "00001111010100000" => rgb <= "000000";
					when "00001111010100001" => rgb <= "000000";
					when "00001111010100010" => rgb <= "000000";
					when "00001111010100011" => rgb <= "000000";
					when "00001111010100100" => rgb <= "000000";
					when "00001111010100101" => rgb <= "000000";
					when "00001111010100110" => rgb <= "000000";
					when "00001111010100111" => rgb <= "000000";
					when "00001111010101000" => rgb <= "000000";
					when "00001111010101001" => rgb <= "000000";
					when "00001111010101010" => rgb <= "000000";
					when "00001111010101011" => rgb <= "000000";
					when "00001111010101100" => rgb <= "000000";
					when "00001111010101101" => rgb <= "000000";
					when "00001111010101110" => rgb <= "000000";
					when "00001111010101111" => rgb <= "000000";
					when "00001111010110000" => rgb <= "000000";
					when "00001111010110001" => rgb <= "000000";
					when "00001111010110010" => rgb <= "000000";
					when "00001111010110011" => rgb <= "000000";
					when "00001111010110100" => rgb <= "000000";
					when "00001111010110101" => rgb <= "000000";
					when "00001111010110110" => rgb <= "000000";
					when "00001111010110111" => rgb <= "000000";
					when "00001111010111000" => rgb <= "000000";
					when "00001111010111001" => rgb <= "000000";
					when "00001111010111010" => rgb <= "000000";
					when "00001111010111011" => rgb <= "000000";
					when "00001111010111100" => rgb <= "000000";
					when "00001111010111101" => rgb <= "000000";
					when "00001111010111110" => rgb <= "000000";
					when "00001111010111111" => rgb <= "000000";
					when "00001111011000000" => rgb <= "000000";
					when "00001111011000001" => rgb <= "000000";
					when "00001111011000010" => rgb <= "000000";
					when "00001111011000011" => rgb <= "000000";
					when "00001111011000100" => rgb <= "000000";
					when "00001111011000101" => rgb <= "000000";
					when "00001111011000110" => rgb <= "000000";
					when "00001111011000111" => rgb <= "000000";
					when "00001111011001000" => rgb <= "000000";
					when "00001111011001001" => rgb <= "000000";
					when "00001111011001010" => rgb <= "000000";
					when "00001111011001011" => rgb <= "000000";
					when "00001111011001100" => rgb <= "000000";
					when "00001111011001101" => rgb <= "000000";
					when "00001111011001110" => rgb <= "000000";
					when "00001111011001111" => rgb <= "000000";
					when "00001111011010000" => rgb <= "000000";
					when "00001111011010001" => rgb <= "000000";
					when "00001111011010010" => rgb <= "000000";
					when "00001111011010011" => rgb <= "000000";
					when "00001111011010100" => rgb <= "000000";
					when "00001111011010101" => rgb <= "000000";
					when "00001111011010110" => rgb <= "000000";
					when "00001111011010111" => rgb <= "000000";
					when "00001111011011000" => rgb <= "000000";
					when "00001111011011001" => rgb <= "000000";
					when "00001111011011010" => rgb <= "000000";
					when "00001111011011011" => rgb <= "000000";
					when "00001111011011100" => rgb <= "000000";
					when "00001111011011101" => rgb <= "000000";
					when "00001111011011110" => rgb <= "000000";
					when "00001111011011111" => rgb <= "000000";
					when "00001111011100000" => rgb <= "000000";
					when "00001111011100001" => rgb <= "000000";
					when "00001111011100010" => rgb <= "000000";
					when "00001111011100011" => rgb <= "000000";
					when "00001111011100100" => rgb <= "000000";
					when "00001111011100101" => rgb <= "000000";
					when "00001111011100110" => rgb <= "000000";
					when "00001111011100111" => rgb <= "000000";
					when "00001111011101000" => rgb <= "000000";
					when "00001111011101001" => rgb <= "000000";
					when "00001111011101010" => rgb <= "000000";
					when "00001111011101011" => rgb <= "000000";
					when "00001111011101100" => rgb <= "000000";
					when "00001111011101101" => rgb <= "000000";
					when "00001111011101110" => rgb <= "000000";
					when "00001111011101111" => rgb <= "000000";
					when "00001111011110000" => rgb <= "000000";
					when "00001111011110001" => rgb <= "000000";
					when "00001111011110010" => rgb <= "000000";
					when "00001111011110011" => rgb <= "000000";
					when "00001111011110100" => rgb <= "000000";
					when "00001111011110101" => rgb <= "000000";
					when "00001111011110110" => rgb <= "000000";
					when "00001111011110111" => rgb <= "000000";
					when "00001111011111000" => rgb <= "000000";
					when "00001111011111001" => rgb <= "000000";
					when "00001111011111010" => rgb <= "000000";
					when "00001111011111011" => rgb <= "000000";
					when "00001111011111100" => rgb <= "000000";
					when "00001111011111101" => rgb <= "000000";
					when "00001111011111110" => rgb <= "000000";
					when "00001111011111111" => rgb <= "000000";
					when "00001111100000000" => rgb <= "000000";
					when "00001111100000001" => rgb <= "000000";
					when "00001111100000010" => rgb <= "000000";
					when "00001111100000011" => rgb <= "000000";
					when "00001111100000100" => rgb <= "000000";
					when "00001111100000101" => rgb <= "000000";
					when "00001111100000110" => rgb <= "000000";
					when "00001111100000111" => rgb <= "000000";
					when "00001111100001000" => rgb <= "000000";
					when "00001111100001001" => rgb <= "000000";
					when "00001111100001010" => rgb <= "000000";
					when "00001111100001011" => rgb <= "000000";
					when "00001111100001100" => rgb <= "000000";
					when "00001111100001101" => rgb <= "000000";
					when "00001111100001110" => rgb <= "000000";
					when "00001111100001111" => rgb <= "000000";
					when "00001111100010000" => rgb <= "000000";
					when "00001111100010001" => rgb <= "000000";
					when "00001111100010010" => rgb <= "000000";
					when "00001111100010011" => rgb <= "000000";
					when "00001111100010100" => rgb <= "000000";
					when "00001111100010101" => rgb <= "000000";
					when "00001111100010110" => rgb <= "000000";
					when "00001111100010111" => rgb <= "000000";
					when "00001111100011000" => rgb <= "000000";
					when "00001111100011001" => rgb <= "000000";
					when "00001111100011010" => rgb <= "000000";
					when "00001111100011011" => rgb <= "000000";
					when "00001111100011100" => rgb <= "000000";
					when "00001111100011101" => rgb <= "000000";
					when "00001111100011110" => rgb <= "000000";
					when "00001111100011111" => rgb <= "000000";
					when "00001111100100000" => rgb <= "000000";
					when "00001111100100001" => rgb <= "000000";
					when "00001111100100010" => rgb <= "000000";
					when "00001111100100011" => rgb <= "000000";
					when "00001111100100100" => rgb <= "000000";
					when "00001111100100101" => rgb <= "000000";
					when "00001111100100110" => rgb <= "000000";
					when "00001111100100111" => rgb <= "000000";
					when "00001111100101000" => rgb <= "000000";
					when "00001111100101001" => rgb <= "000000";
					when "00001111100101010" => rgb <= "000000";
					when "00001111100101011" => rgb <= "000000";
					when "00001111100101100" => rgb <= "000000";
					when "00001111100101101" => rgb <= "000000";
					when "00001111100101110" => rgb <= "000000";
					when "00001111100101111" => rgb <= "000000";
					when "00001111100110000" => rgb <= "000000";
					when "00001111100110001" => rgb <= "000000";
					when "00001111100110010" => rgb <= "000000";
					when "00001111100110011" => rgb <= "000000";
					when "00001111100110100" => rgb <= "000000";
					when "00001111100110101" => rgb <= "000000";
					when "00001111100110110" => rgb <= "000000";
					when "00001111100110111" => rgb <= "000000";
					when "00001111100111000" => rgb <= "000000";
					when "00001111100111001" => rgb <= "000000";
					when "00001111100111010" => rgb <= "000000";
					when "00001111100111011" => rgb <= "000000";
					when "00001111100111100" => rgb <= "000000";
					when "00001111100111101" => rgb <= "000000";
					when "00001111100111110" => rgb <= "000000";
					when "00001111100111111" => rgb <= "000000";
					when "00010000000000000" => rgb <= "000000";
					when "00010000000000001" => rgb <= "000000";
					when "00010000000000010" => rgb <= "000000";
					when "00010000000000011" => rgb <= "000000";
					when "00010000000000100" => rgb <= "000000";
					when "00010000000000101" => rgb <= "000000";
					when "00010000000000110" => rgb <= "000000";
					when "00010000000000111" => rgb <= "000000";
					when "00010000000001000" => rgb <= "000000";
					when "00010000000001001" => rgb <= "000000";
					when "00010000000001010" => rgb <= "000000";
					when "00010000000001011" => rgb <= "000000";
					when "00010000000001100" => rgb <= "000000";
					when "00010000000001101" => rgb <= "000000";
					when "00010000000001110" => rgb <= "000000";
					when "00010000000001111" => rgb <= "000000";
					when "00010000000010000" => rgb <= "000000";
					when "00010000000010001" => rgb <= "000000";
					when "00010000000010010" => rgb <= "000000";
					when "00010000000010011" => rgb <= "000000";
					when "00010000000010100" => rgb <= "000000";
					when "00010000000010101" => rgb <= "000000";
					when "00010000000010110" => rgb <= "000000";
					when "00010000000010111" => rgb <= "000000";
					when "00010000000011000" => rgb <= "000000";
					when "00010000000011001" => rgb <= "000000";
					when "00010000000011010" => rgb <= "000000";
					when "00010000000011011" => rgb <= "000000";
					when "00010000000011100" => rgb <= "000000";
					when "00010000000011101" => rgb <= "000000";
					when "00010000000011110" => rgb <= "000000";
					when "00010000000011111" => rgb <= "000000";
					when "00010000000100000" => rgb <= "000000";
					when "00010000000100001" => rgb <= "000000";
					when "00010000000100010" => rgb <= "000000";
					when "00010000000100011" => rgb <= "000000";
					when "00010000000100100" => rgb <= "000000";
					when "00010000000100101" => rgb <= "000000";
					when "00010000000100110" => rgb <= "000000";
					when "00010000000100111" => rgb <= "000000";
					when "00010000000101000" => rgb <= "000000";
					when "00010000000101001" => rgb <= "000000";
					when "00010000000101010" => rgb <= "000000";
					when "00010000000101011" => rgb <= "000000";
					when "00010000000101100" => rgb <= "000000";
					when "00010000000101101" => rgb <= "000000";
					when "00010000000101110" => rgb <= "000000";
					when "00010000000101111" => rgb <= "000000";
					when "00010000000110000" => rgb <= "000000";
					when "00010000000110001" => rgb <= "000000";
					when "00010000000110010" => rgb <= "000000";
					when "00010000000110011" => rgb <= "000000";
					when "00010000000110100" => rgb <= "000000";
					when "00010000000110101" => rgb <= "000000";
					when "00010000000110110" => rgb <= "000000";
					when "00010000000110111" => rgb <= "000000";
					when "00010000000111000" => rgb <= "000000";
					when "00010000000111001" => rgb <= "000000";
					when "00010000000111010" => rgb <= "000000";
					when "00010000000111011" => rgb <= "000000";
					when "00010000000111100" => rgb <= "000000";
					when "00010000000111101" => rgb <= "000000";
					when "00010000000111110" => rgb <= "000000";
					when "00010000000111111" => rgb <= "000000";
					when "00010000001000000" => rgb <= "000000";
					when "00010000001000001" => rgb <= "000000";
					when "00010000001000010" => rgb <= "000000";
					when "00010000001000011" => rgb <= "000000";
					when "00010000001000100" => rgb <= "000000";
					when "00010000001000101" => rgb <= "000000";
					when "00010000001000110" => rgb <= "000000";
					when "00010000001000111" => rgb <= "000000";
					when "00010000001001000" => rgb <= "000000";
					when "00010000001001001" => rgb <= "000000";
					when "00010000001001010" => rgb <= "000000";
					when "00010000001001011" => rgb <= "000000";
					when "00010000001001100" => rgb <= "000000";
					when "00010000001001101" => rgb <= "000000";
					when "00010000001001110" => rgb <= "000000";
					when "00010000001001111" => rgb <= "000000";
					when "00010000001010000" => rgb <= "000000";
					when "00010000001010001" => rgb <= "000000";
					when "00010000001010010" => rgb <= "000000";
					when "00010000001010011" => rgb <= "000000";
					when "00010000001010100" => rgb <= "000000";
					when "00010000001010101" => rgb <= "000000";
					when "00010000001010110" => rgb <= "000000";
					when "00010000001010111" => rgb <= "000000";
					when "00010000001011000" => rgb <= "000000";
					when "00010000001011001" => rgb <= "000000";
					when "00010000001011010" => rgb <= "000000";
					when "00010000001011011" => rgb <= "000000";
					when "00010000001011100" => rgb <= "000000";
					when "00010000001011101" => rgb <= "000000";
					when "00010000001011110" => rgb <= "000000";
					when "00010000001011111" => rgb <= "000000";
					when "00010000001100000" => rgb <= "000000";
					when "00010000001100001" => rgb <= "000000";
					when "00010000001100010" => rgb <= "000000";
					when "00010000001100011" => rgb <= "000000";
					when "00010000001100100" => rgb <= "000000";
					when "00010000001100101" => rgb <= "000000";
					when "00010000001100110" => rgb <= "000000";
					when "00010000001100111" => rgb <= "000000";
					when "00010000001101000" => rgb <= "000000";
					when "00010000001101001" => rgb <= "000000";
					when "00010000001101010" => rgb <= "000000";
					when "00010000001101011" => rgb <= "000000";
					when "00010000001101100" => rgb <= "000000";
					when "00010000001101101" => rgb <= "000000";
					when "00010000001101110" => rgb <= "000000";
					when "00010000001101111" => rgb <= "000000";
					when "00010000001110000" => rgb <= "000000";
					when "00010000001110001" => rgb <= "000000";
					when "00010000001110010" => rgb <= "000000";
					when "00010000001110011" => rgb <= "000000";
					when "00010000001110100" => rgb <= "000000";
					when "00010000001110101" => rgb <= "000000";
					when "00010000001110110" => rgb <= "000000";
					when "00010000001110111" => rgb <= "000000";
					when "00010000001111000" => rgb <= "000000";
					when "00010000001111001" => rgb <= "000000";
					when "00010000001111010" => rgb <= "000000";
					when "00010000001111011" => rgb <= "000000";
					when "00010000001111100" => rgb <= "000000";
					when "00010000001111101" => rgb <= "000000";
					when "00010000001111110" => rgb <= "000000";
					when "00010000001111111" => rgb <= "000000";
					when "00010000010000000" => rgb <= "000000";
					when "00010000010000001" => rgb <= "000000";
					when "00010000010000010" => rgb <= "000000";
					when "00010000010000011" => rgb <= "000000";
					when "00010000010000100" => rgb <= "000000";
					when "00010000010000101" => rgb <= "000000";
					when "00010000010000110" => rgb <= "000000";
					when "00010000010000111" => rgb <= "000000";
					when "00010000010001000" => rgb <= "000000";
					when "00010000010001001" => rgb <= "000000";
					when "00010000010001010" => rgb <= "000000";
					when "00010000010001011" => rgb <= "000000";
					when "00010000010001100" => rgb <= "000000";
					when "00010000010001101" => rgb <= "000000";
					when "00010000010001110" => rgb <= "000000";
					when "00010000010001111" => rgb <= "000000";
					when "00010000010010000" => rgb <= "000000";
					when "00010000010010001" => rgb <= "000000";
					when "00010000010010010" => rgb <= "000000";
					when "00010000010010011" => rgb <= "000000";
					when "00010000010010100" => rgb <= "000000";
					when "00010000010010101" => rgb <= "000000";
					when "00010000010010110" => rgb <= "000000";
					when "00010000010010111" => rgb <= "000000";
					when "00010000010011000" => rgb <= "000000";
					when "00010000010011001" => rgb <= "000000";
					when "00010000010011010" => rgb <= "000000";
					when "00010000010011011" => rgb <= "000000";
					when "00010000010011100" => rgb <= "000000";
					when "00010000010011101" => rgb <= "000000";
					when "00010000010011110" => rgb <= "000000";
					when "00010000010011111" => rgb <= "000000";
					when "00010000010100000" => rgb <= "000000";
					when "00010000010100001" => rgb <= "000000";
					when "00010000010100010" => rgb <= "000000";
					when "00010000010100011" => rgb <= "000000";
					when "00010000010100100" => rgb <= "000000";
					when "00010000010100101" => rgb <= "000000";
					when "00010000010100110" => rgb <= "000000";
					when "00010000010100111" => rgb <= "000000";
					when "00010000010101000" => rgb <= "000000";
					when "00010000010101001" => rgb <= "000000";
					when "00010000010101010" => rgb <= "000000";
					when "00010000010101011" => rgb <= "000000";
					when "00010000010101100" => rgb <= "000000";
					when "00010000010101101" => rgb <= "000000";
					when "00010000010101110" => rgb <= "000000";
					when "00010000010101111" => rgb <= "000000";
					when "00010000010110000" => rgb <= "000000";
					when "00010000010110001" => rgb <= "000000";
					when "00010000010110010" => rgb <= "000000";
					when "00010000010110011" => rgb <= "000000";
					when "00010000010110100" => rgb <= "000000";
					when "00010000010110101" => rgb <= "000000";
					when "00010000010110110" => rgb <= "000000";
					when "00010000010110111" => rgb <= "000000";
					when "00010000010111000" => rgb <= "000000";
					when "00010000010111001" => rgb <= "000000";
					when "00010000010111010" => rgb <= "000000";
					when "00010000010111011" => rgb <= "000000";
					when "00010000010111100" => rgb <= "000000";
					when "00010000010111101" => rgb <= "000000";
					when "00010000010111110" => rgb <= "000000";
					when "00010000010111111" => rgb <= "000000";
					when "00010000011000000" => rgb <= "000000";
					when "00010000011000001" => rgb <= "000000";
					when "00010000011000010" => rgb <= "000000";
					when "00010000011000011" => rgb <= "000000";
					when "00010000011000100" => rgb <= "000000";
					when "00010000011000101" => rgb <= "000000";
					when "00010000011000110" => rgb <= "000000";
					when "00010000011000111" => rgb <= "000000";
					when "00010000011001000" => rgb <= "000000";
					when "00010000011001001" => rgb <= "000000";
					when "00010000011001010" => rgb <= "000000";
					when "00010000011001011" => rgb <= "000000";
					when "00010000011001100" => rgb <= "000000";
					when "00010000011001101" => rgb <= "000000";
					when "00010000011001110" => rgb <= "000000";
					when "00010000011001111" => rgb <= "000000";
					when "00010000011010000" => rgb <= "000000";
					when "00010000011010001" => rgb <= "000000";
					when "00010000011010010" => rgb <= "000000";
					when "00010000011010011" => rgb <= "000000";
					when "00010000011010100" => rgb <= "000000";
					when "00010000011010101" => rgb <= "000000";
					when "00010000011010110" => rgb <= "000000";
					when "00010000011010111" => rgb <= "000000";
					when "00010000011011000" => rgb <= "000000";
					when "00010000011011001" => rgb <= "000000";
					when "00010000011011010" => rgb <= "000000";
					when "00010000011011011" => rgb <= "000000";
					when "00010000011011100" => rgb <= "000000";
					when "00010000011011101" => rgb <= "000000";
					when "00010000011011110" => rgb <= "000000";
					when "00010000011011111" => rgb <= "000000";
					when "00010000011100000" => rgb <= "000000";
					when "00010000011100001" => rgb <= "000000";
					when "00010000011100010" => rgb <= "000000";
					when "00010000011100011" => rgb <= "000000";
					when "00010000011100100" => rgb <= "000000";
					when "00010000011100101" => rgb <= "000000";
					when "00010000011100110" => rgb <= "000000";
					when "00010000011100111" => rgb <= "000000";
					when "00010000011101000" => rgb <= "000000";
					when "00010000011101001" => rgb <= "000000";
					when "00010000011101010" => rgb <= "000000";
					when "00010000011101011" => rgb <= "000000";
					when "00010000011101100" => rgb <= "000000";
					when "00010000011101101" => rgb <= "000000";
					when "00010000011101110" => rgb <= "000000";
					when "00010000011101111" => rgb <= "000000";
					when "00010000011110000" => rgb <= "000000";
					when "00010000011110001" => rgb <= "000000";
					when "00010000011110010" => rgb <= "000000";
					when "00010000011110011" => rgb <= "000000";
					when "00010000011110100" => rgb <= "000000";
					when "00010000011110101" => rgb <= "000000";
					when "00010000011110110" => rgb <= "000000";
					when "00010000011110111" => rgb <= "000000";
					when "00010000011111000" => rgb <= "000000";
					when "00010000011111001" => rgb <= "000000";
					when "00010000011111010" => rgb <= "000000";
					when "00010000011111011" => rgb <= "000000";
					when "00010000011111100" => rgb <= "000000";
					when "00010000011111101" => rgb <= "000000";
					when "00010000011111110" => rgb <= "000000";
					when "00010000011111111" => rgb <= "000000";
					when "00010000100000000" => rgb <= "000000";
					when "00010000100000001" => rgb <= "000000";
					when "00010000100000010" => rgb <= "000000";
					when "00010000100000011" => rgb <= "000000";
					when "00010000100000100" => rgb <= "000000";
					when "00010000100000101" => rgb <= "000000";
					when "00010000100000110" => rgb <= "000000";
					when "00010000100000111" => rgb <= "000000";
					when "00010000100001000" => rgb <= "000000";
					when "00010000100001001" => rgb <= "000000";
					when "00010000100001010" => rgb <= "000000";
					when "00010000100001011" => rgb <= "000000";
					when "00010000100001100" => rgb <= "000000";
					when "00010000100001101" => rgb <= "000000";
					when "00010000100001110" => rgb <= "000000";
					when "00010000100001111" => rgb <= "000000";
					when "00010000100010000" => rgb <= "000000";
					when "00010000100010001" => rgb <= "000000";
					when "00010000100010010" => rgb <= "000000";
					when "00010000100010011" => rgb <= "000000";
					when "00010000100010100" => rgb <= "000000";
					when "00010000100010101" => rgb <= "000000";
					when "00010000100010110" => rgb <= "000000";
					when "00010000100010111" => rgb <= "000000";
					when "00010000100011000" => rgb <= "000000";
					when "00010000100011001" => rgb <= "000000";
					when "00010000100011010" => rgb <= "000000";
					when "00010000100011011" => rgb <= "000000";
					when "00010000100011100" => rgb <= "000000";
					when "00010000100011101" => rgb <= "000000";
					when "00010000100011110" => rgb <= "000000";
					when "00010000100011111" => rgb <= "000000";
					when "00010000100100000" => rgb <= "000000";
					when "00010000100100001" => rgb <= "000000";
					when "00010000100100010" => rgb <= "000000";
					when "00010000100100011" => rgb <= "000000";
					when "00010000100100100" => rgb <= "000000";
					when "00010000100100101" => rgb <= "000000";
					when "00010000100100110" => rgb <= "000000";
					when "00010000100100111" => rgb <= "000000";
					when "00010000100101000" => rgb <= "000000";
					when "00010000100101001" => rgb <= "000000";
					when "00010000100101010" => rgb <= "000000";
					when "00010000100101011" => rgb <= "000000";
					when "00010000100101100" => rgb <= "000000";
					when "00010000100101101" => rgb <= "000000";
					when "00010000100101110" => rgb <= "000000";
					when "00010000100101111" => rgb <= "000000";
					when "00010000100110000" => rgb <= "000000";
					when "00010000100110001" => rgb <= "000000";
					when "00010000100110010" => rgb <= "000000";
					when "00010000100110011" => rgb <= "000000";
					when "00010000100110100" => rgb <= "000000";
					when "00010000100110101" => rgb <= "000000";
					when "00010000100110110" => rgb <= "000000";
					when "00010000100110111" => rgb <= "000000";
					when "00010000100111000" => rgb <= "000000";
					when "00010000100111001" => rgb <= "000000";
					when "00010000100111010" => rgb <= "000000";
					when "00010000100111011" => rgb <= "000000";
					when "00010000100111100" => rgb <= "000000";
					when "00010000100111101" => rgb <= "000000";
					when "00010000100111110" => rgb <= "000000";
					when "00010000100111111" => rgb <= "000000";
					when "00010001000000000" => rgb <= "000000";
					when "00010001000000001" => rgb <= "000000";
					when "00010001000000010" => rgb <= "000000";
					when "00010001000000011" => rgb <= "000000";
					when "00010001000000100" => rgb <= "000000";
					when "00010001000000101" => rgb <= "000000";
					when "00010001000000110" => rgb <= "000000";
					when "00010001000000111" => rgb <= "000000";
					when "00010001000001000" => rgb <= "000000";
					when "00010001000001001" => rgb <= "000000";
					when "00010001000001010" => rgb <= "000000";
					when "00010001000001011" => rgb <= "000000";
					when "00010001000001100" => rgb <= "000000";
					when "00010001000001101" => rgb <= "000000";
					when "00010001000001110" => rgb <= "000000";
					when "00010001000001111" => rgb <= "000000";
					when "00010001000010000" => rgb <= "000000";
					when "00010001000010001" => rgb <= "000000";
					when "00010001000010010" => rgb <= "000000";
					when "00010001000010011" => rgb <= "000000";
					when "00010001000010100" => rgb <= "000000";
					when "00010001000010101" => rgb <= "000000";
					when "00010001000010110" => rgb <= "000000";
					when "00010001000010111" => rgb <= "000000";
					when "00010001000011000" => rgb <= "000000";
					when "00010001000011001" => rgb <= "000000";
					when "00010001000011010" => rgb <= "000000";
					when "00010001000011011" => rgb <= "000000";
					when "00010001000011100" => rgb <= "000000";
					when "00010001000011101" => rgb <= "000000";
					when "00010001000011110" => rgb <= "000000";
					when "00010001000011111" => rgb <= "000000";
					when "00010001000100000" => rgb <= "000000";
					when "00010001000100001" => rgb <= "000000";
					when "00010001000100010" => rgb <= "000000";
					when "00010001000100011" => rgb <= "000000";
					when "00010001000100100" => rgb <= "000000";
					when "00010001000100101" => rgb <= "000000";
					when "00010001000100110" => rgb <= "000000";
					when "00010001000100111" => rgb <= "000000";
					when "00010001000101000" => rgb <= "000000";
					when "00010001000101001" => rgb <= "000000";
					when "00010001000101010" => rgb <= "000000";
					when "00010001000101011" => rgb <= "000000";
					when "00010001000101100" => rgb <= "000000";
					when "00010001000101101" => rgb <= "000000";
					when "00010001000101110" => rgb <= "000000";
					when "00010001000101111" => rgb <= "000000";
					when "00010001000110000" => rgb <= "000000";
					when "00010001000110001" => rgb <= "000000";
					when "00010001000110010" => rgb <= "000000";
					when "00010001000110011" => rgb <= "000000";
					when "00010001000110100" => rgb <= "000000";
					when "00010001000110101" => rgb <= "000000";
					when "00010001000110110" => rgb <= "000000";
					when "00010001000110111" => rgb <= "000000";
					when "00010001000111000" => rgb <= "000000";
					when "00010001000111001" => rgb <= "000000";
					when "00010001000111010" => rgb <= "000000";
					when "00010001000111011" => rgb <= "000000";
					when "00010001000111100" => rgb <= "000000";
					when "00010001000111101" => rgb <= "000000";
					when "00010001000111110" => rgb <= "000000";
					when "00010001000111111" => rgb <= "000000";
					when "00010001001000000" => rgb <= "000000";
					when "00010001001000001" => rgb <= "000000";
					when "00010001001000010" => rgb <= "000000";
					when "00010001001000011" => rgb <= "000000";
					when "00010001001000100" => rgb <= "000000";
					when "00010001001000101" => rgb <= "000000";
					when "00010001001000110" => rgb <= "000000";
					when "00010001001000111" => rgb <= "000000";
					when "00010001001001000" => rgb <= "000000";
					when "00010001001001001" => rgb <= "000000";
					when "00010001001001010" => rgb <= "000000";
					when "00010001001001011" => rgb <= "000000";
					when "00010001001001100" => rgb <= "000000";
					when "00010001001001101" => rgb <= "000000";
					when "00010001001001110" => rgb <= "000000";
					when "00010001001001111" => rgb <= "000000";
					when "00010001001010000" => rgb <= "000000";
					when "00010001001010001" => rgb <= "000000";
					when "00010001001010010" => rgb <= "000000";
					when "00010001001010011" => rgb <= "000000";
					when "00010001001010100" => rgb <= "000000";
					when "00010001001010101" => rgb <= "000000";
					when "00010001001010110" => rgb <= "000000";
					when "00010001001010111" => rgb <= "000000";
					when "00010001001011000" => rgb <= "000000";
					when "00010001001011001" => rgb <= "000000";
					when "00010001001011010" => rgb <= "000000";
					when "00010001001011011" => rgb <= "000000";
					when "00010001001011100" => rgb <= "000000";
					when "00010001001011101" => rgb <= "000000";
					when "00010001001011110" => rgb <= "000000";
					when "00010001001011111" => rgb <= "000000";
					when "00010001001100000" => rgb <= "000000";
					when "00010001001100001" => rgb <= "000000";
					when "00010001001100010" => rgb <= "000000";
					when "00010001001100011" => rgb <= "000000";
					when "00010001001100100" => rgb <= "000000";
					when "00010001001100101" => rgb <= "000000";
					when "00010001001100110" => rgb <= "000000";
					when "00010001001100111" => rgb <= "000000";
					when "00010001001101000" => rgb <= "000000";
					when "00010001001101001" => rgb <= "000000";
					when "00010001001101010" => rgb <= "000000";
					when "00010001001101011" => rgb <= "000000";
					when "00010001001101100" => rgb <= "000000";
					when "00010001001101101" => rgb <= "000000";
					when "00010001001101110" => rgb <= "000000";
					when "00010001001101111" => rgb <= "000000";
					when "00010001001110000" => rgb <= "000000";
					when "00010001001110001" => rgb <= "000000";
					when "00010001001110010" => rgb <= "000000";
					when "00010001001110011" => rgb <= "000000";
					when "00010001001110100" => rgb <= "000000";
					when "00010001001110101" => rgb <= "000000";
					when "00010001001110110" => rgb <= "000000";
					when "00010001001110111" => rgb <= "000000";
					when "00010001001111000" => rgb <= "000000";
					when "00010001001111001" => rgb <= "000000";
					when "00010001001111010" => rgb <= "000000";
					when "00010001001111011" => rgb <= "000000";
					when "00010001001111100" => rgb <= "000000";
					when "00010001001111101" => rgb <= "100100";
					when "00010001001111110" => rgb <= "101000";
					when "00010001001111111" => rgb <= "101000";
					when "00010001010000000" => rgb <= "101000";
					when "00010001010000001" => rgb <= "101000";
					when "00010001010000010" => rgb <= "101000";
					when "00010001010000011" => rgb <= "101000";
					when "00010001010000100" => rgb <= "101000";
					when "00010001010000101" => rgb <= "101000";
					when "00010001010000110" => rgb <= "101000";
					when "00010001010000111" => rgb <= "101000";
					when "00010001010001000" => rgb <= "101000";
					when "00010001010001001" => rgb <= "101000";
					when "00010001010001010" => rgb <= "101000";
					when "00010001010001011" => rgb <= "101000";
					when "00010001010001100" => rgb <= "101000";
					when "00010001010001101" => rgb <= "101000";
					when "00010001010001110" => rgb <= "101000";
					when "00010001010001111" => rgb <= "101000";
					when "00010001010010000" => rgb <= "101000";
					when "00010001010010001" => rgb <= "101000";
					when "00010001010010010" => rgb <= "101000";
					when "00010001010010011" => rgb <= "101000";
					when "00010001010010100" => rgb <= "101000";
					when "00010001010010101" => rgb <= "101000";
					when "00010001010010110" => rgb <= "101000";
					when "00010001010010111" => rgb <= "101000";
					when "00010001010011000" => rgb <= "101000";
					when "00010001010011001" => rgb <= "101000";
					when "00010001010011010" => rgb <= "101000";
					when "00010001010011011" => rgb <= "101000";
					when "00010001010011100" => rgb <= "101000";
					when "00010001010011101" => rgb <= "101000";
					when "00010001010011110" => rgb <= "101000";
					when "00010001010011111" => rgb <= "101000";
					when "00010001010100000" => rgb <= "101000";
					when "00010001010100001" => rgb <= "101000";
					when "00010001010100010" => rgb <= "101000";
					when "00010001010100011" => rgb <= "101000";
					when "00010001010100100" => rgb <= "101000";
					when "00010001010100101" => rgb <= "101000";
					when "00010001010100110" => rgb <= "101000";
					when "00010001010100111" => rgb <= "101000";
					when "00010001010101000" => rgb <= "101000";
					when "00010001010101001" => rgb <= "101000";
					when "00010001010101010" => rgb <= "101000";
					when "00010001010101011" => rgb <= "101000";
					when "00010001010101100" => rgb <= "101000";
					when "00010001010101101" => rgb <= "101000";
					when "00010001010101110" => rgb <= "101000";
					when "00010001010101111" => rgb <= "101000";
					when "00010001010110000" => rgb <= "101000";
					when "00010001010110001" => rgb <= "101000";
					when "00010001010110010" => rgb <= "101000";
					when "00010001010110011" => rgb <= "101000";
					when "00010001010110100" => rgb <= "101000";
					when "00010001010110101" => rgb <= "101000";
					when "00010001010110110" => rgb <= "100100";
					when "00010001010110111" => rgb <= "100100";
					when "00010001010111000" => rgb <= "100100";
					when "00010001010111001" => rgb <= "100100";
					when "00010001010111010" => rgb <= "100100";
					when "00010001010111011" => rgb <= "100100";
					when "00010001010111100" => rgb <= "100100";
					when "00010001010111101" => rgb <= "100100";
					when "00010001010111110" => rgb <= "100100";
					when "00010001010111111" => rgb <= "100100";
					when "00010001011000000" => rgb <= "010100";
					when "00010001011000001" => rgb <= "000000";
					when "00010001011000010" => rgb <= "000000";
					when "00010001011000011" => rgb <= "000000";
					when "00010001011000100" => rgb <= "000000";
					when "00010001011000101" => rgb <= "000000";
					when "00010001011000110" => rgb <= "000000";
					when "00010001011000111" => rgb <= "000000";
					when "00010001011001000" => rgb <= "000000";
					when "00010001011001001" => rgb <= "000000";
					when "00010001011001010" => rgb <= "000000";
					when "00010001011001011" => rgb <= "000000";
					when "00010001011001100" => rgb <= "000000";
					when "00010001011001101" => rgb <= "000000";
					when "00010001011001110" => rgb <= "000000";
					when "00010001011001111" => rgb <= "000000";
					when "00010001011010000" => rgb <= "000000";
					when "00010001011010001" => rgb <= "000000";
					when "00010001011010010" => rgb <= "000000";
					when "00010001011010011" => rgb <= "000000";
					when "00010001011010100" => rgb <= "000000";
					when "00010001011010101" => rgb <= "000000";
					when "00010001011010110" => rgb <= "000000";
					when "00010001011010111" => rgb <= "000000";
					when "00010001011011000" => rgb <= "000000";
					when "00010001011011001" => rgb <= "000000";
					when "00010001011011010" => rgb <= "000000";
					when "00010001011011011" => rgb <= "000000";
					when "00010001011011100" => rgb <= "000000";
					when "00010001011011101" => rgb <= "000000";
					when "00010001011011110" => rgb <= "000000";
					when "00010001011011111" => rgb <= "000000";
					when "00010001011100000" => rgb <= "000000";
					when "00010001011100001" => rgb <= "000000";
					when "00010001011100010" => rgb <= "000000";
					when "00010001011100011" => rgb <= "000000";
					when "00010001011100100" => rgb <= "000000";
					when "00010001011100101" => rgb <= "000000";
					when "00010001011100110" => rgb <= "000000";
					when "00010001011100111" => rgb <= "000000";
					when "00010001011101000" => rgb <= "000000";
					when "00010001011101001" => rgb <= "000000";
					when "00010001011101010" => rgb <= "000000";
					when "00010001011101011" => rgb <= "000000";
					when "00010001011101100" => rgb <= "000000";
					when "00010001011101101" => rgb <= "000000";
					when "00010001011101110" => rgb <= "000000";
					when "00010001011101111" => rgb <= "000000";
					when "00010001011110000" => rgb <= "000000";
					when "00010001011110001" => rgb <= "000000";
					when "00010001011110010" => rgb <= "000000";
					when "00010001011110011" => rgb <= "000000";
					when "00010001011110100" => rgb <= "000000";
					when "00010001011110101" => rgb <= "000000";
					when "00010001011110110" => rgb <= "000000";
					when "00010001011110111" => rgb <= "000000";
					when "00010001011111000" => rgb <= "000000";
					when "00010001011111001" => rgb <= "000000";
					when "00010001011111010" => rgb <= "000000";
					when "00010001011111011" => rgb <= "000000";
					when "00010001011111100" => rgb <= "000000";
					when "00010001011111101" => rgb <= "000000";
					when "00010001011111110" => rgb <= "000000";
					when "00010001011111111" => rgb <= "000000";
					when "00010001100000000" => rgb <= "000000";
					when "00010001100000001" => rgb <= "000000";
					when "00010001100000010" => rgb <= "000000";
					when "00010001100000011" => rgb <= "000000";
					when "00010001100000100" => rgb <= "000000";
					when "00010001100000101" => rgb <= "000000";
					when "00010001100000110" => rgb <= "000000";
					when "00010001100000111" => rgb <= "000000";
					when "00010001100001000" => rgb <= "000000";
					when "00010001100001001" => rgb <= "000000";
					when "00010001100001010" => rgb <= "000000";
					when "00010001100001011" => rgb <= "000000";
					when "00010001100001100" => rgb <= "000000";
					when "00010001100001101" => rgb <= "000000";
					when "00010001100001110" => rgb <= "000000";
					when "00010001100001111" => rgb <= "000000";
					when "00010001100010000" => rgb <= "000000";
					when "00010001100010001" => rgb <= "000000";
					when "00010001100010010" => rgb <= "000000";
					when "00010001100010011" => rgb <= "000000";
					when "00010001100010100" => rgb <= "000000";
					when "00010001100010101" => rgb <= "000000";
					when "00010001100010110" => rgb <= "000000";
					when "00010001100010111" => rgb <= "000000";
					when "00010001100011000" => rgb <= "000000";
					when "00010001100011001" => rgb <= "000000";
					when "00010001100011010" => rgb <= "000000";
					when "00010001100011011" => rgb <= "000000";
					when "00010001100011100" => rgb <= "000000";
					when "00010001100011101" => rgb <= "000000";
					when "00010001100011110" => rgb <= "000000";
					when "00010001100011111" => rgb <= "000000";
					when "00010001100100000" => rgb <= "000000";
					when "00010001100100001" => rgb <= "000000";
					when "00010001100100010" => rgb <= "000000";
					when "00010001100100011" => rgb <= "000000";
					when "00010001100100100" => rgb <= "000000";
					when "00010001100100101" => rgb <= "000000";
					when "00010001100100110" => rgb <= "000000";
					when "00010001100100111" => rgb <= "000000";
					when "00010001100101000" => rgb <= "000000";
					when "00010001100101001" => rgb <= "000000";
					when "00010001100101010" => rgb <= "000000";
					when "00010001100101011" => rgb <= "000000";
					when "00010001100101100" => rgb <= "000000";
					when "00010001100101101" => rgb <= "000000";
					when "00010001100101110" => rgb <= "000000";
					when "00010001100101111" => rgb <= "000000";
					when "00010001100110000" => rgb <= "000000";
					when "00010001100110001" => rgb <= "000000";
					when "00010001100110010" => rgb <= "000000";
					when "00010001100110011" => rgb <= "000000";
					when "00010001100110100" => rgb <= "000000";
					when "00010001100110101" => rgb <= "000000";
					when "00010001100110110" => rgb <= "000000";
					when "00010001100110111" => rgb <= "000000";
					when "00010001100111000" => rgb <= "000000";
					when "00010001100111001" => rgb <= "000000";
					when "00010001100111010" => rgb <= "000000";
					when "00010001100111011" => rgb <= "000000";
					when "00010001100111100" => rgb <= "000000";
					when "00010001100111101" => rgb <= "000000";
					when "00010001100111110" => rgb <= "000000";
					when "00010001100111111" => rgb <= "000000";
					when "00010010000000000" => rgb <= "000000";
					when "00010010000000001" => rgb <= "000000";
					when "00010010000000010" => rgb <= "000000";
					when "00010010000000011" => rgb <= "000000";
					when "00010010000000100" => rgb <= "000000";
					when "00010010000000101" => rgb <= "000000";
					when "00010010000000110" => rgb <= "000000";
					when "00010010000000111" => rgb <= "000000";
					when "00010010000001000" => rgb <= "000000";
					when "00010010000001001" => rgb <= "000000";
					when "00010010000001010" => rgb <= "000000";
					when "00010010000001011" => rgb <= "000000";
					when "00010010000001100" => rgb <= "000000";
					when "00010010000001101" => rgb <= "000000";
					when "00010010000001110" => rgb <= "000000";
					when "00010010000001111" => rgb <= "000000";
					when "00010010000010000" => rgb <= "000000";
					when "00010010000010001" => rgb <= "000000";
					when "00010010000010010" => rgb <= "000000";
					when "00010010000010011" => rgb <= "000000";
					when "00010010000010100" => rgb <= "000000";
					when "00010010000010101" => rgb <= "000000";
					when "00010010000010110" => rgb <= "000000";
					when "00010010000010111" => rgb <= "000000";
					when "00010010000011000" => rgb <= "000000";
					when "00010010000011001" => rgb <= "000000";
					when "00010010000011010" => rgb <= "000000";
					when "00010010000011011" => rgb <= "000000";
					when "00010010000011100" => rgb <= "000000";
					when "00010010000011101" => rgb <= "000000";
					when "00010010000011110" => rgb <= "000000";
					when "00010010000011111" => rgb <= "000000";
					when "00010010000100000" => rgb <= "000000";
					when "00010010000100001" => rgb <= "000000";
					when "00010010000100010" => rgb <= "000000";
					when "00010010000100011" => rgb <= "000000";
					when "00010010000100100" => rgb <= "000000";
					when "00010010000100101" => rgb <= "000000";
					when "00010010000100110" => rgb <= "000000";
					when "00010010000100111" => rgb <= "000000";
					when "00010010000101000" => rgb <= "000000";
					when "00010010000101001" => rgb <= "000000";
					when "00010010000101010" => rgb <= "000000";
					when "00010010000101011" => rgb <= "000000";
					when "00010010000101100" => rgb <= "000000";
					when "00010010000101101" => rgb <= "000000";
					when "00010010000101110" => rgb <= "000000";
					when "00010010000101111" => rgb <= "000000";
					when "00010010000110000" => rgb <= "000000";
					when "00010010000110001" => rgb <= "000000";
					when "00010010000110010" => rgb <= "000000";
					when "00010010000110011" => rgb <= "000000";
					when "00010010000110100" => rgb <= "000000";
					when "00010010000110101" => rgb <= "000000";
					when "00010010000110110" => rgb <= "000000";
					when "00010010000110111" => rgb <= "000000";
					when "00010010000111000" => rgb <= "000000";
					when "00010010000111001" => rgb <= "000000";
					when "00010010000111010" => rgb <= "000000";
					when "00010010000111011" => rgb <= "000000";
					when "00010010000111100" => rgb <= "000000";
					when "00010010000111101" => rgb <= "000000";
					when "00010010000111110" => rgb <= "000000";
					when "00010010000111111" => rgb <= "000000";
					when "00010010001000000" => rgb <= "000000";
					when "00010010001000001" => rgb <= "000000";
					when "00010010001000010" => rgb <= "000000";
					when "00010010001000011" => rgb <= "000000";
					when "00010010001000100" => rgb <= "000000";
					when "00010010001000101" => rgb <= "000000";
					when "00010010001000110" => rgb <= "000000";
					when "00010010001000111" => rgb <= "000000";
					when "00010010001001000" => rgb <= "000000";
					when "00010010001001001" => rgb <= "000000";
					when "00010010001001010" => rgb <= "000000";
					when "00010010001001011" => rgb <= "000000";
					when "00010010001001100" => rgb <= "000000";
					when "00010010001001101" => rgb <= "000000";
					when "00010010001001110" => rgb <= "000000";
					when "00010010001001111" => rgb <= "000000";
					when "00010010001010000" => rgb <= "000000";
					when "00010010001010001" => rgb <= "000000";
					when "00010010001010010" => rgb <= "000000";
					when "00010010001010011" => rgb <= "000000";
					when "00010010001010100" => rgb <= "000000";
					when "00010010001010101" => rgb <= "000000";
					when "00010010001010110" => rgb <= "000000";
					when "00010010001010111" => rgb <= "000000";
					when "00010010001011000" => rgb <= "000000";
					when "00010010001011001" => rgb <= "000000";
					when "00010010001011010" => rgb <= "000000";
					when "00010010001011011" => rgb <= "000000";
					when "00010010001011100" => rgb <= "000000";
					when "00010010001011101" => rgb <= "000000";
					when "00010010001011110" => rgb <= "000000";
					when "00010010001011111" => rgb <= "000000";
					when "00010010001100000" => rgb <= "000000";
					when "00010010001100001" => rgb <= "000000";
					when "00010010001100010" => rgb <= "000000";
					when "00010010001100011" => rgb <= "000000";
					when "00010010001100100" => rgb <= "000000";
					when "00010010001100101" => rgb <= "000000";
					when "00010010001100110" => rgb <= "000000";
					when "00010010001100111" => rgb <= "000000";
					when "00010010001101000" => rgb <= "000000";
					when "00010010001101001" => rgb <= "000000";
					when "00010010001101010" => rgb <= "000000";
					when "00010010001101011" => rgb <= "000000";
					when "00010010001101100" => rgb <= "000000";
					when "00010010001101101" => rgb <= "000000";
					when "00010010001101110" => rgb <= "000000";
					when "00010010001101111" => rgb <= "000000";
					when "00010010001110000" => rgb <= "000000";
					when "00010010001110001" => rgb <= "000000";
					when "00010010001110010" => rgb <= "000000";
					when "00010010001110011" => rgb <= "000000";
					when "00010010001110100" => rgb <= "000000";
					when "00010010001110101" => rgb <= "000000";
					when "00010010001110110" => rgb <= "000000";
					when "00010010001110111" => rgb <= "000000";
					when "00010010001111000" => rgb <= "000000";
					when "00010010001111001" => rgb <= "000000";
					when "00010010001111010" => rgb <= "000000";
					when "00010010001111011" => rgb <= "000000";
					when "00010010001111100" => rgb <= "000000";
					when "00010010001111101" => rgb <= "101000";
					when "00010010001111110" => rgb <= "101000";
					when "00010010001111111" => rgb <= "101000";
					when "00010010010000000" => rgb <= "101000";
					when "00010010010000001" => rgb <= "101000";
					when "00010010010000010" => rgb <= "101000";
					when "00010010010000011" => rgb <= "101000";
					when "00010010010000100" => rgb <= "101000";
					when "00010010010000101" => rgb <= "101000";
					when "00010010010000110" => rgb <= "101000";
					when "00010010010000111" => rgb <= "101000";
					when "00010010010001000" => rgb <= "101000";
					when "00010010010001001" => rgb <= "101000";
					when "00010010010001010" => rgb <= "101000";
					when "00010010010001011" => rgb <= "101000";
					when "00010010010001100" => rgb <= "101000";
					when "00010010010001101" => rgb <= "101000";
					when "00010010010001110" => rgb <= "101000";
					when "00010010010001111" => rgb <= "101000";
					when "00010010010010000" => rgb <= "101000";
					when "00010010010010001" => rgb <= "101000";
					when "00010010010010010" => rgb <= "101000";
					when "00010010010010011" => rgb <= "101000";
					when "00010010010010100" => rgb <= "101000";
					when "00010010010010101" => rgb <= "101000";
					when "00010010010010110" => rgb <= "101000";
					when "00010010010010111" => rgb <= "101000";
					when "00010010010011000" => rgb <= "101000";
					when "00010010010011001" => rgb <= "101000";
					when "00010010010011010" => rgb <= "101000";
					when "00010010010011011" => rgb <= "101000";
					when "00010010010011100" => rgb <= "101000";
					when "00010010010011101" => rgb <= "101000";
					when "00010010010011110" => rgb <= "101000";
					when "00010010010011111" => rgb <= "101000";
					when "00010010010100000" => rgb <= "101000";
					when "00010010010100001" => rgb <= "101000";
					when "00010010010100010" => rgb <= "101000";
					when "00010010010100011" => rgb <= "101000";
					when "00010010010100100" => rgb <= "101000";
					when "00010010010100101" => rgb <= "101000";
					when "00010010010100110" => rgb <= "101000";
					when "00010010010100111" => rgb <= "101000";
					when "00010010010101000" => rgb <= "101000";
					when "00010010010101001" => rgb <= "101000";
					when "00010010010101010" => rgb <= "101000";
					when "00010010010101011" => rgb <= "101000";
					when "00010010010101100" => rgb <= "101000";
					when "00010010010101101" => rgb <= "101000";
					when "00010010010101110" => rgb <= "101000";
					when "00010010010101111" => rgb <= "101000";
					when "00010010010110000" => rgb <= "101000";
					when "00010010010110001" => rgb <= "101000";
					when "00010010010110010" => rgb <= "111000";
					when "00010010010110011" => rgb <= "101000";
					when "00010010010110100" => rgb <= "101000";
					when "00010010010110101" => rgb <= "101000";
					when "00010010010110110" => rgb <= "101000";
					when "00010010010110111" => rgb <= "101000";
					when "00010010010111000" => rgb <= "101000";
					when "00010010010111001" => rgb <= "101000";
					when "00010010010111010" => rgb <= "101000";
					when "00010010010111011" => rgb <= "101000";
					when "00010010010111100" => rgb <= "101000";
					when "00010010010111101" => rgb <= "101000";
					when "00010010010111110" => rgb <= "101000";
					when "00010010010111111" => rgb <= "101000";
					when "00010010011000000" => rgb <= "101000";
					when "00010010011000001" => rgb <= "000000";
					when "00010010011000010" => rgb <= "000000";
					when "00010010011000011" => rgb <= "000000";
					when "00010010011000100" => rgb <= "000000";
					when "00010010011000101" => rgb <= "000000";
					when "00010010011000110" => rgb <= "000000";
					when "00010010011000111" => rgb <= "000000";
					when "00010010011001000" => rgb <= "000000";
					when "00010010011001001" => rgb <= "000000";
					when "00010010011001010" => rgb <= "000000";
					when "00010010011001011" => rgb <= "000000";
					when "00010010011001100" => rgb <= "000000";
					when "00010010011001101" => rgb <= "000000";
					when "00010010011001110" => rgb <= "000000";
					when "00010010011001111" => rgb <= "000000";
					when "00010010011010000" => rgb <= "000000";
					when "00010010011010001" => rgb <= "000000";
					when "00010010011010010" => rgb <= "000000";
					when "00010010011010011" => rgb <= "000000";
					when "00010010011010100" => rgb <= "000000";
					when "00010010011010101" => rgb <= "000000";
					when "00010010011010110" => rgb <= "000000";
					when "00010010011010111" => rgb <= "000000";
					when "00010010011011000" => rgb <= "000000";
					when "00010010011011001" => rgb <= "000000";
					when "00010010011011010" => rgb <= "000000";
					when "00010010011011011" => rgb <= "000000";
					when "00010010011011100" => rgb <= "000000";
					when "00010010011011101" => rgb <= "000000";
					when "00010010011011110" => rgb <= "000000";
					when "00010010011011111" => rgb <= "000000";
					when "00010010011100000" => rgb <= "000000";
					when "00010010011100001" => rgb <= "000000";
					when "00010010011100010" => rgb <= "000000";
					when "00010010011100011" => rgb <= "000000";
					when "00010010011100100" => rgb <= "000000";
					when "00010010011100101" => rgb <= "000000";
					when "00010010011100110" => rgb <= "000000";
					when "00010010011100111" => rgb <= "000000";
					when "00010010011101000" => rgb <= "000000";
					when "00010010011101001" => rgb <= "000000";
					when "00010010011101010" => rgb <= "000000";
					when "00010010011101011" => rgb <= "000000";
					when "00010010011101100" => rgb <= "000000";
					when "00010010011101101" => rgb <= "000000";
					when "00010010011101110" => rgb <= "000000";
					when "00010010011101111" => rgb <= "000000";
					when "00010010011110000" => rgb <= "000000";
					when "00010010011110001" => rgb <= "000000";
					when "00010010011110010" => rgb <= "000000";
					when "00010010011110011" => rgb <= "000000";
					when "00010010011110100" => rgb <= "000000";
					when "00010010011110101" => rgb <= "000000";
					when "00010010011110110" => rgb <= "000000";
					when "00010010011110111" => rgb <= "000000";
					when "00010010011111000" => rgb <= "000000";
					when "00010010011111001" => rgb <= "000000";
					when "00010010011111010" => rgb <= "000000";
					when "00010010011111011" => rgb <= "000000";
					when "00010010011111100" => rgb <= "000000";
					when "00010010011111101" => rgb <= "000000";
					when "00010010011111110" => rgb <= "000000";
					when "00010010011111111" => rgb <= "000000";
					when "00010010100000000" => rgb <= "000000";
					when "00010010100000001" => rgb <= "000000";
					when "00010010100000010" => rgb <= "000000";
					when "00010010100000011" => rgb <= "000000";
					when "00010010100000100" => rgb <= "000000";
					when "00010010100000101" => rgb <= "000000";
					when "00010010100000110" => rgb <= "000000";
					when "00010010100000111" => rgb <= "000000";
					when "00010010100001000" => rgb <= "000000";
					when "00010010100001001" => rgb <= "000000";
					when "00010010100001010" => rgb <= "000000";
					when "00010010100001011" => rgb <= "000000";
					when "00010010100001100" => rgb <= "000000";
					when "00010010100001101" => rgb <= "000000";
					when "00010010100001110" => rgb <= "000000";
					when "00010010100001111" => rgb <= "000000";
					when "00010010100010000" => rgb <= "000000";
					when "00010010100010001" => rgb <= "000000";
					when "00010010100010010" => rgb <= "000000";
					when "00010010100010011" => rgb <= "000000";
					when "00010010100010100" => rgb <= "000000";
					when "00010010100010101" => rgb <= "000000";
					when "00010010100010110" => rgb <= "000000";
					when "00010010100010111" => rgb <= "000000";
					when "00010010100011000" => rgb <= "000000";
					when "00010010100011001" => rgb <= "000000";
					when "00010010100011010" => rgb <= "000000";
					when "00010010100011011" => rgb <= "000000";
					when "00010010100011100" => rgb <= "000000";
					when "00010010100011101" => rgb <= "000000";
					when "00010010100011110" => rgb <= "000000";
					when "00010010100011111" => rgb <= "000000";
					when "00010010100100000" => rgb <= "000000";
					when "00010010100100001" => rgb <= "000000";
					when "00010010100100010" => rgb <= "000000";
					when "00010010100100011" => rgb <= "000000";
					when "00010010100100100" => rgb <= "000000";
					when "00010010100100101" => rgb <= "000000";
					when "00010010100100110" => rgb <= "000000";
					when "00010010100100111" => rgb <= "000000";
					when "00010010100101000" => rgb <= "000000";
					when "00010010100101001" => rgb <= "000000";
					when "00010010100101010" => rgb <= "000000";
					when "00010010100101011" => rgb <= "000000";
					when "00010010100101100" => rgb <= "000000";
					when "00010010100101101" => rgb <= "000000";
					when "00010010100101110" => rgb <= "000000";
					when "00010010100101111" => rgb <= "000000";
					when "00010010100110000" => rgb <= "000000";
					when "00010010100110001" => rgb <= "000000";
					when "00010010100110010" => rgb <= "000000";
					when "00010010100110011" => rgb <= "000000";
					when "00010010100110100" => rgb <= "000000";
					when "00010010100110101" => rgb <= "000000";
					when "00010010100110110" => rgb <= "000000";
					when "00010010100110111" => rgb <= "000000";
					when "00010010100111000" => rgb <= "000000";
					when "00010010100111001" => rgb <= "000000";
					when "00010010100111010" => rgb <= "000000";
					when "00010010100111011" => rgb <= "000000";
					when "00010010100111100" => rgb <= "000000";
					when "00010010100111101" => rgb <= "000000";
					when "00010010100111110" => rgb <= "000000";
					when "00010010100111111" => rgb <= "000000";
					when "00010011000000000" => rgb <= "000000";
					when "00010011000000001" => rgb <= "000000";
					when "00010011000000010" => rgb <= "000000";
					when "00010011000000011" => rgb <= "000000";
					when "00010011000000100" => rgb <= "000000";
					when "00010011000000101" => rgb <= "000000";
					when "00010011000000110" => rgb <= "000000";
					when "00010011000000111" => rgb <= "000000";
					when "00010011000001000" => rgb <= "000000";
					when "00010011000001001" => rgb <= "000000";
					when "00010011000001010" => rgb <= "000000";
					when "00010011000001011" => rgb <= "000000";
					when "00010011000001100" => rgb <= "000000";
					when "00010011000001101" => rgb <= "000000";
					when "00010011000001110" => rgb <= "000000";
					when "00010011000001111" => rgb <= "000000";
					when "00010011000010000" => rgb <= "000000";
					when "00010011000010001" => rgb <= "000000";
					when "00010011000010010" => rgb <= "000000";
					when "00010011000010011" => rgb <= "000000";
					when "00010011000010100" => rgb <= "000000";
					when "00010011000010101" => rgb <= "000000";
					when "00010011000010110" => rgb <= "000000";
					when "00010011000010111" => rgb <= "000000";
					when "00010011000011000" => rgb <= "000000";
					when "00010011000011001" => rgb <= "000000";
					when "00010011000011010" => rgb <= "000000";
					when "00010011000011011" => rgb <= "000000";
					when "00010011000011100" => rgb <= "000000";
					when "00010011000011101" => rgb <= "000000";
					when "00010011000011110" => rgb <= "000000";
					when "00010011000011111" => rgb <= "000000";
					when "00010011000100000" => rgb <= "000000";
					when "00010011000100001" => rgb <= "000000";
					when "00010011000100010" => rgb <= "000000";
					when "00010011000100011" => rgb <= "000000";
					when "00010011000100100" => rgb <= "000000";
					when "00010011000100101" => rgb <= "000000";
					when "00010011000100110" => rgb <= "000000";
					when "00010011000100111" => rgb <= "000000";
					when "00010011000101000" => rgb <= "000000";
					when "00010011000101001" => rgb <= "000000";
					when "00010011000101010" => rgb <= "000000";
					when "00010011000101011" => rgb <= "000000";
					when "00010011000101100" => rgb <= "000000";
					when "00010011000101101" => rgb <= "000000";
					when "00010011000101110" => rgb <= "000000";
					when "00010011000101111" => rgb <= "000000";
					when "00010011000110000" => rgb <= "000000";
					when "00010011000110001" => rgb <= "000000";
					when "00010011000110010" => rgb <= "000000";
					when "00010011000110011" => rgb <= "000000";
					when "00010011000110100" => rgb <= "000000";
					when "00010011000110101" => rgb <= "000000";
					when "00010011000110110" => rgb <= "000000";
					when "00010011000110111" => rgb <= "000000";
					when "00010011000111000" => rgb <= "000000";
					when "00010011000111001" => rgb <= "000000";
					when "00010011000111010" => rgb <= "000000";
					when "00010011000111011" => rgb <= "000000";
					when "00010011000111100" => rgb <= "000000";
					when "00010011000111101" => rgb <= "000000";
					when "00010011000111110" => rgb <= "000000";
					when "00010011000111111" => rgb <= "000000";
					when "00010011001000000" => rgb <= "000000";
					when "00010011001000001" => rgb <= "000000";
					when "00010011001000010" => rgb <= "000000";
					when "00010011001000011" => rgb <= "000000";
					when "00010011001000100" => rgb <= "000000";
					when "00010011001000101" => rgb <= "000000";
					when "00010011001000110" => rgb <= "000000";
					when "00010011001000111" => rgb <= "000000";
					when "00010011001001000" => rgb <= "000000";
					when "00010011001001001" => rgb <= "000000";
					when "00010011001001010" => rgb <= "000000";
					when "00010011001001011" => rgb <= "000000";
					when "00010011001001100" => rgb <= "000000";
					when "00010011001001101" => rgb <= "000000";
					when "00010011001001110" => rgb <= "000000";
					when "00010011001001111" => rgb <= "000000";
					when "00010011001010000" => rgb <= "000000";
					when "00010011001010001" => rgb <= "000000";
					when "00010011001010010" => rgb <= "000000";
					when "00010011001010011" => rgb <= "000000";
					when "00010011001010100" => rgb <= "000000";
					when "00010011001010101" => rgb <= "000000";
					when "00010011001010110" => rgb <= "000000";
					when "00010011001010111" => rgb <= "000000";
					when "00010011001011000" => rgb <= "000000";
					when "00010011001011001" => rgb <= "000000";
					when "00010011001011010" => rgb <= "000000";
					when "00010011001011011" => rgb <= "000000";
					when "00010011001011100" => rgb <= "000000";
					when "00010011001011101" => rgb <= "000000";
					when "00010011001011110" => rgb <= "000000";
					when "00010011001011111" => rgb <= "000000";
					when "00010011001100000" => rgb <= "000000";
					when "00010011001100001" => rgb <= "000000";
					when "00010011001100010" => rgb <= "000000";
					when "00010011001100011" => rgb <= "000000";
					when "00010011001100100" => rgb <= "000000";
					when "00010011001100101" => rgb <= "000000";
					when "00010011001100110" => rgb <= "000000";
					when "00010011001100111" => rgb <= "000000";
					when "00010011001101000" => rgb <= "000000";
					when "00010011001101001" => rgb <= "000000";
					when "00010011001101010" => rgb <= "000000";
					when "00010011001101011" => rgb <= "000000";
					when "00010011001101100" => rgb <= "000000";
					when "00010011001101101" => rgb <= "000000";
					when "00010011001101110" => rgb <= "000000";
					when "00010011001101111" => rgb <= "000000";
					when "00010011001110000" => rgb <= "000000";
					when "00010011001110001" => rgb <= "000000";
					when "00010011001110010" => rgb <= "000000";
					when "00010011001110011" => rgb <= "000000";
					when "00010011001110100" => rgb <= "000000";
					when "00010011001110101" => rgb <= "000000";
					when "00010011001110110" => rgb <= "000000";
					when "00010011001110111" => rgb <= "000000";
					when "00010011001111000" => rgb <= "000000";
					when "00010011001111001" => rgb <= "000000";
					when "00010011001111010" => rgb <= "000000";
					when "00010011001111011" => rgb <= "000000";
					when "00010011001111100" => rgb <= "000000";
					when "00010011001111101" => rgb <= "101000";
					when "00010011001111110" => rgb <= "101000";
					when "00010011001111111" => rgb <= "101000";
					when "00010011010000000" => rgb <= "101000";
					when "00010011010000001" => rgb <= "101000";
					when "00010011010000010" => rgb <= "101000";
					when "00010011010000011" => rgb <= "101000";
					when "00010011010000100" => rgb <= "101000";
					when "00010011010000101" => rgb <= "101000";
					when "00010011010000110" => rgb <= "101000";
					when "00010011010000111" => rgb <= "101000";
					when "00010011010001000" => rgb <= "101000";
					when "00010011010001001" => rgb <= "101000";
					when "00010011010001010" => rgb <= "101000";
					when "00010011010001011" => rgb <= "101000";
					when "00010011010001100" => rgb <= "101000";
					when "00010011010001101" => rgb <= "101000";
					when "00010011010001110" => rgb <= "101000";
					when "00010011010001111" => rgb <= "101000";
					when "00010011010010000" => rgb <= "101000";
					when "00010011010010001" => rgb <= "101000";
					when "00010011010010010" => rgb <= "101000";
					when "00010011010010011" => rgb <= "101000";
					when "00010011010010100" => rgb <= "101000";
					when "00010011010010101" => rgb <= "101000";
					when "00010011010010110" => rgb <= "101000";
					when "00010011010010111" => rgb <= "101000";
					when "00010011010011000" => rgb <= "101000";
					when "00010011010011001" => rgb <= "101000";
					when "00010011010011010" => rgb <= "101000";
					when "00010011010011011" => rgb <= "101000";
					when "00010011010011100" => rgb <= "101000";
					when "00010011010011101" => rgb <= "101000";
					when "00010011010011110" => rgb <= "101000";
					when "00010011010011111" => rgb <= "101000";
					when "00010011010100000" => rgb <= "101000";
					when "00010011010100001" => rgb <= "101000";
					when "00010011010100010" => rgb <= "101000";
					when "00010011010100011" => rgb <= "101000";
					when "00010011010100100" => rgb <= "101000";
					when "00010011010100101" => rgb <= "101000";
					when "00010011010100110" => rgb <= "101000";
					when "00010011010100111" => rgb <= "101000";
					when "00010011010101000" => rgb <= "101000";
					when "00010011010101001" => rgb <= "101000";
					when "00010011010101010" => rgb <= "101000";
					when "00010011010101011" => rgb <= "101000";
					when "00010011010101100" => rgb <= "101000";
					when "00010011010101101" => rgb <= "101000";
					when "00010011010101110" => rgb <= "101000";
					when "00010011010101111" => rgb <= "101000";
					when "00010011010110000" => rgb <= "101000";
					when "00010011010110001" => rgb <= "101000";
					when "00010011010110010" => rgb <= "101000";
					when "00010011010110011" => rgb <= "101000";
					when "00010011010110100" => rgb <= "101000";
					when "00010011010110101" => rgb <= "101000";
					when "00010011010110110" => rgb <= "101000";
					when "00010011010110111" => rgb <= "101000";
					when "00010011010111000" => rgb <= "101000";
					when "00010011010111001" => rgb <= "101000";
					when "00010011010111010" => rgb <= "101000";
					when "00010011010111011" => rgb <= "101000";
					when "00010011010111100" => rgb <= "101000";
					when "00010011010111101" => rgb <= "101000";
					when "00010011010111110" => rgb <= "101000";
					when "00010011010111111" => rgb <= "101000";
					when "00010011011000000" => rgb <= "101000";
					when "00010011011000001" => rgb <= "000000";
					when "00010011011000010" => rgb <= "000000";
					when "00010011011000011" => rgb <= "000000";
					when "00010011011000100" => rgb <= "000000";
					when "00010011011000101" => rgb <= "000000";
					when "00010011011000110" => rgb <= "000000";
					when "00010011011000111" => rgb <= "000000";
					when "00010011011001000" => rgb <= "000000";
					when "00010011011001001" => rgb <= "000000";
					when "00010011011001010" => rgb <= "000000";
					when "00010011011001011" => rgb <= "000000";
					when "00010011011001100" => rgb <= "000000";
					when "00010011011001101" => rgb <= "000000";
					when "00010011011001110" => rgb <= "000000";
					when "00010011011001111" => rgb <= "000000";
					when "00010011011010000" => rgb <= "000000";
					when "00010011011010001" => rgb <= "000000";
					when "00010011011010010" => rgb <= "000000";
					when "00010011011010011" => rgb <= "000000";
					when "00010011011010100" => rgb <= "000000";
					when "00010011011010101" => rgb <= "000000";
					when "00010011011010110" => rgb <= "000000";
					when "00010011011010111" => rgb <= "000000";
					when "00010011011011000" => rgb <= "000000";
					when "00010011011011001" => rgb <= "000000";
					when "00010011011011010" => rgb <= "000000";
					when "00010011011011011" => rgb <= "000000";
					when "00010011011011100" => rgb <= "000000";
					when "00010011011011101" => rgb <= "000000";
					when "00010011011011110" => rgb <= "000000";
					when "00010011011011111" => rgb <= "000000";
					when "00010011011100000" => rgb <= "000000";
					when "00010011011100001" => rgb <= "000000";
					when "00010011011100010" => rgb <= "000000";
					when "00010011011100011" => rgb <= "000000";
					when "00010011011100100" => rgb <= "000000";
					when "00010011011100101" => rgb <= "000000";
					when "00010011011100110" => rgb <= "000000";
					when "00010011011100111" => rgb <= "000000";
					when "00010011011101000" => rgb <= "000000";
					when "00010011011101001" => rgb <= "000000";
					when "00010011011101010" => rgb <= "000000";
					when "00010011011101011" => rgb <= "000000";
					when "00010011011101100" => rgb <= "000000";
					when "00010011011101101" => rgb <= "000000";
					when "00010011011101110" => rgb <= "000000";
					when "00010011011101111" => rgb <= "000000";
					when "00010011011110000" => rgb <= "000000";
					when "00010011011110001" => rgb <= "000000";
					when "00010011011110010" => rgb <= "000000";
					when "00010011011110011" => rgb <= "000000";
					when "00010011011110100" => rgb <= "000000";
					when "00010011011110101" => rgb <= "000000";
					when "00010011011110110" => rgb <= "000000";
					when "00010011011110111" => rgb <= "000000";
					when "00010011011111000" => rgb <= "000000";
					when "00010011011111001" => rgb <= "000000";
					when "00010011011111010" => rgb <= "000000";
					when "00010011011111011" => rgb <= "000000";
					when "00010011011111100" => rgb <= "000000";
					when "00010011011111101" => rgb <= "000000";
					when "00010011011111110" => rgb <= "000000";
					when "00010011011111111" => rgb <= "000000";
					when "00010011100000000" => rgb <= "000000";
					when "00010011100000001" => rgb <= "000000";
					when "00010011100000010" => rgb <= "000000";
					when "00010011100000011" => rgb <= "000000";
					when "00010011100000100" => rgb <= "000000";
					when "00010011100000101" => rgb <= "000000";
					when "00010011100000110" => rgb <= "000000";
					when "00010011100000111" => rgb <= "000000";
					when "00010011100001000" => rgb <= "000000";
					when "00010011100001001" => rgb <= "000000";
					when "00010011100001010" => rgb <= "000000";
					when "00010011100001011" => rgb <= "000000";
					when "00010011100001100" => rgb <= "000000";
					when "00010011100001101" => rgb <= "000000";
					when "00010011100001110" => rgb <= "000000";
					when "00010011100001111" => rgb <= "000000";
					when "00010011100010000" => rgb <= "000000";
					when "00010011100010001" => rgb <= "000000";
					when "00010011100010010" => rgb <= "000000";
					when "00010011100010011" => rgb <= "000000";
					when "00010011100010100" => rgb <= "000000";
					when "00010011100010101" => rgb <= "000000";
					when "00010011100010110" => rgb <= "000000";
					when "00010011100010111" => rgb <= "000000";
					when "00010011100011000" => rgb <= "000000";
					when "00010011100011001" => rgb <= "000000";
					when "00010011100011010" => rgb <= "000000";
					when "00010011100011011" => rgb <= "000000";
					when "00010011100011100" => rgb <= "000000";
					when "00010011100011101" => rgb <= "000000";
					when "00010011100011110" => rgb <= "000000";
					when "00010011100011111" => rgb <= "000000";
					when "00010011100100000" => rgb <= "000000";
					when "00010011100100001" => rgb <= "000000";
					when "00010011100100010" => rgb <= "000000";
					when "00010011100100011" => rgb <= "000000";
					when "00010011100100100" => rgb <= "000000";
					when "00010011100100101" => rgb <= "000000";
					when "00010011100100110" => rgb <= "000000";
					when "00010011100100111" => rgb <= "000000";
					when "00010011100101000" => rgb <= "000000";
					when "00010011100101001" => rgb <= "000000";
					when "00010011100101010" => rgb <= "000000";
					when "00010011100101011" => rgb <= "000000";
					when "00010011100101100" => rgb <= "000000";
					when "00010011100101101" => rgb <= "000000";
					when "00010011100101110" => rgb <= "000000";
					when "00010011100101111" => rgb <= "000000";
					when "00010011100110000" => rgb <= "000000";
					when "00010011100110001" => rgb <= "000000";
					when "00010011100110010" => rgb <= "000000";
					when "00010011100110011" => rgb <= "000000";
					when "00010011100110100" => rgb <= "000000";
					when "00010011100110101" => rgb <= "000000";
					when "00010011100110110" => rgb <= "000000";
					when "00010011100110111" => rgb <= "000000";
					when "00010011100111000" => rgb <= "000000";
					when "00010011100111001" => rgb <= "000000";
					when "00010011100111010" => rgb <= "000000";
					when "00010011100111011" => rgb <= "000000";
					when "00010011100111100" => rgb <= "000000";
					when "00010011100111101" => rgb <= "000000";
					when "00010011100111110" => rgb <= "000000";
					when "00010011100111111" => rgb <= "000000";
					when "00010100000000000" => rgb <= "000000";
					when "00010100000000001" => rgb <= "000000";
					when "00010100000000010" => rgb <= "000000";
					when "00010100000000011" => rgb <= "000000";
					when "00010100000000100" => rgb <= "000000";
					when "00010100000000101" => rgb <= "000000";
					when "00010100000000110" => rgb <= "000000";
					when "00010100000000111" => rgb <= "000000";
					when "00010100000001000" => rgb <= "000000";
					when "00010100000001001" => rgb <= "000000";
					when "00010100000001010" => rgb <= "000000";
					when "00010100000001011" => rgb <= "000000";
					when "00010100000001100" => rgb <= "000000";
					when "00010100000001101" => rgb <= "000000";
					when "00010100000001110" => rgb <= "000000";
					when "00010100000001111" => rgb <= "000000";
					when "00010100000010000" => rgb <= "000000";
					when "00010100000010001" => rgb <= "000000";
					when "00010100000010010" => rgb <= "000000";
					when "00010100000010011" => rgb <= "000000";
					when "00010100000010100" => rgb <= "000000";
					when "00010100000010101" => rgb <= "000000";
					when "00010100000010110" => rgb <= "000000";
					when "00010100000010111" => rgb <= "000000";
					when "00010100000011000" => rgb <= "000000";
					when "00010100000011001" => rgb <= "000000";
					when "00010100000011010" => rgb <= "000000";
					when "00010100000011011" => rgb <= "000000";
					when "00010100000011100" => rgb <= "000000";
					when "00010100000011101" => rgb <= "000000";
					when "00010100000011110" => rgb <= "000000";
					when "00010100000011111" => rgb <= "000000";
					when "00010100000100000" => rgb <= "000000";
					when "00010100000100001" => rgb <= "000000";
					when "00010100000100010" => rgb <= "000000";
					when "00010100000100011" => rgb <= "000000";
					when "00010100000100100" => rgb <= "000000";
					when "00010100000100101" => rgb <= "000000";
					when "00010100000100110" => rgb <= "000000";
					when "00010100000100111" => rgb <= "000000";
					when "00010100000101000" => rgb <= "000000";
					when "00010100000101001" => rgb <= "000000";
					when "00010100000101010" => rgb <= "000000";
					when "00010100000101011" => rgb <= "000000";
					when "00010100000101100" => rgb <= "000000";
					when "00010100000101101" => rgb <= "000000";
					when "00010100000101110" => rgb <= "000000";
					when "00010100000101111" => rgb <= "000000";
					when "00010100000110000" => rgb <= "000000";
					when "00010100000110001" => rgb <= "000000";
					when "00010100000110010" => rgb <= "000000";
					when "00010100000110011" => rgb <= "000000";
					when "00010100000110100" => rgb <= "000000";
					when "00010100000110101" => rgb <= "000000";
					when "00010100000110110" => rgb <= "000000";
					when "00010100000110111" => rgb <= "000000";
					when "00010100000111000" => rgb <= "000000";
					when "00010100000111001" => rgb <= "000000";
					when "00010100000111010" => rgb <= "000000";
					when "00010100000111011" => rgb <= "000000";
					when "00010100000111100" => rgb <= "000000";
					when "00010100000111101" => rgb <= "000000";
					when "00010100000111110" => rgb <= "000000";
					when "00010100000111111" => rgb <= "000000";
					when "00010100001000000" => rgb <= "000000";
					when "00010100001000001" => rgb <= "000000";
					when "00010100001000010" => rgb <= "000000";
					when "00010100001000011" => rgb <= "000000";
					when "00010100001000100" => rgb <= "000000";
					when "00010100001000101" => rgb <= "000000";
					when "00010100001000110" => rgb <= "000000";
					when "00010100001000111" => rgb <= "000000";
					when "00010100001001000" => rgb <= "000000";
					when "00010100001001001" => rgb <= "000000";
					when "00010100001001010" => rgb <= "000000";
					when "00010100001001011" => rgb <= "000000";
					when "00010100001001100" => rgb <= "000000";
					when "00010100001001101" => rgb <= "000000";
					when "00010100001001110" => rgb <= "000000";
					when "00010100001001111" => rgb <= "000000";
					when "00010100001010000" => rgb <= "000000";
					when "00010100001010001" => rgb <= "000000";
					when "00010100001010010" => rgb <= "000000";
					when "00010100001010011" => rgb <= "000000";
					when "00010100001010100" => rgb <= "000000";
					when "00010100001010101" => rgb <= "000000";
					when "00010100001010110" => rgb <= "000000";
					when "00010100001010111" => rgb <= "000000";
					when "00010100001011000" => rgb <= "000000";
					when "00010100001011001" => rgb <= "000000";
					when "00010100001011010" => rgb <= "000000";
					when "00010100001011011" => rgb <= "000000";
					when "00010100001011100" => rgb <= "000000";
					when "00010100001011101" => rgb <= "000000";
					when "00010100001011110" => rgb <= "000000";
					when "00010100001011111" => rgb <= "000000";
					when "00010100001100000" => rgb <= "000000";
					when "00010100001100001" => rgb <= "000000";
					when "00010100001100010" => rgb <= "000000";
					when "00010100001100011" => rgb <= "000000";
					when "00010100001100100" => rgb <= "000000";
					when "00010100001100101" => rgb <= "000000";
					when "00010100001100110" => rgb <= "000000";
					when "00010100001100111" => rgb <= "000000";
					when "00010100001101000" => rgb <= "000000";
					when "00010100001101001" => rgb <= "000000";
					when "00010100001101010" => rgb <= "000000";
					when "00010100001101011" => rgb <= "000000";
					when "00010100001101100" => rgb <= "000000";
					when "00010100001101101" => rgb <= "000000";
					when "00010100001101110" => rgb <= "000000";
					when "00010100001101111" => rgb <= "000000";
					when "00010100001110000" => rgb <= "000000";
					when "00010100001110001" => rgb <= "000000";
					when "00010100001110010" => rgb <= "000000";
					when "00010100001110011" => rgb <= "000000";
					when "00010100001110100" => rgb <= "000000";
					when "00010100001110101" => rgb <= "000000";
					when "00010100001110110" => rgb <= "000000";
					when "00010100001110111" => rgb <= "000000";
					when "00010100001111000" => rgb <= "000000";
					when "00010100001111001" => rgb <= "000000";
					when "00010100001111010" => rgb <= "000000";
					when "00010100001111011" => rgb <= "000000";
					when "00010100001111100" => rgb <= "000000";
					when "00010100001111101" => rgb <= "101000";
					when "00010100001111110" => rgb <= "101000";
					when "00010100001111111" => rgb <= "101000";
					when "00010100010000000" => rgb <= "101000";
					when "00010100010000001" => rgb <= "101000";
					when "00010100010000010" => rgb <= "101000";
					when "00010100010000011" => rgb <= "101000";
					when "00010100010000100" => rgb <= "101000";
					when "00010100010000101" => rgb <= "101000";
					when "00010100010000110" => rgb <= "101000";
					when "00010100010000111" => rgb <= "101000";
					when "00010100010001000" => rgb <= "101000";
					when "00010100010001001" => rgb <= "101000";
					when "00010100010001010" => rgb <= "101000";
					when "00010100010001011" => rgb <= "101000";
					when "00010100010001100" => rgb <= "101000";
					when "00010100010001101" => rgb <= "101000";
					when "00010100010001110" => rgb <= "101000";
					when "00010100010001111" => rgb <= "101000";
					when "00010100010010000" => rgb <= "101000";
					when "00010100010010001" => rgb <= "101000";
					when "00010100010010010" => rgb <= "101000";
					when "00010100010010011" => rgb <= "101000";
					when "00010100010010100" => rgb <= "101000";
					when "00010100010010101" => rgb <= "101000";
					when "00010100010010110" => rgb <= "101000";
					when "00010100010010111" => rgb <= "101000";
					when "00010100010011000" => rgb <= "101000";
					when "00010100010011001" => rgb <= "101000";
					when "00010100010011010" => rgb <= "101000";
					when "00010100010011011" => rgb <= "101000";
					when "00010100010011100" => rgb <= "101000";
					when "00010100010011101" => rgb <= "101000";
					when "00010100010011110" => rgb <= "101000";
					when "00010100010011111" => rgb <= "101000";
					when "00010100010100000" => rgb <= "101000";
					when "00010100010100001" => rgb <= "101000";
					when "00010100010100010" => rgb <= "101000";
					when "00010100010100011" => rgb <= "101000";
					when "00010100010100100" => rgb <= "101000";
					when "00010100010100101" => rgb <= "101000";
					when "00010100010100110" => rgb <= "101000";
					when "00010100010100111" => rgb <= "101000";
					when "00010100010101000" => rgb <= "101000";
					when "00010100010101001" => rgb <= "101000";
					when "00010100010101010" => rgb <= "101000";
					when "00010100010101011" => rgb <= "101000";
					when "00010100010101100" => rgb <= "101000";
					when "00010100010101101" => rgb <= "101000";
					when "00010100010101110" => rgb <= "101000";
					when "00010100010101111" => rgb <= "101000";
					when "00010100010110000" => rgb <= "101000";
					when "00010100010110001" => rgb <= "101000";
					when "00010100010110010" => rgb <= "101000";
					when "00010100010110011" => rgb <= "101000";
					when "00010100010110100" => rgb <= "101000";
					when "00010100010110101" => rgb <= "101000";
					when "00010100010110110" => rgb <= "101000";
					when "00010100010110111" => rgb <= "101000";
					when "00010100010111000" => rgb <= "101000";
					when "00010100010111001" => rgb <= "101000";
					when "00010100010111010" => rgb <= "101000";
					when "00010100010111011" => rgb <= "101000";
					when "00010100010111100" => rgb <= "101000";
					when "00010100010111101" => rgb <= "101000";
					when "00010100010111110" => rgb <= "101000";
					when "00010100010111111" => rgb <= "101000";
					when "00010100011000000" => rgb <= "100100";
					when "00010100011000001" => rgb <= "000000";
					when "00010100011000010" => rgb <= "000000";
					when "00010100011000011" => rgb <= "000000";
					when "00010100011000100" => rgb <= "000000";
					when "00010100011000101" => rgb <= "000000";
					when "00010100011000110" => rgb <= "000000";
					when "00010100011000111" => rgb <= "000000";
					when "00010100011001000" => rgb <= "000000";
					when "00010100011001001" => rgb <= "000000";
					when "00010100011001010" => rgb <= "000000";
					when "00010100011001011" => rgb <= "000000";
					when "00010100011001100" => rgb <= "000000";
					when "00010100011001101" => rgb <= "000000";
					when "00010100011001110" => rgb <= "000000";
					when "00010100011001111" => rgb <= "000000";
					when "00010100011010000" => rgb <= "000000";
					when "00010100011010001" => rgb <= "000000";
					when "00010100011010010" => rgb <= "000000";
					when "00010100011010011" => rgb <= "000000";
					when "00010100011010100" => rgb <= "000000";
					when "00010100011010101" => rgb <= "000000";
					when "00010100011010110" => rgb <= "000000";
					when "00010100011010111" => rgb <= "000000";
					when "00010100011011000" => rgb <= "000000";
					when "00010100011011001" => rgb <= "000000";
					when "00010100011011010" => rgb <= "000000";
					when "00010100011011011" => rgb <= "000000";
					when "00010100011011100" => rgb <= "000000";
					when "00010100011011101" => rgb <= "000000";
					when "00010100011011110" => rgb <= "000000";
					when "00010100011011111" => rgb <= "000000";
					when "00010100011100000" => rgb <= "000000";
					when "00010100011100001" => rgb <= "000000";
					when "00010100011100010" => rgb <= "000000";
					when "00010100011100011" => rgb <= "000000";
					when "00010100011100100" => rgb <= "000000";
					when "00010100011100101" => rgb <= "000000";
					when "00010100011100110" => rgb <= "000000";
					when "00010100011100111" => rgb <= "000000";
					when "00010100011101000" => rgb <= "000000";
					when "00010100011101001" => rgb <= "000000";
					when "00010100011101010" => rgb <= "000000";
					when "00010100011101011" => rgb <= "000000";
					when "00010100011101100" => rgb <= "000000";
					when "00010100011101101" => rgb <= "000000";
					when "00010100011101110" => rgb <= "000000";
					when "00010100011101111" => rgb <= "000000";
					when "00010100011110000" => rgb <= "000000";
					when "00010100011110001" => rgb <= "000000";
					when "00010100011110010" => rgb <= "000000";
					when "00010100011110011" => rgb <= "000000";
					when "00010100011110100" => rgb <= "000000";
					when "00010100011110101" => rgb <= "000000";
					when "00010100011110110" => rgb <= "000000";
					when "00010100011110111" => rgb <= "000000";
					when "00010100011111000" => rgb <= "000000";
					when "00010100011111001" => rgb <= "000000";
					when "00010100011111010" => rgb <= "000000";
					when "00010100011111011" => rgb <= "000000";
					when "00010100011111100" => rgb <= "000000";
					when "00010100011111101" => rgb <= "000000";
					when "00010100011111110" => rgb <= "000000";
					when "00010100011111111" => rgb <= "000000";
					when "00010100100000000" => rgb <= "000000";
					when "00010100100000001" => rgb <= "000000";
					when "00010100100000010" => rgb <= "000000";
					when "00010100100000011" => rgb <= "000000";
					when "00010100100000100" => rgb <= "000000";
					when "00010100100000101" => rgb <= "000000";
					when "00010100100000110" => rgb <= "000000";
					when "00010100100000111" => rgb <= "000000";
					when "00010100100001000" => rgb <= "000000";
					when "00010100100001001" => rgb <= "000000";
					when "00010100100001010" => rgb <= "000000";
					when "00010100100001011" => rgb <= "000000";
					when "00010100100001100" => rgb <= "000000";
					when "00010100100001101" => rgb <= "000000";
					when "00010100100001110" => rgb <= "000000";
					when "00010100100001111" => rgb <= "000000";
					when "00010100100010000" => rgb <= "000000";
					when "00010100100010001" => rgb <= "000000";
					when "00010100100010010" => rgb <= "000000";
					when "00010100100010011" => rgb <= "000000";
					when "00010100100010100" => rgb <= "000000";
					when "00010100100010101" => rgb <= "000000";
					when "00010100100010110" => rgb <= "000000";
					when "00010100100010111" => rgb <= "000000";
					when "00010100100011000" => rgb <= "000000";
					when "00010100100011001" => rgb <= "000000";
					when "00010100100011010" => rgb <= "000000";
					when "00010100100011011" => rgb <= "000000";
					when "00010100100011100" => rgb <= "000000";
					when "00010100100011101" => rgb <= "000000";
					when "00010100100011110" => rgb <= "000000";
					when "00010100100011111" => rgb <= "000000";
					when "00010100100100000" => rgb <= "000000";
					when "00010100100100001" => rgb <= "000000";
					when "00010100100100010" => rgb <= "000000";
					when "00010100100100011" => rgb <= "000000";
					when "00010100100100100" => rgb <= "000000";
					when "00010100100100101" => rgb <= "000000";
					when "00010100100100110" => rgb <= "000000";
					when "00010100100100111" => rgb <= "000000";
					when "00010100100101000" => rgb <= "000000";
					when "00010100100101001" => rgb <= "000000";
					when "00010100100101010" => rgb <= "000000";
					when "00010100100101011" => rgb <= "000000";
					when "00010100100101100" => rgb <= "000000";
					when "00010100100101101" => rgb <= "000000";
					when "00010100100101110" => rgb <= "000000";
					when "00010100100101111" => rgb <= "000000";
					when "00010100100110000" => rgb <= "000000";
					when "00010100100110001" => rgb <= "000000";
					when "00010100100110010" => rgb <= "000000";
					when "00010100100110011" => rgb <= "000000";
					when "00010100100110100" => rgb <= "000000";
					when "00010100100110101" => rgb <= "000000";
					when "00010100100110110" => rgb <= "000000";
					when "00010100100110111" => rgb <= "000000";
					when "00010100100111000" => rgb <= "000000";
					when "00010100100111001" => rgb <= "000000";
					when "00010100100111010" => rgb <= "000000";
					when "00010100100111011" => rgb <= "000000";
					when "00010100100111100" => rgb <= "000000";
					when "00010100100111101" => rgb <= "000000";
					when "00010100100111110" => rgb <= "000000";
					when "00010100100111111" => rgb <= "000000";
					when "00010101000000000" => rgb <= "000000";
					when "00010101000000001" => rgb <= "000000";
					when "00010101000000010" => rgb <= "000000";
					when "00010101000000011" => rgb <= "000000";
					when "00010101000000100" => rgb <= "000000";
					when "00010101000000101" => rgb <= "000000";
					when "00010101000000110" => rgb <= "000000";
					when "00010101000000111" => rgb <= "000000";
					when "00010101000001000" => rgb <= "000000";
					when "00010101000001001" => rgb <= "000000";
					when "00010101000001010" => rgb <= "000000";
					when "00010101000001011" => rgb <= "000000";
					when "00010101000001100" => rgb <= "000000";
					when "00010101000001101" => rgb <= "000000";
					when "00010101000001110" => rgb <= "000000";
					when "00010101000001111" => rgb <= "000000";
					when "00010101000010000" => rgb <= "000000";
					when "00010101000010001" => rgb <= "000000";
					when "00010101000010010" => rgb <= "000000";
					when "00010101000010011" => rgb <= "000000";
					when "00010101000010100" => rgb <= "000000";
					when "00010101000010101" => rgb <= "000000";
					when "00010101000010110" => rgb <= "000000";
					when "00010101000010111" => rgb <= "000000";
					when "00010101000011000" => rgb <= "000000";
					when "00010101000011001" => rgb <= "000000";
					when "00010101000011010" => rgb <= "000000";
					when "00010101000011011" => rgb <= "000000";
					when "00010101000011100" => rgb <= "000000";
					when "00010101000011101" => rgb <= "000000";
					when "00010101000011110" => rgb <= "000000";
					when "00010101000011111" => rgb <= "000000";
					when "00010101000100000" => rgb <= "000000";
					when "00010101000100001" => rgb <= "000000";
					when "00010101000100010" => rgb <= "000000";
					when "00010101000100011" => rgb <= "000000";
					when "00010101000100100" => rgb <= "000000";
					when "00010101000100101" => rgb <= "000000";
					when "00010101000100110" => rgb <= "000000";
					when "00010101000100111" => rgb <= "000000";
					when "00010101000101000" => rgb <= "000000";
					when "00010101000101001" => rgb <= "000000";
					when "00010101000101010" => rgb <= "000000";
					when "00010101000101011" => rgb <= "000000";
					when "00010101000101100" => rgb <= "000000";
					when "00010101000101101" => rgb <= "000000";
					when "00010101000101110" => rgb <= "000000";
					when "00010101000101111" => rgb <= "000000";
					when "00010101000110000" => rgb <= "000000";
					when "00010101000110001" => rgb <= "000000";
					when "00010101000110010" => rgb <= "000000";
					when "00010101000110011" => rgb <= "000000";
					when "00010101000110100" => rgb <= "000000";
					when "00010101000110101" => rgb <= "000000";
					when "00010101000110110" => rgb <= "000000";
					when "00010101000110111" => rgb <= "000000";
					when "00010101000111000" => rgb <= "000000";
					when "00010101000111001" => rgb <= "000000";
					when "00010101000111010" => rgb <= "000000";
					when "00010101000111011" => rgb <= "000000";
					when "00010101000111100" => rgb <= "000000";
					when "00010101000111101" => rgb <= "000000";
					when "00010101000111110" => rgb <= "000000";
					when "00010101000111111" => rgb <= "000000";
					when "00010101001000000" => rgb <= "000000";
					when "00010101001000001" => rgb <= "000000";
					when "00010101001000010" => rgb <= "000000";
					when "00010101001000011" => rgb <= "000000";
					when "00010101001000100" => rgb <= "000000";
					when "00010101001000101" => rgb <= "000000";
					when "00010101001000110" => rgb <= "000000";
					when "00010101001000111" => rgb <= "000000";
					when "00010101001001000" => rgb <= "000000";
					when "00010101001001001" => rgb <= "000000";
					when "00010101001001010" => rgb <= "000000";
					when "00010101001001011" => rgb <= "000000";
					when "00010101001001100" => rgb <= "000000";
					when "00010101001001101" => rgb <= "000000";
					when "00010101001001110" => rgb <= "000000";
					when "00010101001001111" => rgb <= "000000";
					when "00010101001010000" => rgb <= "000000";
					when "00010101001010001" => rgb <= "000000";
					when "00010101001010010" => rgb <= "000000";
					when "00010101001010011" => rgb <= "000000";
					when "00010101001010100" => rgb <= "000000";
					when "00010101001010101" => rgb <= "000000";
					when "00010101001010110" => rgb <= "000000";
					when "00010101001010111" => rgb <= "000000";
					when "00010101001011000" => rgb <= "000000";
					when "00010101001011001" => rgb <= "000000";
					when "00010101001011010" => rgb <= "000000";
					when "00010101001011011" => rgb <= "000000";
					when "00010101001011100" => rgb <= "000000";
					when "00010101001011101" => rgb <= "000000";
					when "00010101001011110" => rgb <= "000000";
					when "00010101001011111" => rgb <= "000000";
					when "00010101001100000" => rgb <= "000000";
					when "00010101001100001" => rgb <= "000000";
					when "00010101001100010" => rgb <= "000000";
					when "00010101001100011" => rgb <= "000000";
					when "00010101001100100" => rgb <= "000000";
					when "00010101001100101" => rgb <= "000000";
					when "00010101001100110" => rgb <= "000000";
					when "00010101001100111" => rgb <= "000000";
					when "00010101001101000" => rgb <= "000000";
					when "00010101001101001" => rgb <= "000000";
					when "00010101001101010" => rgb <= "000000";
					when "00010101001101011" => rgb <= "000000";
					when "00010101001101100" => rgb <= "000000";
					when "00010101001101101" => rgb <= "000000";
					when "00010101001101110" => rgb <= "000000";
					when "00010101001101111" => rgb <= "000000";
					when "00010101001110000" => rgb <= "000000";
					when "00010101001110001" => rgb <= "000000";
					when "00010101001110010" => rgb <= "000000";
					when "00010101001110011" => rgb <= "000000";
					when "00010101001110100" => rgb <= "000000";
					when "00010101001110101" => rgb <= "000000";
					when "00010101001110110" => rgb <= "000000";
					when "00010101001110111" => rgb <= "000000";
					when "00010101001111000" => rgb <= "000000";
					when "00010101001111001" => rgb <= "000000";
					when "00010101001111010" => rgb <= "000000";
					when "00010101001111011" => rgb <= "000000";
					when "00010101001111100" => rgb <= "000000";
					when "00010101001111101" => rgb <= "101000";
					when "00010101001111110" => rgb <= "101000";
					when "00010101001111111" => rgb <= "101000";
					when "00010101010000000" => rgb <= "101000";
					when "00010101010000001" => rgb <= "101000";
					when "00010101010000010" => rgb <= "101000";
					when "00010101010000011" => rgb <= "101000";
					when "00010101010000100" => rgb <= "101000";
					when "00010101010000101" => rgb <= "101000";
					when "00010101010000110" => rgb <= "101000";
					when "00010101010000111" => rgb <= "101000";
					when "00010101010001000" => rgb <= "101000";
					when "00010101010001001" => rgb <= "101000";
					when "00010101010001010" => rgb <= "101000";
					when "00010101010001011" => rgb <= "101000";
					when "00010101010001100" => rgb <= "101000";
					when "00010101010001101" => rgb <= "101000";
					when "00010101010001110" => rgb <= "101000";
					when "00010101010001111" => rgb <= "101000";
					when "00010101010010000" => rgb <= "101000";
					when "00010101010010001" => rgb <= "101000";
					when "00010101010010010" => rgb <= "101000";
					when "00010101010010011" => rgb <= "101000";
					when "00010101010010100" => rgb <= "101000";
					when "00010101010010101" => rgb <= "101000";
					when "00010101010010110" => rgb <= "101000";
					when "00010101010010111" => rgb <= "101000";
					when "00010101010011000" => rgb <= "101000";
					when "00010101010011001" => rgb <= "101000";
					when "00010101010011010" => rgb <= "101000";
					when "00010101010011011" => rgb <= "101000";
					when "00010101010011100" => rgb <= "101000";
					when "00010101010011101" => rgb <= "101000";
					when "00010101010011110" => rgb <= "101000";
					when "00010101010011111" => rgb <= "101000";
					when "00010101010100000" => rgb <= "101000";
					when "00010101010100001" => rgb <= "101000";
					when "00010101010100010" => rgb <= "101000";
					when "00010101010100011" => rgb <= "101000";
					when "00010101010100100" => rgb <= "101000";
					when "00010101010100101" => rgb <= "101000";
					when "00010101010100110" => rgb <= "101000";
					when "00010101010100111" => rgb <= "101000";
					when "00010101010101000" => rgb <= "101000";
					when "00010101010101001" => rgb <= "101000";
					when "00010101010101010" => rgb <= "101000";
					when "00010101010101011" => rgb <= "101000";
					when "00010101010101100" => rgb <= "101000";
					when "00010101010101101" => rgb <= "101000";
					when "00010101010101110" => rgb <= "101000";
					when "00010101010101111" => rgb <= "101000";
					when "00010101010110000" => rgb <= "101000";
					when "00010101010110001" => rgb <= "101000";
					when "00010101010110010" => rgb <= "101000";
					when "00010101010110011" => rgb <= "101000";
					when "00010101010110100" => rgb <= "101000";
					when "00010101010110101" => rgb <= "101000";
					when "00010101010110110" => rgb <= "101000";
					when "00010101010110111" => rgb <= "101000";
					when "00010101010111000" => rgb <= "101000";
					when "00010101010111001" => rgb <= "101000";
					when "00010101010111010" => rgb <= "101000";
					when "00010101010111011" => rgb <= "101000";
					when "00010101010111100" => rgb <= "101000";
					when "00010101010111101" => rgb <= "101000";
					when "00010101010111110" => rgb <= "101000";
					when "00010101010111111" => rgb <= "101000";
					when "00010101011000000" => rgb <= "100100";
					when "00010101011000001" => rgb <= "000000";
					when "00010101011000010" => rgb <= "000000";
					when "00010101011000011" => rgb <= "000000";
					when "00010101011000100" => rgb <= "000000";
					when "00010101011000101" => rgb <= "000000";
					when "00010101011000110" => rgb <= "000000";
					when "00010101011000111" => rgb <= "000000";
					when "00010101011001000" => rgb <= "000000";
					when "00010101011001001" => rgb <= "000000";
					when "00010101011001010" => rgb <= "000000";
					when "00010101011001011" => rgb <= "000000";
					when "00010101011001100" => rgb <= "000000";
					when "00010101011001101" => rgb <= "000000";
					when "00010101011001110" => rgb <= "000000";
					when "00010101011001111" => rgb <= "000000";
					when "00010101011010000" => rgb <= "000000";
					when "00010101011010001" => rgb <= "000000";
					when "00010101011010010" => rgb <= "000000";
					when "00010101011010011" => rgb <= "000000";
					when "00010101011010100" => rgb <= "000000";
					when "00010101011010101" => rgb <= "000000";
					when "00010101011010110" => rgb <= "000000";
					when "00010101011010111" => rgb <= "000000";
					when "00010101011011000" => rgb <= "000000";
					when "00010101011011001" => rgb <= "000000";
					when "00010101011011010" => rgb <= "000000";
					when "00010101011011011" => rgb <= "000000";
					when "00010101011011100" => rgb <= "000000";
					when "00010101011011101" => rgb <= "000000";
					when "00010101011011110" => rgb <= "000000";
					when "00010101011011111" => rgb <= "000000";
					when "00010101011100000" => rgb <= "000000";
					when "00010101011100001" => rgb <= "000000";
					when "00010101011100010" => rgb <= "000000";
					when "00010101011100011" => rgb <= "000000";
					when "00010101011100100" => rgb <= "000000";
					when "00010101011100101" => rgb <= "000000";
					when "00010101011100110" => rgb <= "000000";
					when "00010101011100111" => rgb <= "000000";
					when "00010101011101000" => rgb <= "000000";
					when "00010101011101001" => rgb <= "000000";
					when "00010101011101010" => rgb <= "000000";
					when "00010101011101011" => rgb <= "000000";
					when "00010101011101100" => rgb <= "000000";
					when "00010101011101101" => rgb <= "000000";
					when "00010101011101110" => rgb <= "000000";
					when "00010101011101111" => rgb <= "000000";
					when "00010101011110000" => rgb <= "000000";
					when "00010101011110001" => rgb <= "000000";
					when "00010101011110010" => rgb <= "000000";
					when "00010101011110011" => rgb <= "000000";
					when "00010101011110100" => rgb <= "000000";
					when "00010101011110101" => rgb <= "000000";
					when "00010101011110110" => rgb <= "000000";
					when "00010101011110111" => rgb <= "000000";
					when "00010101011111000" => rgb <= "000000";
					when "00010101011111001" => rgb <= "000000";
					when "00010101011111010" => rgb <= "000000";
					when "00010101011111011" => rgb <= "000000";
					when "00010101011111100" => rgb <= "000000";
					when "00010101011111101" => rgb <= "000000";
					when "00010101011111110" => rgb <= "000000";
					when "00010101011111111" => rgb <= "000000";
					when "00010101100000000" => rgb <= "000000";
					when "00010101100000001" => rgb <= "000000";
					when "00010101100000010" => rgb <= "000000";
					when "00010101100000011" => rgb <= "000000";
					when "00010101100000100" => rgb <= "000000";
					when "00010101100000101" => rgb <= "000000";
					when "00010101100000110" => rgb <= "000000";
					when "00010101100000111" => rgb <= "000000";
					when "00010101100001000" => rgb <= "000000";
					when "00010101100001001" => rgb <= "000000";
					when "00010101100001010" => rgb <= "000000";
					when "00010101100001011" => rgb <= "000000";
					when "00010101100001100" => rgb <= "000000";
					when "00010101100001101" => rgb <= "000000";
					when "00010101100001110" => rgb <= "000000";
					when "00010101100001111" => rgb <= "000000";
					when "00010101100010000" => rgb <= "000000";
					when "00010101100010001" => rgb <= "000000";
					when "00010101100010010" => rgb <= "000000";
					when "00010101100010011" => rgb <= "000000";
					when "00010101100010100" => rgb <= "000000";
					when "00010101100010101" => rgb <= "000000";
					when "00010101100010110" => rgb <= "000000";
					when "00010101100010111" => rgb <= "000000";
					when "00010101100011000" => rgb <= "000000";
					when "00010101100011001" => rgb <= "000000";
					when "00010101100011010" => rgb <= "000000";
					when "00010101100011011" => rgb <= "000000";
					when "00010101100011100" => rgb <= "000000";
					when "00010101100011101" => rgb <= "000000";
					when "00010101100011110" => rgb <= "000000";
					when "00010101100011111" => rgb <= "000000";
					when "00010101100100000" => rgb <= "000000";
					when "00010101100100001" => rgb <= "000000";
					when "00010101100100010" => rgb <= "000000";
					when "00010101100100011" => rgb <= "000000";
					when "00010101100100100" => rgb <= "000000";
					when "00010101100100101" => rgb <= "000000";
					when "00010101100100110" => rgb <= "000000";
					when "00010101100100111" => rgb <= "000000";
					when "00010101100101000" => rgb <= "000000";
					when "00010101100101001" => rgb <= "000000";
					when "00010101100101010" => rgb <= "000000";
					when "00010101100101011" => rgb <= "000000";
					when "00010101100101100" => rgb <= "000000";
					when "00010101100101101" => rgb <= "000000";
					when "00010101100101110" => rgb <= "000000";
					when "00010101100101111" => rgb <= "000000";
					when "00010101100110000" => rgb <= "000000";
					when "00010101100110001" => rgb <= "000000";
					when "00010101100110010" => rgb <= "000000";
					when "00010101100110011" => rgb <= "000000";
					when "00010101100110100" => rgb <= "000000";
					when "00010101100110101" => rgb <= "000000";
					when "00010101100110110" => rgb <= "000000";
					when "00010101100110111" => rgb <= "000000";
					when "00010101100111000" => rgb <= "000000";
					when "00010101100111001" => rgb <= "000000";
					when "00010101100111010" => rgb <= "000000";
					when "00010101100111011" => rgb <= "000000";
					when "00010101100111100" => rgb <= "000000";
					when "00010101100111101" => rgb <= "000000";
					when "00010101100111110" => rgb <= "000000";
					when "00010101100111111" => rgb <= "000000";
					when "00010110000000000" => rgb <= "000000";
					when "00010110000000001" => rgb <= "000000";
					when "00010110000000010" => rgb <= "000000";
					when "00010110000000011" => rgb <= "000000";
					when "00010110000000100" => rgb <= "000000";
					when "00010110000000101" => rgb <= "000000";
					when "00010110000000110" => rgb <= "000000";
					when "00010110000000111" => rgb <= "000000";
					when "00010110000001000" => rgb <= "000000";
					when "00010110000001001" => rgb <= "000000";
					when "00010110000001010" => rgb <= "000000";
					when "00010110000001011" => rgb <= "000000";
					when "00010110000001100" => rgb <= "000000";
					when "00010110000001101" => rgb <= "000000";
					when "00010110000001110" => rgb <= "000000";
					when "00010110000001111" => rgb <= "000000";
					when "00010110000010000" => rgb <= "000000";
					when "00010110000010001" => rgb <= "000000";
					when "00010110000010010" => rgb <= "000000";
					when "00010110000010011" => rgb <= "000000";
					when "00010110000010100" => rgb <= "000000";
					when "00010110000010101" => rgb <= "000000";
					when "00010110000010110" => rgb <= "000000";
					when "00010110000010111" => rgb <= "000000";
					when "00010110000011000" => rgb <= "000000";
					when "00010110000011001" => rgb <= "000000";
					when "00010110000011010" => rgb <= "000000";
					when "00010110000011011" => rgb <= "000000";
					when "00010110000011100" => rgb <= "000000";
					when "00010110000011101" => rgb <= "000000";
					when "00010110000011110" => rgb <= "000000";
					when "00010110000011111" => rgb <= "000000";
					when "00010110000100000" => rgb <= "000000";
					when "00010110000100001" => rgb <= "000000";
					when "00010110000100010" => rgb <= "000000";
					when "00010110000100011" => rgb <= "000000";
					when "00010110000100100" => rgb <= "000000";
					when "00010110000100101" => rgb <= "000000";
					when "00010110000100110" => rgb <= "000000";
					when "00010110000100111" => rgb <= "000000";
					when "00010110000101000" => rgb <= "000000";
					when "00010110000101001" => rgb <= "000000";
					when "00010110000101010" => rgb <= "000000";
					when "00010110000101011" => rgb <= "000000";
					when "00010110000101100" => rgb <= "000000";
					when "00010110000101101" => rgb <= "000000";
					when "00010110000101110" => rgb <= "000000";
					when "00010110000101111" => rgb <= "000000";
					when "00010110000110000" => rgb <= "000000";
					when "00010110000110001" => rgb <= "000000";
					when "00010110000110010" => rgb <= "000000";
					when "00010110000110011" => rgb <= "000000";
					when "00010110000110100" => rgb <= "000000";
					when "00010110000110101" => rgb <= "000000";
					when "00010110000110110" => rgb <= "000000";
					when "00010110000110111" => rgb <= "000000";
					when "00010110000111000" => rgb <= "000000";
					when "00010110000111001" => rgb <= "000000";
					when "00010110000111010" => rgb <= "000000";
					when "00010110000111011" => rgb <= "000000";
					when "00010110000111100" => rgb <= "000000";
					when "00010110000111101" => rgb <= "000000";
					when "00010110000111110" => rgb <= "000000";
					when "00010110000111111" => rgb <= "000000";
					when "00010110001000000" => rgb <= "000000";
					when "00010110001000001" => rgb <= "000000";
					when "00010110001000010" => rgb <= "000000";
					when "00010110001000011" => rgb <= "000000";
					when "00010110001000100" => rgb <= "000000";
					when "00010110001000101" => rgb <= "000000";
					when "00010110001000110" => rgb <= "000000";
					when "00010110001000111" => rgb <= "000000";
					when "00010110001001000" => rgb <= "000000";
					when "00010110001001001" => rgb <= "000000";
					when "00010110001001010" => rgb <= "000000";
					when "00010110001001011" => rgb <= "000000";
					when "00010110001001100" => rgb <= "000000";
					when "00010110001001101" => rgb <= "000000";
					when "00010110001001110" => rgb <= "000000";
					when "00010110001001111" => rgb <= "000000";
					when "00010110001010000" => rgb <= "000000";
					when "00010110001010001" => rgb <= "000000";
					when "00010110001010010" => rgb <= "000000";
					when "00010110001010011" => rgb <= "000000";
					when "00010110001010100" => rgb <= "000000";
					when "00010110001010101" => rgb <= "000000";
					when "00010110001010110" => rgb <= "000000";
					when "00010110001010111" => rgb <= "000000";
					when "00010110001011000" => rgb <= "000000";
					when "00010110001011001" => rgb <= "000000";
					when "00010110001011010" => rgb <= "000000";
					when "00010110001011011" => rgb <= "000000";
					when "00010110001011100" => rgb <= "000000";
					when "00010110001011101" => rgb <= "000000";
					when "00010110001011110" => rgb <= "000000";
					when "00010110001011111" => rgb <= "000000";
					when "00010110001100000" => rgb <= "000000";
					when "00010110001100001" => rgb <= "000000";
					when "00010110001100010" => rgb <= "000000";
					when "00010110001100011" => rgb <= "000000";
					when "00010110001100100" => rgb <= "000000";
					when "00010110001100101" => rgb <= "000000";
					when "00010110001100110" => rgb <= "000000";
					when "00010110001100111" => rgb <= "000000";
					when "00010110001101000" => rgb <= "000000";
					when "00010110001101001" => rgb <= "000000";
					when "00010110001101010" => rgb <= "000000";
					when "00010110001101011" => rgb <= "000000";
					when "00010110001101100" => rgb <= "000000";
					when "00010110001101101" => rgb <= "000000";
					when "00010110001101110" => rgb <= "000000";
					when "00010110001101111" => rgb <= "000000";
					when "00010110001110000" => rgb <= "000000";
					when "00010110001110001" => rgb <= "000000";
					when "00010110001110010" => rgb <= "000000";
					when "00010110001110011" => rgb <= "000000";
					when "00010110001110100" => rgb <= "000000";
					when "00010110001110101" => rgb <= "000000";
					when "00010110001110110" => rgb <= "000000";
					when "00010110001110111" => rgb <= "000000";
					when "00010110001111000" => rgb <= "000000";
					when "00010110001111001" => rgb <= "000000";
					when "00010110001111010" => rgb <= "000000";
					when "00010110001111011" => rgb <= "000000";
					when "00010110001111100" => rgb <= "000000";
					when "00010110001111101" => rgb <= "101000";
					when "00010110001111110" => rgb <= "101000";
					when "00010110001111111" => rgb <= "101000";
					when "00010110010000000" => rgb <= "101000";
					when "00010110010000001" => rgb <= "101000";
					when "00010110010000010" => rgb <= "101000";
					when "00010110010000011" => rgb <= "101000";
					when "00010110010000100" => rgb <= "101000";
					when "00010110010000101" => rgb <= "101000";
					when "00010110010000110" => rgb <= "101000";
					when "00010110010000111" => rgb <= "101000";
					when "00010110010001000" => rgb <= "101000";
					when "00010110010001001" => rgb <= "101000";
					when "00010110010001010" => rgb <= "101000";
					when "00010110010001011" => rgb <= "101000";
					when "00010110010001100" => rgb <= "101000";
					when "00010110010001101" => rgb <= "101000";
					when "00010110010001110" => rgb <= "101000";
					when "00010110010001111" => rgb <= "101000";
					when "00010110010010000" => rgb <= "101000";
					when "00010110010010001" => rgb <= "101000";
					when "00010110010010010" => rgb <= "101000";
					when "00010110010010011" => rgb <= "101000";
					when "00010110010010100" => rgb <= "101000";
					when "00010110010010101" => rgb <= "101000";
					when "00010110010010110" => rgb <= "101000";
					when "00010110010010111" => rgb <= "101000";
					when "00010110010011000" => rgb <= "101000";
					when "00010110010011001" => rgb <= "101000";
					when "00010110010011010" => rgb <= "101000";
					when "00010110010011011" => rgb <= "101000";
					when "00010110010011100" => rgb <= "101000";
					when "00010110010011101" => rgb <= "101000";
					when "00010110010011110" => rgb <= "101000";
					when "00010110010011111" => rgb <= "101000";
					when "00010110010100000" => rgb <= "101000";
					when "00010110010100001" => rgb <= "101000";
					when "00010110010100010" => rgb <= "101000";
					when "00010110010100011" => rgb <= "101000";
					when "00010110010100100" => rgb <= "101000";
					when "00010110010100101" => rgb <= "101000";
					when "00010110010100110" => rgb <= "101000";
					when "00010110010100111" => rgb <= "101000";
					when "00010110010101000" => rgb <= "101000";
					when "00010110010101001" => rgb <= "101000";
					when "00010110010101010" => rgb <= "101000";
					when "00010110010101011" => rgb <= "101000";
					when "00010110010101100" => rgb <= "101000";
					when "00010110010101101" => rgb <= "101000";
					when "00010110010101110" => rgb <= "101000";
					when "00010110010101111" => rgb <= "101000";
					when "00010110010110000" => rgb <= "101000";
					when "00010110010110001" => rgb <= "101000";
					when "00010110010110010" => rgb <= "101000";
					when "00010110010110011" => rgb <= "101000";
					when "00010110010110100" => rgb <= "101000";
					when "00010110010110101" => rgb <= "101000";
					when "00010110010110110" => rgb <= "101000";
					when "00010110010110111" => rgb <= "101000";
					when "00010110010111000" => rgb <= "101000";
					when "00010110010111001" => rgb <= "101000";
					when "00010110010111010" => rgb <= "101000";
					when "00010110010111011" => rgb <= "101000";
					when "00010110010111100" => rgb <= "101000";
					when "00010110010111101" => rgb <= "101000";
					when "00010110010111110" => rgb <= "101000";
					when "00010110010111111" => rgb <= "101000";
					when "00010110011000000" => rgb <= "100100";
					when "00010110011000001" => rgb <= "000000";
					when "00010110011000010" => rgb <= "000000";
					when "00010110011000011" => rgb <= "000000";
					when "00010110011000100" => rgb <= "000000";
					when "00010110011000101" => rgb <= "000000";
					when "00010110011000110" => rgb <= "000000";
					when "00010110011000111" => rgb <= "000000";
					when "00010110011001000" => rgb <= "000000";
					when "00010110011001001" => rgb <= "000000";
					when "00010110011001010" => rgb <= "000000";
					when "00010110011001011" => rgb <= "000000";
					when "00010110011001100" => rgb <= "000000";
					when "00010110011001101" => rgb <= "000000";
					when "00010110011001110" => rgb <= "000000";
					when "00010110011001111" => rgb <= "000000";
					when "00010110011010000" => rgb <= "000000";
					when "00010110011010001" => rgb <= "000000";
					when "00010110011010010" => rgb <= "000000";
					when "00010110011010011" => rgb <= "000000";
					when "00010110011010100" => rgb <= "000000";
					when "00010110011010101" => rgb <= "000000";
					when "00010110011010110" => rgb <= "000000";
					when "00010110011010111" => rgb <= "000000";
					when "00010110011011000" => rgb <= "000000";
					when "00010110011011001" => rgb <= "000000";
					when "00010110011011010" => rgb <= "000000";
					when "00010110011011011" => rgb <= "000000";
					when "00010110011011100" => rgb <= "000000";
					when "00010110011011101" => rgb <= "000000";
					when "00010110011011110" => rgb <= "000000";
					when "00010110011011111" => rgb <= "000000";
					when "00010110011100000" => rgb <= "000000";
					when "00010110011100001" => rgb <= "000000";
					when "00010110011100010" => rgb <= "000000";
					when "00010110011100011" => rgb <= "000000";
					when "00010110011100100" => rgb <= "000000";
					when "00010110011100101" => rgb <= "000000";
					when "00010110011100110" => rgb <= "000000";
					when "00010110011100111" => rgb <= "000000";
					when "00010110011101000" => rgb <= "000000";
					when "00010110011101001" => rgb <= "000000";
					when "00010110011101010" => rgb <= "000000";
					when "00010110011101011" => rgb <= "000000";
					when "00010110011101100" => rgb <= "000000";
					when "00010110011101101" => rgb <= "000000";
					when "00010110011101110" => rgb <= "000000";
					when "00010110011101111" => rgb <= "000000";
					when "00010110011110000" => rgb <= "000000";
					when "00010110011110001" => rgb <= "000000";
					when "00010110011110010" => rgb <= "000000";
					when "00010110011110011" => rgb <= "000000";
					when "00010110011110100" => rgb <= "000000";
					when "00010110011110101" => rgb <= "000000";
					when "00010110011110110" => rgb <= "000000";
					when "00010110011110111" => rgb <= "000000";
					when "00010110011111000" => rgb <= "000000";
					when "00010110011111001" => rgb <= "000000";
					when "00010110011111010" => rgb <= "000000";
					when "00010110011111011" => rgb <= "000000";
					when "00010110011111100" => rgb <= "000000";
					when "00010110011111101" => rgb <= "000000";
					when "00010110011111110" => rgb <= "000000";
					when "00010110011111111" => rgb <= "000000";
					when "00010110100000000" => rgb <= "000000";
					when "00010110100000001" => rgb <= "000000";
					when "00010110100000010" => rgb <= "000000";
					when "00010110100000011" => rgb <= "000000";
					when "00010110100000100" => rgb <= "000000";
					when "00010110100000101" => rgb <= "000000";
					when "00010110100000110" => rgb <= "000000";
					when "00010110100000111" => rgb <= "000000";
					when "00010110100001000" => rgb <= "000000";
					when "00010110100001001" => rgb <= "000000";
					when "00010110100001010" => rgb <= "000000";
					when "00010110100001011" => rgb <= "000000";
					when "00010110100001100" => rgb <= "000000";
					when "00010110100001101" => rgb <= "000000";
					when "00010110100001110" => rgb <= "000000";
					when "00010110100001111" => rgb <= "000000";
					when "00010110100010000" => rgb <= "000000";
					when "00010110100010001" => rgb <= "000000";
					when "00010110100010010" => rgb <= "000000";
					when "00010110100010011" => rgb <= "000000";
					when "00010110100010100" => rgb <= "000000";
					when "00010110100010101" => rgb <= "000000";
					when "00010110100010110" => rgb <= "000000";
					when "00010110100010111" => rgb <= "000000";
					when "00010110100011000" => rgb <= "000000";
					when "00010110100011001" => rgb <= "000000";
					when "00010110100011010" => rgb <= "000000";
					when "00010110100011011" => rgb <= "000000";
					when "00010110100011100" => rgb <= "000000";
					when "00010110100011101" => rgb <= "000000";
					when "00010110100011110" => rgb <= "000000";
					when "00010110100011111" => rgb <= "000000";
					when "00010110100100000" => rgb <= "000000";
					when "00010110100100001" => rgb <= "000000";
					when "00010110100100010" => rgb <= "000000";
					when "00010110100100011" => rgb <= "000000";
					when "00010110100100100" => rgb <= "000000";
					when "00010110100100101" => rgb <= "000000";
					when "00010110100100110" => rgb <= "000000";
					when "00010110100100111" => rgb <= "000000";
					when "00010110100101000" => rgb <= "000000";
					when "00010110100101001" => rgb <= "000000";
					when "00010110100101010" => rgb <= "000000";
					when "00010110100101011" => rgb <= "000000";
					when "00010110100101100" => rgb <= "000000";
					when "00010110100101101" => rgb <= "000000";
					when "00010110100101110" => rgb <= "000000";
					when "00010110100101111" => rgb <= "000000";
					when "00010110100110000" => rgb <= "000000";
					when "00010110100110001" => rgb <= "000000";
					when "00010110100110010" => rgb <= "000000";
					when "00010110100110011" => rgb <= "000000";
					when "00010110100110100" => rgb <= "000000";
					when "00010110100110101" => rgb <= "000000";
					when "00010110100110110" => rgb <= "000000";
					when "00010110100110111" => rgb <= "000000";
					when "00010110100111000" => rgb <= "000000";
					when "00010110100111001" => rgb <= "000000";
					when "00010110100111010" => rgb <= "000000";
					when "00010110100111011" => rgb <= "000000";
					when "00010110100111100" => rgb <= "000000";
					when "00010110100111101" => rgb <= "000000";
					when "00010110100111110" => rgb <= "000000";
					when "00010110100111111" => rgb <= "000000";
					when "00010111000000000" => rgb <= "000000";
					when "00010111000000001" => rgb <= "000000";
					when "00010111000000010" => rgb <= "000000";
					when "00010111000000011" => rgb <= "000000";
					when "00010111000000100" => rgb <= "000000";
					when "00010111000000101" => rgb <= "000000";
					when "00010111000000110" => rgb <= "000000";
					when "00010111000000111" => rgb <= "000000";
					when "00010111000001000" => rgb <= "000000";
					when "00010111000001001" => rgb <= "000000";
					when "00010111000001010" => rgb <= "000000";
					when "00010111000001011" => rgb <= "000000";
					when "00010111000001100" => rgb <= "000000";
					when "00010111000001101" => rgb <= "000000";
					when "00010111000001110" => rgb <= "000000";
					when "00010111000001111" => rgb <= "000000";
					when "00010111000010000" => rgb <= "000000";
					when "00010111000010001" => rgb <= "000000";
					when "00010111000010010" => rgb <= "000000";
					when "00010111000010011" => rgb <= "000000";
					when "00010111000010100" => rgb <= "000000";
					when "00010111000010101" => rgb <= "000000";
					when "00010111000010110" => rgb <= "000000";
					when "00010111000010111" => rgb <= "000000";
					when "00010111000011000" => rgb <= "000000";
					when "00010111000011001" => rgb <= "000000";
					when "00010111000011010" => rgb <= "000000";
					when "00010111000011011" => rgb <= "000000";
					when "00010111000011100" => rgb <= "000000";
					when "00010111000011101" => rgb <= "000000";
					when "00010111000011110" => rgb <= "000000";
					when "00010111000011111" => rgb <= "000000";
					when "00010111000100000" => rgb <= "000000";
					when "00010111000100001" => rgb <= "000000";
					when "00010111000100010" => rgb <= "000000";
					when "00010111000100011" => rgb <= "000000";
					when "00010111000100100" => rgb <= "000000";
					when "00010111000100101" => rgb <= "000000";
					when "00010111000100110" => rgb <= "000000";
					when "00010111000100111" => rgb <= "000000";
					when "00010111000101000" => rgb <= "000000";
					when "00010111000101001" => rgb <= "000000";
					when "00010111000101010" => rgb <= "000000";
					when "00010111000101011" => rgb <= "000000";
					when "00010111000101100" => rgb <= "000000";
					when "00010111000101101" => rgb <= "000000";
					when "00010111000101110" => rgb <= "000000";
					when "00010111000101111" => rgb <= "000000";
					when "00010111000110000" => rgb <= "000000";
					when "00010111000110001" => rgb <= "000000";
					when "00010111000110010" => rgb <= "000000";
					when "00010111000110011" => rgb <= "000000";
					when "00010111000110100" => rgb <= "000000";
					when "00010111000110101" => rgb <= "000000";
					when "00010111000110110" => rgb <= "000000";
					when "00010111000110111" => rgb <= "000000";
					when "00010111000111000" => rgb <= "000000";
					when "00010111000111001" => rgb <= "000000";
					when "00010111000111010" => rgb <= "000000";
					when "00010111000111011" => rgb <= "000000";
					when "00010111000111100" => rgb <= "000000";
					when "00010111000111101" => rgb <= "000000";
					when "00010111000111110" => rgb <= "000000";
					when "00010111000111111" => rgb <= "000000";
					when "00010111001000000" => rgb <= "000000";
					when "00010111001000001" => rgb <= "000000";
					when "00010111001000010" => rgb <= "000000";
					when "00010111001000011" => rgb <= "000000";
					when "00010111001000100" => rgb <= "000000";
					when "00010111001000101" => rgb <= "000000";
					when "00010111001000110" => rgb <= "000000";
					when "00010111001000111" => rgb <= "000000";
					when "00010111001001000" => rgb <= "000000";
					when "00010111001001001" => rgb <= "000000";
					when "00010111001001010" => rgb <= "000000";
					when "00010111001001011" => rgb <= "000000";
					when "00010111001001100" => rgb <= "000000";
					when "00010111001001101" => rgb <= "000000";
					when "00010111001001110" => rgb <= "000000";
					when "00010111001001111" => rgb <= "000000";
					when "00010111001010000" => rgb <= "000000";
					when "00010111001010001" => rgb <= "000000";
					when "00010111001010010" => rgb <= "000000";
					when "00010111001010011" => rgb <= "000000";
					when "00010111001010100" => rgb <= "000000";
					when "00010111001010101" => rgb <= "000000";
					when "00010111001010110" => rgb <= "000000";
					when "00010111001010111" => rgb <= "000000";
					when "00010111001011000" => rgb <= "000000";
					when "00010111001011001" => rgb <= "000000";
					when "00010111001011010" => rgb <= "000000";
					when "00010111001011011" => rgb <= "000000";
					when "00010111001011100" => rgb <= "000000";
					when "00010111001011101" => rgb <= "000000";
					when "00010111001011110" => rgb <= "000000";
					when "00010111001011111" => rgb <= "000000";
					when "00010111001100000" => rgb <= "000000";
					when "00010111001100001" => rgb <= "000000";
					when "00010111001100010" => rgb <= "000000";
					when "00010111001100011" => rgb <= "000000";
					when "00010111001100100" => rgb <= "000000";
					when "00010111001100101" => rgb <= "000000";
					when "00010111001100110" => rgb <= "000000";
					when "00010111001100111" => rgb <= "000000";
					when "00010111001101000" => rgb <= "000000";
					when "00010111001101001" => rgb <= "000000";
					when "00010111001101010" => rgb <= "000000";
					when "00010111001101011" => rgb <= "000000";
					when "00010111001101100" => rgb <= "000000";
					when "00010111001101101" => rgb <= "000000";
					when "00010111001101110" => rgb <= "000000";
					when "00010111001101111" => rgb <= "000000";
					when "00010111001110000" => rgb <= "000000";
					when "00010111001110001" => rgb <= "000000";
					when "00010111001110010" => rgb <= "000000";
					when "00010111001110011" => rgb <= "000000";
					when "00010111001110100" => rgb <= "000000";
					when "00010111001110101" => rgb <= "000000";
					when "00010111001110110" => rgb <= "000000";
					when "00010111001110111" => rgb <= "000000";
					when "00010111001111000" => rgb <= "000000";
					when "00010111001111001" => rgb <= "000000";
					when "00010111001111010" => rgb <= "000000";
					when "00010111001111011" => rgb <= "000000";
					when "00010111001111100" => rgb <= "000000";
					when "00010111001111101" => rgb <= "101000";
					when "00010111001111110" => rgb <= "101000";
					when "00010111001111111" => rgb <= "101000";
					when "00010111010000000" => rgb <= "101000";
					when "00010111010000001" => rgb <= "101000";
					when "00010111010000010" => rgb <= "101000";
					when "00010111010000011" => rgb <= "101000";
					when "00010111010000100" => rgb <= "101000";
					when "00010111010000101" => rgb <= "101000";
					when "00010111010000110" => rgb <= "101000";
					when "00010111010000111" => rgb <= "101000";
					when "00010111010001000" => rgb <= "101000";
					when "00010111010001001" => rgb <= "101000";
					when "00010111010001010" => rgb <= "101000";
					when "00010111010001011" => rgb <= "101000";
					when "00010111010001100" => rgb <= "101000";
					when "00010111010001101" => rgb <= "101000";
					when "00010111010001110" => rgb <= "101000";
					when "00010111010001111" => rgb <= "101000";
					when "00010111010010000" => rgb <= "101000";
					when "00010111010010001" => rgb <= "101000";
					when "00010111010010010" => rgb <= "101000";
					when "00010111010010011" => rgb <= "101000";
					when "00010111010010100" => rgb <= "101000";
					when "00010111010010101" => rgb <= "101000";
					when "00010111010010110" => rgb <= "101000";
					when "00010111010010111" => rgb <= "101000";
					when "00010111010011000" => rgb <= "101000";
					when "00010111010011001" => rgb <= "101000";
					when "00010111010011010" => rgb <= "101000";
					when "00010111010011011" => rgb <= "101000";
					when "00010111010011100" => rgb <= "101000";
					when "00010111010011101" => rgb <= "101000";
					when "00010111010011110" => rgb <= "101000";
					when "00010111010011111" => rgb <= "101000";
					when "00010111010100000" => rgb <= "101000";
					when "00010111010100001" => rgb <= "101000";
					when "00010111010100010" => rgb <= "101000";
					when "00010111010100011" => rgb <= "101000";
					when "00010111010100100" => rgb <= "101000";
					when "00010111010100101" => rgb <= "101000";
					when "00010111010100110" => rgb <= "101000";
					when "00010111010100111" => rgb <= "101000";
					when "00010111010101000" => rgb <= "101000";
					when "00010111010101001" => rgb <= "101000";
					when "00010111010101010" => rgb <= "101000";
					when "00010111010101011" => rgb <= "101000";
					when "00010111010101100" => rgb <= "101000";
					when "00010111010101101" => rgb <= "101000";
					when "00010111010101110" => rgb <= "101000";
					when "00010111010101111" => rgb <= "101000";
					when "00010111010110000" => rgb <= "101000";
					when "00010111010110001" => rgb <= "101000";
					when "00010111010110010" => rgb <= "101000";
					when "00010111010110011" => rgb <= "101000";
					when "00010111010110100" => rgb <= "101000";
					when "00010111010110101" => rgb <= "101000";
					when "00010111010110110" => rgb <= "101000";
					when "00010111010110111" => rgb <= "101000";
					when "00010111010111000" => rgb <= "101000";
					when "00010111010111001" => rgb <= "101000";
					when "00010111010111010" => rgb <= "101000";
					when "00010111010111011" => rgb <= "101000";
					when "00010111010111100" => rgb <= "101000";
					when "00010111010111101" => rgb <= "101000";
					when "00010111010111110" => rgb <= "101000";
					when "00010111010111111" => rgb <= "101000";
					when "00010111011000000" => rgb <= "101000";
					when "00010111011000001" => rgb <= "000000";
					when "00010111011000010" => rgb <= "000000";
					when "00010111011000011" => rgb <= "000000";
					when "00010111011000100" => rgb <= "000000";
					when "00010111011000101" => rgb <= "000000";
					when "00010111011000110" => rgb <= "000000";
					when "00010111011000111" => rgb <= "000000";
					when "00010111011001000" => rgb <= "000000";
					when "00010111011001001" => rgb <= "000000";
					when "00010111011001010" => rgb <= "000000";
					when "00010111011001011" => rgb <= "000000";
					when "00010111011001100" => rgb <= "000000";
					when "00010111011001101" => rgb <= "000000";
					when "00010111011001110" => rgb <= "000000";
					when "00010111011001111" => rgb <= "000000";
					when "00010111011010000" => rgb <= "000000";
					when "00010111011010001" => rgb <= "000000";
					when "00010111011010010" => rgb <= "000000";
					when "00010111011010011" => rgb <= "000000";
					when "00010111011010100" => rgb <= "000000";
					when "00010111011010101" => rgb <= "000000";
					when "00010111011010110" => rgb <= "000000";
					when "00010111011010111" => rgb <= "000000";
					when "00010111011011000" => rgb <= "000000";
					when "00010111011011001" => rgb <= "000000";
					when "00010111011011010" => rgb <= "000000";
					when "00010111011011011" => rgb <= "000000";
					when "00010111011011100" => rgb <= "000000";
					when "00010111011011101" => rgb <= "000000";
					when "00010111011011110" => rgb <= "000000";
					when "00010111011011111" => rgb <= "000000";
					when "00010111011100000" => rgb <= "000000";
					when "00010111011100001" => rgb <= "000000";
					when "00010111011100010" => rgb <= "000000";
					when "00010111011100011" => rgb <= "000000";
					when "00010111011100100" => rgb <= "000000";
					when "00010111011100101" => rgb <= "000000";
					when "00010111011100110" => rgb <= "000000";
					when "00010111011100111" => rgb <= "000000";
					when "00010111011101000" => rgb <= "000000";
					when "00010111011101001" => rgb <= "000000";
					when "00010111011101010" => rgb <= "000000";
					when "00010111011101011" => rgb <= "000000";
					when "00010111011101100" => rgb <= "000000";
					when "00010111011101101" => rgb <= "000000";
					when "00010111011101110" => rgb <= "000000";
					when "00010111011101111" => rgb <= "000000";
					when "00010111011110000" => rgb <= "000000";
					when "00010111011110001" => rgb <= "000000";
					when "00010111011110010" => rgb <= "000000";
					when "00010111011110011" => rgb <= "000000";
					when "00010111011110100" => rgb <= "000000";
					when "00010111011110101" => rgb <= "000000";
					when "00010111011110110" => rgb <= "000000";
					when "00010111011110111" => rgb <= "000000";
					when "00010111011111000" => rgb <= "000000";
					when "00010111011111001" => rgb <= "000000";
					when "00010111011111010" => rgb <= "000000";
					when "00010111011111011" => rgb <= "000000";
					when "00010111011111100" => rgb <= "000000";
					when "00010111011111101" => rgb <= "000000";
					when "00010111011111110" => rgb <= "000000";
					when "00010111011111111" => rgb <= "000000";
					when "00010111100000000" => rgb <= "000000";
					when "00010111100000001" => rgb <= "000000";
					when "00010111100000010" => rgb <= "000000";
					when "00010111100000011" => rgb <= "000000";
					when "00010111100000100" => rgb <= "000000";
					when "00010111100000101" => rgb <= "000000";
					when "00010111100000110" => rgb <= "000000";
					when "00010111100000111" => rgb <= "000000";
					when "00010111100001000" => rgb <= "000000";
					when "00010111100001001" => rgb <= "000000";
					when "00010111100001010" => rgb <= "000000";
					when "00010111100001011" => rgb <= "000000";
					when "00010111100001100" => rgb <= "000000";
					when "00010111100001101" => rgb <= "000000";
					when "00010111100001110" => rgb <= "000000";
					when "00010111100001111" => rgb <= "000000";
					when "00010111100010000" => rgb <= "000000";
					when "00010111100010001" => rgb <= "000000";
					when "00010111100010010" => rgb <= "000000";
					when "00010111100010011" => rgb <= "000000";
					when "00010111100010100" => rgb <= "000000";
					when "00010111100010101" => rgb <= "000000";
					when "00010111100010110" => rgb <= "000000";
					when "00010111100010111" => rgb <= "000000";
					when "00010111100011000" => rgb <= "000000";
					when "00010111100011001" => rgb <= "000000";
					when "00010111100011010" => rgb <= "000000";
					when "00010111100011011" => rgb <= "000000";
					when "00010111100011100" => rgb <= "000000";
					when "00010111100011101" => rgb <= "000000";
					when "00010111100011110" => rgb <= "000000";
					when "00010111100011111" => rgb <= "000000";
					when "00010111100100000" => rgb <= "000000";
					when "00010111100100001" => rgb <= "000000";
					when "00010111100100010" => rgb <= "000000";
					when "00010111100100011" => rgb <= "000000";
					when "00010111100100100" => rgb <= "000000";
					when "00010111100100101" => rgb <= "000000";
					when "00010111100100110" => rgb <= "000000";
					when "00010111100100111" => rgb <= "000000";
					when "00010111100101000" => rgb <= "000000";
					when "00010111100101001" => rgb <= "000000";
					when "00010111100101010" => rgb <= "000000";
					when "00010111100101011" => rgb <= "000000";
					when "00010111100101100" => rgb <= "000000";
					when "00010111100101101" => rgb <= "000000";
					when "00010111100101110" => rgb <= "000000";
					when "00010111100101111" => rgb <= "000000";
					when "00010111100110000" => rgb <= "000000";
					when "00010111100110001" => rgb <= "000000";
					when "00010111100110010" => rgb <= "000000";
					when "00010111100110011" => rgb <= "000000";
					when "00010111100110100" => rgb <= "000000";
					when "00010111100110101" => rgb <= "000000";
					when "00010111100110110" => rgb <= "000000";
					when "00010111100110111" => rgb <= "000000";
					when "00010111100111000" => rgb <= "000000";
					when "00010111100111001" => rgb <= "000000";
					when "00010111100111010" => rgb <= "000000";
					when "00010111100111011" => rgb <= "000000";
					when "00010111100111100" => rgb <= "000000";
					when "00010111100111101" => rgb <= "000000";
					when "00010111100111110" => rgb <= "000000";
					when "00010111100111111" => rgb <= "000000";
					when "00011000000000000" => rgb <= "000000";
					when "00011000000000001" => rgb <= "000000";
					when "00011000000000010" => rgb <= "000000";
					when "00011000000000011" => rgb <= "000000";
					when "00011000000000100" => rgb <= "000000";
					when "00011000000000101" => rgb <= "000000";
					when "00011000000000110" => rgb <= "000000";
					when "00011000000000111" => rgb <= "000000";
					when "00011000000001000" => rgb <= "000000";
					when "00011000000001001" => rgb <= "000000";
					when "00011000000001010" => rgb <= "000000";
					when "00011000000001011" => rgb <= "000000";
					when "00011000000001100" => rgb <= "000000";
					when "00011000000001101" => rgb <= "000000";
					when "00011000000001110" => rgb <= "000000";
					when "00011000000001111" => rgb <= "000000";
					when "00011000000010000" => rgb <= "000000";
					when "00011000000010001" => rgb <= "000000";
					when "00011000000010010" => rgb <= "000000";
					when "00011000000010011" => rgb <= "000000";
					when "00011000000010100" => rgb <= "000000";
					when "00011000000010101" => rgb <= "000000";
					when "00011000000010110" => rgb <= "000000";
					when "00011000000010111" => rgb <= "000000";
					when "00011000000011000" => rgb <= "000000";
					when "00011000000011001" => rgb <= "000000";
					when "00011000000011010" => rgb <= "000000";
					when "00011000000011011" => rgb <= "000000";
					when "00011000000011100" => rgb <= "000000";
					when "00011000000011101" => rgb <= "000000";
					when "00011000000011110" => rgb <= "000000";
					when "00011000000011111" => rgb <= "000000";
					when "00011000000100000" => rgb <= "000000";
					when "00011000000100001" => rgb <= "000000";
					when "00011000000100010" => rgb <= "000000";
					when "00011000000100011" => rgb <= "000000";
					when "00011000000100100" => rgb <= "000000";
					when "00011000000100101" => rgb <= "000000";
					when "00011000000100110" => rgb <= "000000";
					when "00011000000100111" => rgb <= "000000";
					when "00011000000101000" => rgb <= "000000";
					when "00011000000101001" => rgb <= "000000";
					when "00011000000101010" => rgb <= "000000";
					when "00011000000101011" => rgb <= "000000";
					when "00011000000101100" => rgb <= "000000";
					when "00011000000101101" => rgb <= "000000";
					when "00011000000101110" => rgb <= "000000";
					when "00011000000101111" => rgb <= "000000";
					when "00011000000110000" => rgb <= "000000";
					when "00011000000110001" => rgb <= "000000";
					when "00011000000110010" => rgb <= "000000";
					when "00011000000110011" => rgb <= "000000";
					when "00011000000110100" => rgb <= "000000";
					when "00011000000110101" => rgb <= "000000";
					when "00011000000110110" => rgb <= "000000";
					when "00011000000110111" => rgb <= "000000";
					when "00011000000111000" => rgb <= "000000";
					when "00011000000111001" => rgb <= "000000";
					when "00011000000111010" => rgb <= "000000";
					when "00011000000111011" => rgb <= "000000";
					when "00011000000111100" => rgb <= "000000";
					when "00011000000111101" => rgb <= "000000";
					when "00011000000111110" => rgb <= "000000";
					when "00011000000111111" => rgb <= "000000";
					when "00011000001000000" => rgb <= "000000";
					when "00011000001000001" => rgb <= "000000";
					when "00011000001000010" => rgb <= "000000";
					when "00011000001000011" => rgb <= "000000";
					when "00011000001000100" => rgb <= "000000";
					when "00011000001000101" => rgb <= "000000";
					when "00011000001000110" => rgb <= "000000";
					when "00011000001000111" => rgb <= "000000";
					when "00011000001001000" => rgb <= "000000";
					when "00011000001001001" => rgb <= "000000";
					when "00011000001001010" => rgb <= "000000";
					when "00011000001001011" => rgb <= "000000";
					when "00011000001001100" => rgb <= "000000";
					when "00011000001001101" => rgb <= "000000";
					when "00011000001001110" => rgb <= "000000";
					when "00011000001001111" => rgb <= "000000";
					when "00011000001010000" => rgb <= "000000";
					when "00011000001010001" => rgb <= "000000";
					when "00011000001010010" => rgb <= "000000";
					when "00011000001010011" => rgb <= "000000";
					when "00011000001010100" => rgb <= "000000";
					when "00011000001010101" => rgb <= "000000";
					when "00011000001010110" => rgb <= "000000";
					when "00011000001010111" => rgb <= "000000";
					when "00011000001011000" => rgb <= "000000";
					when "00011000001011001" => rgb <= "000000";
					when "00011000001011010" => rgb <= "000000";
					when "00011000001011011" => rgb <= "000000";
					when "00011000001011100" => rgb <= "000000";
					when "00011000001011101" => rgb <= "000000";
					when "00011000001011110" => rgb <= "000000";
					when "00011000001011111" => rgb <= "000000";
					when "00011000001100000" => rgb <= "000000";
					when "00011000001100001" => rgb <= "000000";
					when "00011000001100010" => rgb <= "000000";
					when "00011000001100011" => rgb <= "000000";
					when "00011000001100100" => rgb <= "000000";
					when "00011000001100101" => rgb <= "000000";
					when "00011000001100110" => rgb <= "000000";
					when "00011000001100111" => rgb <= "000000";
					when "00011000001101000" => rgb <= "000000";
					when "00011000001101001" => rgb <= "000000";
					when "00011000001101010" => rgb <= "000000";
					when "00011000001101011" => rgb <= "000000";
					when "00011000001101100" => rgb <= "000000";
					when "00011000001101101" => rgb <= "000000";
					when "00011000001101110" => rgb <= "000000";
					when "00011000001101111" => rgb <= "000000";
					when "00011000001110000" => rgb <= "000000";
					when "00011000001110001" => rgb <= "000000";
					when "00011000001110010" => rgb <= "000000";
					when "00011000001110011" => rgb <= "000000";
					when "00011000001110100" => rgb <= "000000";
					when "00011000001110101" => rgb <= "000000";
					when "00011000001110110" => rgb <= "000000";
					when "00011000001110111" => rgb <= "000000";
					when "00011000001111000" => rgb <= "000000";
					when "00011000001111001" => rgb <= "000000";
					when "00011000001111010" => rgb <= "000000";
					when "00011000001111011" => rgb <= "000000";
					when "00011000001111100" => rgb <= "000000";
					when "00011000001111101" => rgb <= "101000";
					when "00011000001111110" => rgb <= "101000";
					when "00011000001111111" => rgb <= "101000";
					when "00011000010000000" => rgb <= "101000";
					when "00011000010000001" => rgb <= "101000";
					when "00011000010000010" => rgb <= "101000";
					when "00011000010000011" => rgb <= "101000";
					when "00011000010000100" => rgb <= "101000";
					when "00011000010000101" => rgb <= "101000";
					when "00011000010000110" => rgb <= "101000";
					when "00011000010000111" => rgb <= "101000";
					when "00011000010001000" => rgb <= "101000";
					when "00011000010001001" => rgb <= "101000";
					when "00011000010001010" => rgb <= "101000";
					when "00011000010001011" => rgb <= "101000";
					when "00011000010001100" => rgb <= "101000";
					when "00011000010001101" => rgb <= "101000";
					when "00011000010001110" => rgb <= "101000";
					when "00011000010001111" => rgb <= "101000";
					when "00011000010010000" => rgb <= "101000";
					when "00011000010010001" => rgb <= "101000";
					when "00011000010010010" => rgb <= "101000";
					when "00011000010010011" => rgb <= "101000";
					when "00011000010010100" => rgb <= "101000";
					when "00011000010010101" => rgb <= "101000";
					when "00011000010010110" => rgb <= "101000";
					when "00011000010010111" => rgb <= "101000";
					when "00011000010011000" => rgb <= "101000";
					when "00011000010011001" => rgb <= "101000";
					when "00011000010011010" => rgb <= "101000";
					when "00011000010011011" => rgb <= "101000";
					when "00011000010011100" => rgb <= "101000";
					when "00011000010011101" => rgb <= "101000";
					when "00011000010011110" => rgb <= "101000";
					when "00011000010011111" => rgb <= "101000";
					when "00011000010100000" => rgb <= "101000";
					when "00011000010100001" => rgb <= "101000";
					when "00011000010100010" => rgb <= "101000";
					when "00011000010100011" => rgb <= "101000";
					when "00011000010100100" => rgb <= "101000";
					when "00011000010100101" => rgb <= "101000";
					when "00011000010100110" => rgb <= "101000";
					when "00011000010100111" => rgb <= "101000";
					when "00011000010101000" => rgb <= "101000";
					when "00011000010101001" => rgb <= "101000";
					when "00011000010101010" => rgb <= "101000";
					when "00011000010101011" => rgb <= "101000";
					when "00011000010101100" => rgb <= "101000";
					when "00011000010101101" => rgb <= "101000";
					when "00011000010101110" => rgb <= "101000";
					when "00011000010101111" => rgb <= "101000";
					when "00011000010110000" => rgb <= "101000";
					when "00011000010110001" => rgb <= "101000";
					when "00011000010110010" => rgb <= "101000";
					when "00011000010110011" => rgb <= "101000";
					when "00011000010110100" => rgb <= "101000";
					when "00011000010110101" => rgb <= "101000";
					when "00011000010110110" => rgb <= "101000";
					when "00011000010110111" => rgb <= "101000";
					when "00011000010111000" => rgb <= "101000";
					when "00011000010111001" => rgb <= "101000";
					when "00011000010111010" => rgb <= "101000";
					when "00011000010111011" => rgb <= "101000";
					when "00011000010111100" => rgb <= "101000";
					when "00011000010111101" => rgb <= "101000";
					when "00011000010111110" => rgb <= "101000";
					when "00011000010111111" => rgb <= "101000";
					when "00011000011000000" => rgb <= "100100";
					when "00011000011000001" => rgb <= "000000";
					when "00011000011000010" => rgb <= "000000";
					when "00011000011000011" => rgb <= "000000";
					when "00011000011000100" => rgb <= "000000";
					when "00011000011000101" => rgb <= "000000";
					when "00011000011000110" => rgb <= "000000";
					when "00011000011000111" => rgb <= "000000";
					when "00011000011001000" => rgb <= "000000";
					when "00011000011001001" => rgb <= "000000";
					when "00011000011001010" => rgb <= "000000";
					when "00011000011001011" => rgb <= "000000";
					when "00011000011001100" => rgb <= "000000";
					when "00011000011001101" => rgb <= "000000";
					when "00011000011001110" => rgb <= "000000";
					when "00011000011001111" => rgb <= "000000";
					when "00011000011010000" => rgb <= "000000";
					when "00011000011010001" => rgb <= "000000";
					when "00011000011010010" => rgb <= "000000";
					when "00011000011010011" => rgb <= "000000";
					when "00011000011010100" => rgb <= "000000";
					when "00011000011010101" => rgb <= "000000";
					when "00011000011010110" => rgb <= "000000";
					when "00011000011010111" => rgb <= "000000";
					when "00011000011011000" => rgb <= "000000";
					when "00011000011011001" => rgb <= "000000";
					when "00011000011011010" => rgb <= "000000";
					when "00011000011011011" => rgb <= "000000";
					when "00011000011011100" => rgb <= "000000";
					when "00011000011011101" => rgb <= "000000";
					when "00011000011011110" => rgb <= "000000";
					when "00011000011011111" => rgb <= "000000";
					when "00011000011100000" => rgb <= "000000";
					when "00011000011100001" => rgb <= "000000";
					when "00011000011100010" => rgb <= "000000";
					when "00011000011100011" => rgb <= "000000";
					when "00011000011100100" => rgb <= "000000";
					when "00011000011100101" => rgb <= "000000";
					when "00011000011100110" => rgb <= "000000";
					when "00011000011100111" => rgb <= "000000";
					when "00011000011101000" => rgb <= "000000";
					when "00011000011101001" => rgb <= "000000";
					when "00011000011101010" => rgb <= "000000";
					when "00011000011101011" => rgb <= "000000";
					when "00011000011101100" => rgb <= "000000";
					when "00011000011101101" => rgb <= "000000";
					when "00011000011101110" => rgb <= "000000";
					when "00011000011101111" => rgb <= "000000";
					when "00011000011110000" => rgb <= "000000";
					when "00011000011110001" => rgb <= "000000";
					when "00011000011110010" => rgb <= "000000";
					when "00011000011110011" => rgb <= "000000";
					when "00011000011110100" => rgb <= "000000";
					when "00011000011110101" => rgb <= "000000";
					when "00011000011110110" => rgb <= "000000";
					when "00011000011110111" => rgb <= "000000";
					when "00011000011111000" => rgb <= "000000";
					when "00011000011111001" => rgb <= "000000";
					when "00011000011111010" => rgb <= "000000";
					when "00011000011111011" => rgb <= "000000";
					when "00011000011111100" => rgb <= "000000";
					when "00011000011111101" => rgb <= "000000";
					when "00011000011111110" => rgb <= "000000";
					when "00011000011111111" => rgb <= "000000";
					when "00011000100000000" => rgb <= "000000";
					when "00011000100000001" => rgb <= "000000";
					when "00011000100000010" => rgb <= "000000";
					when "00011000100000011" => rgb <= "000000";
					when "00011000100000100" => rgb <= "000000";
					when "00011000100000101" => rgb <= "000000";
					when "00011000100000110" => rgb <= "000000";
					when "00011000100000111" => rgb <= "000000";
					when "00011000100001000" => rgb <= "000000";
					when "00011000100001001" => rgb <= "000000";
					when "00011000100001010" => rgb <= "000000";
					when "00011000100001011" => rgb <= "000000";
					when "00011000100001100" => rgb <= "000000";
					when "00011000100001101" => rgb <= "000000";
					when "00011000100001110" => rgb <= "000000";
					when "00011000100001111" => rgb <= "000000";
					when "00011000100010000" => rgb <= "000000";
					when "00011000100010001" => rgb <= "000000";
					when "00011000100010010" => rgb <= "000000";
					when "00011000100010011" => rgb <= "000000";
					when "00011000100010100" => rgb <= "000000";
					when "00011000100010101" => rgb <= "000000";
					when "00011000100010110" => rgb <= "000000";
					when "00011000100010111" => rgb <= "000000";
					when "00011000100011000" => rgb <= "000000";
					when "00011000100011001" => rgb <= "000000";
					when "00011000100011010" => rgb <= "000000";
					when "00011000100011011" => rgb <= "000000";
					when "00011000100011100" => rgb <= "000000";
					when "00011000100011101" => rgb <= "000000";
					when "00011000100011110" => rgb <= "000000";
					when "00011000100011111" => rgb <= "000000";
					when "00011000100100000" => rgb <= "000000";
					when "00011000100100001" => rgb <= "000000";
					when "00011000100100010" => rgb <= "000000";
					when "00011000100100011" => rgb <= "000000";
					when "00011000100100100" => rgb <= "000000";
					when "00011000100100101" => rgb <= "000000";
					when "00011000100100110" => rgb <= "000000";
					when "00011000100100111" => rgb <= "000000";
					when "00011000100101000" => rgb <= "000000";
					when "00011000100101001" => rgb <= "000000";
					when "00011000100101010" => rgb <= "000000";
					when "00011000100101011" => rgb <= "000000";
					when "00011000100101100" => rgb <= "000000";
					when "00011000100101101" => rgb <= "000000";
					when "00011000100101110" => rgb <= "000000";
					when "00011000100101111" => rgb <= "000000";
					when "00011000100110000" => rgb <= "000000";
					when "00011000100110001" => rgb <= "000000";
					when "00011000100110010" => rgb <= "000000";
					when "00011000100110011" => rgb <= "000000";
					when "00011000100110100" => rgb <= "000000";
					when "00011000100110101" => rgb <= "000000";
					when "00011000100110110" => rgb <= "000000";
					when "00011000100110111" => rgb <= "000000";
					when "00011000100111000" => rgb <= "000000";
					when "00011000100111001" => rgb <= "000000";
					when "00011000100111010" => rgb <= "000000";
					when "00011000100111011" => rgb <= "000000";
					when "00011000100111100" => rgb <= "000000";
					when "00011000100111101" => rgb <= "000000";
					when "00011000100111110" => rgb <= "000000";
					when "00011000100111111" => rgb <= "000000";
					when "00011001000000000" => rgb <= "000000";
					when "00011001000000001" => rgb <= "000000";
					when "00011001000000010" => rgb <= "000000";
					when "00011001000000011" => rgb <= "000000";
					when "00011001000000100" => rgb <= "000000";
					when "00011001000000101" => rgb <= "000000";
					when "00011001000000110" => rgb <= "000000";
					when "00011001000000111" => rgb <= "000000";
					when "00011001000001000" => rgb <= "000000";
					when "00011001000001001" => rgb <= "000000";
					when "00011001000001010" => rgb <= "000000";
					when "00011001000001011" => rgb <= "000000";
					when "00011001000001100" => rgb <= "000000";
					when "00011001000001101" => rgb <= "000000";
					when "00011001000001110" => rgb <= "000000";
					when "00011001000001111" => rgb <= "000000";
					when "00011001000010000" => rgb <= "000000";
					when "00011001000010001" => rgb <= "000000";
					when "00011001000010010" => rgb <= "000000";
					when "00011001000010011" => rgb <= "000000";
					when "00011001000010100" => rgb <= "000000";
					when "00011001000010101" => rgb <= "000000";
					when "00011001000010110" => rgb <= "000000";
					when "00011001000010111" => rgb <= "000000";
					when "00011001000011000" => rgb <= "000000";
					when "00011001000011001" => rgb <= "000000";
					when "00011001000011010" => rgb <= "000000";
					when "00011001000011011" => rgb <= "000000";
					when "00011001000011100" => rgb <= "000000";
					when "00011001000011101" => rgb <= "000000";
					when "00011001000011110" => rgb <= "000000";
					when "00011001000011111" => rgb <= "000000";
					when "00011001000100000" => rgb <= "000000";
					when "00011001000100001" => rgb <= "000000";
					when "00011001000100010" => rgb <= "000000";
					when "00011001000100011" => rgb <= "000000";
					when "00011001000100100" => rgb <= "000000";
					when "00011001000100101" => rgb <= "000000";
					when "00011001000100110" => rgb <= "000000";
					when "00011001000100111" => rgb <= "000000";
					when "00011001000101000" => rgb <= "000000";
					when "00011001000101001" => rgb <= "000000";
					when "00011001000101010" => rgb <= "000000";
					when "00011001000101011" => rgb <= "000000";
					when "00011001000101100" => rgb <= "000000";
					when "00011001000101101" => rgb <= "000000";
					when "00011001000101110" => rgb <= "000000";
					when "00011001000101111" => rgb <= "000000";
					when "00011001000110000" => rgb <= "000000";
					when "00011001000110001" => rgb <= "000000";
					when "00011001000110010" => rgb <= "000000";
					when "00011001000110011" => rgb <= "000000";
					when "00011001000110100" => rgb <= "000000";
					when "00011001000110101" => rgb <= "000000";
					when "00011001000110110" => rgb <= "000000";
					when "00011001000110111" => rgb <= "000000";
					when "00011001000111000" => rgb <= "000000";
					when "00011001000111001" => rgb <= "000000";
					when "00011001000111010" => rgb <= "000000";
					when "00011001000111011" => rgb <= "000000";
					when "00011001000111100" => rgb <= "000000";
					when "00011001000111101" => rgb <= "000000";
					when "00011001000111110" => rgb <= "000000";
					when "00011001000111111" => rgb <= "000000";
					when "00011001001000000" => rgb <= "000000";
					when "00011001001000001" => rgb <= "000000";
					when "00011001001000010" => rgb <= "000000";
					when "00011001001000011" => rgb <= "000000";
					when "00011001001000100" => rgb <= "000000";
					when "00011001001000101" => rgb <= "000000";
					when "00011001001000110" => rgb <= "000000";
					when "00011001001000111" => rgb <= "000000";
					when "00011001001001000" => rgb <= "000000";
					when "00011001001001001" => rgb <= "000000";
					when "00011001001001010" => rgb <= "000000";
					when "00011001001001011" => rgb <= "000000";
					when "00011001001001100" => rgb <= "000000";
					when "00011001001001101" => rgb <= "000000";
					when "00011001001001110" => rgb <= "000000";
					when "00011001001001111" => rgb <= "000000";
					when "00011001001010000" => rgb <= "000000";
					when "00011001001010001" => rgb <= "000000";
					when "00011001001010010" => rgb <= "000000";
					when "00011001001010011" => rgb <= "000000";
					when "00011001001010100" => rgb <= "000000";
					when "00011001001010101" => rgb <= "000000";
					when "00011001001010110" => rgb <= "000000";
					when "00011001001010111" => rgb <= "000000";
					when "00011001001011000" => rgb <= "000000";
					when "00011001001011001" => rgb <= "000000";
					when "00011001001011010" => rgb <= "000000";
					when "00011001001011011" => rgb <= "000000";
					when "00011001001011100" => rgb <= "000000";
					when "00011001001011101" => rgb <= "000000";
					when "00011001001011110" => rgb <= "000000";
					when "00011001001011111" => rgb <= "000000";
					when "00011001001100000" => rgb <= "000000";
					when "00011001001100001" => rgb <= "000000";
					when "00011001001100010" => rgb <= "000000";
					when "00011001001100011" => rgb <= "000000";
					when "00011001001100100" => rgb <= "000000";
					when "00011001001100101" => rgb <= "000000";
					when "00011001001100110" => rgb <= "000000";
					when "00011001001100111" => rgb <= "000000";
					when "00011001001101000" => rgb <= "000000";
					when "00011001001101001" => rgb <= "000000";
					when "00011001001101010" => rgb <= "000000";
					when "00011001001101011" => rgb <= "000000";
					when "00011001001101100" => rgb <= "000000";
					when "00011001001101101" => rgb <= "000000";
					when "00011001001101110" => rgb <= "000000";
					when "00011001001101111" => rgb <= "000000";
					when "00011001001110000" => rgb <= "000000";
					when "00011001001110001" => rgb <= "000000";
					when "00011001001110010" => rgb <= "000000";
					when "00011001001110011" => rgb <= "000000";
					when "00011001001110100" => rgb <= "000000";
					when "00011001001110101" => rgb <= "000000";
					when "00011001001110110" => rgb <= "000000";
					when "00011001001110111" => rgb <= "000000";
					when "00011001001111000" => rgb <= "000000";
					when "00011001001111001" => rgb <= "000000";
					when "00011001001111010" => rgb <= "000000";
					when "00011001001111011" => rgb <= "000000";
					when "00011001001111100" => rgb <= "000000";
					when "00011001001111101" => rgb <= "101000";
					when "00011001001111110" => rgb <= "101000";
					when "00011001001111111" => rgb <= "101000";
					when "00011001010000000" => rgb <= "101000";
					when "00011001010000001" => rgb <= "101000";
					when "00011001010000010" => rgb <= "101000";
					when "00011001010000011" => rgb <= "101000";
					when "00011001010000100" => rgb <= "101000";
					when "00011001010000101" => rgb <= "101000";
					when "00011001010000110" => rgb <= "101000";
					when "00011001010000111" => rgb <= "101000";
					when "00011001010001000" => rgb <= "101000";
					when "00011001010001001" => rgb <= "101000";
					when "00011001010001010" => rgb <= "101000";
					when "00011001010001011" => rgb <= "101000";
					when "00011001010001100" => rgb <= "101000";
					when "00011001010001101" => rgb <= "101000";
					when "00011001010001110" => rgb <= "101000";
					when "00011001010001111" => rgb <= "101000";
					when "00011001010010000" => rgb <= "101000";
					when "00011001010010001" => rgb <= "101000";
					when "00011001010010010" => rgb <= "101000";
					when "00011001010010011" => rgb <= "101000";
					when "00011001010010100" => rgb <= "101000";
					when "00011001010010101" => rgb <= "101000";
					when "00011001010010110" => rgb <= "101000";
					when "00011001010010111" => rgb <= "101000";
					when "00011001010011000" => rgb <= "101000";
					when "00011001010011001" => rgb <= "101000";
					when "00011001010011010" => rgb <= "101000";
					when "00011001010011011" => rgb <= "101000";
					when "00011001010011100" => rgb <= "101000";
					when "00011001010011101" => rgb <= "101000";
					when "00011001010011110" => rgb <= "101000";
					when "00011001010011111" => rgb <= "101000";
					when "00011001010100000" => rgb <= "101000";
					when "00011001010100001" => rgb <= "101000";
					when "00011001010100010" => rgb <= "101000";
					when "00011001010100011" => rgb <= "101000";
					when "00011001010100100" => rgb <= "101000";
					when "00011001010100101" => rgb <= "101000";
					when "00011001010100110" => rgb <= "101000";
					when "00011001010100111" => rgb <= "101000";
					when "00011001010101000" => rgb <= "101000";
					when "00011001010101001" => rgb <= "101000";
					when "00011001010101010" => rgb <= "101000";
					when "00011001010101011" => rgb <= "101000";
					when "00011001010101100" => rgb <= "101000";
					when "00011001010101101" => rgb <= "101000";
					when "00011001010101110" => rgb <= "101000";
					when "00011001010101111" => rgb <= "101000";
					when "00011001010110000" => rgb <= "101000";
					when "00011001010110001" => rgb <= "101000";
					when "00011001010110010" => rgb <= "101000";
					when "00011001010110011" => rgb <= "101000";
					when "00011001010110100" => rgb <= "101000";
					when "00011001010110101" => rgb <= "101000";
					when "00011001010110110" => rgb <= "101000";
					when "00011001010110111" => rgb <= "101000";
					when "00011001010111000" => rgb <= "101000";
					when "00011001010111001" => rgb <= "101000";
					when "00011001010111010" => rgb <= "101000";
					when "00011001010111011" => rgb <= "101000";
					when "00011001010111100" => rgb <= "101000";
					when "00011001010111101" => rgb <= "101000";
					when "00011001010111110" => rgb <= "101000";
					when "00011001010111111" => rgb <= "101000";
					when "00011001011000000" => rgb <= "100100";
					when "00011001011000001" => rgb <= "000000";
					when "00011001011000010" => rgb <= "000000";
					when "00011001011000011" => rgb <= "000000";
					when "00011001011000100" => rgb <= "000000";
					when "00011001011000101" => rgb <= "000000";
					when "00011001011000110" => rgb <= "000000";
					when "00011001011000111" => rgb <= "000000";
					when "00011001011001000" => rgb <= "000000";
					when "00011001011001001" => rgb <= "000000";
					when "00011001011001010" => rgb <= "000000";
					when "00011001011001011" => rgb <= "000000";
					when "00011001011001100" => rgb <= "000000";
					when "00011001011001101" => rgb <= "000000";
					when "00011001011001110" => rgb <= "000000";
					when "00011001011001111" => rgb <= "000000";
					when "00011001011010000" => rgb <= "000000";
					when "00011001011010001" => rgb <= "000000";
					when "00011001011010010" => rgb <= "000000";
					when "00011001011010011" => rgb <= "000000";
					when "00011001011010100" => rgb <= "000000";
					when "00011001011010101" => rgb <= "000000";
					when "00011001011010110" => rgb <= "000000";
					when "00011001011010111" => rgb <= "000000";
					when "00011001011011000" => rgb <= "000000";
					when "00011001011011001" => rgb <= "000000";
					when "00011001011011010" => rgb <= "000000";
					when "00011001011011011" => rgb <= "000000";
					when "00011001011011100" => rgb <= "000000";
					when "00011001011011101" => rgb <= "000000";
					when "00011001011011110" => rgb <= "000000";
					when "00011001011011111" => rgb <= "000000";
					when "00011001011100000" => rgb <= "000000";
					when "00011001011100001" => rgb <= "000000";
					when "00011001011100010" => rgb <= "000000";
					when "00011001011100011" => rgb <= "000000";
					when "00011001011100100" => rgb <= "000000";
					when "00011001011100101" => rgb <= "000000";
					when "00011001011100110" => rgb <= "000000";
					when "00011001011100111" => rgb <= "000000";
					when "00011001011101000" => rgb <= "000000";
					when "00011001011101001" => rgb <= "000000";
					when "00011001011101010" => rgb <= "000000";
					when "00011001011101011" => rgb <= "000000";
					when "00011001011101100" => rgb <= "000000";
					when "00011001011101101" => rgb <= "000000";
					when "00011001011101110" => rgb <= "000000";
					when "00011001011101111" => rgb <= "000000";
					when "00011001011110000" => rgb <= "000000";
					when "00011001011110001" => rgb <= "000000";
					when "00011001011110010" => rgb <= "000000";
					when "00011001011110011" => rgb <= "000000";
					when "00011001011110100" => rgb <= "000000";
					when "00011001011110101" => rgb <= "000000";
					when "00011001011110110" => rgb <= "000000";
					when "00011001011110111" => rgb <= "000000";
					when "00011001011111000" => rgb <= "000000";
					when "00011001011111001" => rgb <= "000000";
					when "00011001011111010" => rgb <= "000000";
					when "00011001011111011" => rgb <= "000000";
					when "00011001011111100" => rgb <= "000000";
					when "00011001011111101" => rgb <= "000000";
					when "00011001011111110" => rgb <= "000000";
					when "00011001011111111" => rgb <= "000000";
					when "00011001100000000" => rgb <= "000000";
					when "00011001100000001" => rgb <= "000000";
					when "00011001100000010" => rgb <= "000000";
					when "00011001100000011" => rgb <= "000000";
					when "00011001100000100" => rgb <= "000000";
					when "00011001100000101" => rgb <= "000000";
					when "00011001100000110" => rgb <= "000000";
					when "00011001100000111" => rgb <= "000000";
					when "00011001100001000" => rgb <= "000000";
					when "00011001100001001" => rgb <= "000000";
					when "00011001100001010" => rgb <= "000000";
					when "00011001100001011" => rgb <= "000000";
					when "00011001100001100" => rgb <= "000000";
					when "00011001100001101" => rgb <= "000000";
					when "00011001100001110" => rgb <= "000000";
					when "00011001100001111" => rgb <= "000000";
					when "00011001100010000" => rgb <= "000000";
					when "00011001100010001" => rgb <= "000000";
					when "00011001100010010" => rgb <= "000000";
					when "00011001100010011" => rgb <= "000000";
					when "00011001100010100" => rgb <= "000000";
					when "00011001100010101" => rgb <= "000000";
					when "00011001100010110" => rgb <= "000000";
					when "00011001100010111" => rgb <= "000000";
					when "00011001100011000" => rgb <= "000000";
					when "00011001100011001" => rgb <= "000000";
					when "00011001100011010" => rgb <= "000000";
					when "00011001100011011" => rgb <= "000000";
					when "00011001100011100" => rgb <= "000000";
					when "00011001100011101" => rgb <= "000000";
					when "00011001100011110" => rgb <= "000000";
					when "00011001100011111" => rgb <= "000000";
					when "00011001100100000" => rgb <= "000000";
					when "00011001100100001" => rgb <= "000000";
					when "00011001100100010" => rgb <= "000000";
					when "00011001100100011" => rgb <= "000000";
					when "00011001100100100" => rgb <= "000000";
					when "00011001100100101" => rgb <= "000000";
					when "00011001100100110" => rgb <= "000000";
					when "00011001100100111" => rgb <= "000000";
					when "00011001100101000" => rgb <= "000000";
					when "00011001100101001" => rgb <= "000000";
					when "00011001100101010" => rgb <= "000000";
					when "00011001100101011" => rgb <= "000000";
					when "00011001100101100" => rgb <= "000000";
					when "00011001100101101" => rgb <= "000000";
					when "00011001100101110" => rgb <= "000000";
					when "00011001100101111" => rgb <= "000000";
					when "00011001100110000" => rgb <= "000000";
					when "00011001100110001" => rgb <= "000000";
					when "00011001100110010" => rgb <= "000000";
					when "00011001100110011" => rgb <= "000000";
					when "00011001100110100" => rgb <= "000000";
					when "00011001100110101" => rgb <= "000000";
					when "00011001100110110" => rgb <= "000000";
					when "00011001100110111" => rgb <= "000000";
					when "00011001100111000" => rgb <= "000000";
					when "00011001100111001" => rgb <= "000000";
					when "00011001100111010" => rgb <= "000000";
					when "00011001100111011" => rgb <= "000000";
					when "00011001100111100" => rgb <= "000000";
					when "00011001100111101" => rgb <= "000000";
					when "00011001100111110" => rgb <= "000000";
					when "00011001100111111" => rgb <= "000000";
					when "00011010000000000" => rgb <= "000000";
					when "00011010000000001" => rgb <= "000000";
					when "00011010000000010" => rgb <= "000000";
					when "00011010000000011" => rgb <= "000000";
					when "00011010000000100" => rgb <= "000000";
					when "00011010000000101" => rgb <= "000000";
					when "00011010000000110" => rgb <= "000000";
					when "00011010000000111" => rgb <= "000000";
					when "00011010000001000" => rgb <= "000000";
					when "00011010000001001" => rgb <= "000000";
					when "00011010000001010" => rgb <= "000000";
					when "00011010000001011" => rgb <= "000000";
					when "00011010000001100" => rgb <= "000000";
					when "00011010000001101" => rgb <= "000000";
					when "00011010000001110" => rgb <= "000000";
					when "00011010000001111" => rgb <= "000000";
					when "00011010000010000" => rgb <= "000000";
					when "00011010000010001" => rgb <= "000000";
					when "00011010000010010" => rgb <= "000000";
					when "00011010000010011" => rgb <= "000000";
					when "00011010000010100" => rgb <= "000000";
					when "00011010000010101" => rgb <= "000000";
					when "00011010000010110" => rgb <= "000000";
					when "00011010000010111" => rgb <= "000000";
					when "00011010000011000" => rgb <= "000000";
					when "00011010000011001" => rgb <= "000000";
					when "00011010000011010" => rgb <= "000000";
					when "00011010000011011" => rgb <= "000000";
					when "00011010000011100" => rgb <= "000000";
					when "00011010000011101" => rgb <= "000000";
					when "00011010000011110" => rgb <= "000000";
					when "00011010000011111" => rgb <= "000000";
					when "00011010000100000" => rgb <= "000000";
					when "00011010000100001" => rgb <= "000000";
					when "00011010000100010" => rgb <= "000000";
					when "00011010000100011" => rgb <= "000000";
					when "00011010000100100" => rgb <= "000000";
					when "00011010000100101" => rgb <= "000000";
					when "00011010000100110" => rgb <= "000000";
					when "00011010000100111" => rgb <= "000000";
					when "00011010000101000" => rgb <= "000000";
					when "00011010000101001" => rgb <= "000000";
					when "00011010000101010" => rgb <= "000000";
					when "00011010000101011" => rgb <= "000000";
					when "00011010000101100" => rgb <= "000000";
					when "00011010000101101" => rgb <= "000000";
					when "00011010000101110" => rgb <= "000000";
					when "00011010000101111" => rgb <= "000000";
					when "00011010000110000" => rgb <= "000000";
					when "00011010000110001" => rgb <= "000000";
					when "00011010000110010" => rgb <= "000000";
					when "00011010000110011" => rgb <= "000000";
					when "00011010000110100" => rgb <= "000000";
					when "00011010000110101" => rgb <= "000000";
					when "00011010000110110" => rgb <= "000000";
					when "00011010000110111" => rgb <= "000000";
					when "00011010000111000" => rgb <= "000000";
					when "00011010000111001" => rgb <= "000000";
					when "00011010000111010" => rgb <= "000000";
					when "00011010000111011" => rgb <= "000000";
					when "00011010000111100" => rgb <= "000000";
					when "00011010000111101" => rgb <= "000000";
					when "00011010000111110" => rgb <= "000000";
					when "00011010000111111" => rgb <= "000000";
					when "00011010001000000" => rgb <= "000000";
					when "00011010001000001" => rgb <= "000000";
					when "00011010001000010" => rgb <= "000000";
					when "00011010001000011" => rgb <= "000000";
					when "00011010001000100" => rgb <= "000000";
					when "00011010001000101" => rgb <= "000000";
					when "00011010001000110" => rgb <= "000000";
					when "00011010001000111" => rgb <= "000000";
					when "00011010001001000" => rgb <= "000000";
					when "00011010001001001" => rgb <= "000000";
					when "00011010001001010" => rgb <= "000000";
					when "00011010001001011" => rgb <= "000000";
					when "00011010001001100" => rgb <= "000000";
					when "00011010001001101" => rgb <= "000000";
					when "00011010001001110" => rgb <= "000000";
					when "00011010001001111" => rgb <= "000000";
					when "00011010001010000" => rgb <= "000000";
					when "00011010001010001" => rgb <= "000000";
					when "00011010001010010" => rgb <= "000000";
					when "00011010001010011" => rgb <= "000000";
					when "00011010001010100" => rgb <= "000000";
					when "00011010001010101" => rgb <= "000000";
					when "00011010001010110" => rgb <= "000000";
					when "00011010001010111" => rgb <= "000000";
					when "00011010001011000" => rgb <= "000000";
					when "00011010001011001" => rgb <= "000000";
					when "00011010001011010" => rgb <= "000000";
					when "00011010001011011" => rgb <= "000000";
					when "00011010001011100" => rgb <= "000000";
					when "00011010001011101" => rgb <= "000000";
					when "00011010001011110" => rgb <= "000000";
					when "00011010001011111" => rgb <= "000000";
					when "00011010001100000" => rgb <= "000000";
					when "00011010001100001" => rgb <= "000000";
					when "00011010001100010" => rgb <= "000000";
					when "00011010001100011" => rgb <= "000000";
					when "00011010001100100" => rgb <= "000000";
					when "00011010001100101" => rgb <= "000000";
					when "00011010001100110" => rgb <= "000000";
					when "00011010001100111" => rgb <= "000000";
					when "00011010001101000" => rgb <= "000000";
					when "00011010001101001" => rgb <= "000000";
					when "00011010001101010" => rgb <= "000000";
					when "00011010001101011" => rgb <= "000000";
					when "00011010001101100" => rgb <= "000000";
					when "00011010001101101" => rgb <= "000000";
					when "00011010001101110" => rgb <= "000000";
					when "00011010001101111" => rgb <= "000000";
					when "00011010001110000" => rgb <= "000000";
					when "00011010001110001" => rgb <= "000000";
					when "00011010001110010" => rgb <= "000000";
					when "00011010001110011" => rgb <= "000000";
					when "00011010001110100" => rgb <= "000000";
					when "00011010001110101" => rgb <= "000000";
					when "00011010001110110" => rgb <= "000000";
					when "00011010001110111" => rgb <= "000000";
					when "00011010001111000" => rgb <= "000000";
					when "00011010001111001" => rgb <= "000000";
					when "00011010001111010" => rgb <= "000000";
					when "00011010001111011" => rgb <= "000000";
					when "00011010001111100" => rgb <= "000000";
					when "00011010001111101" => rgb <= "101000";
					when "00011010001111110" => rgb <= "101000";
					when "00011010001111111" => rgb <= "101000";
					when "00011010010000000" => rgb <= "101000";
					when "00011010010000001" => rgb <= "101000";
					when "00011010010000010" => rgb <= "101000";
					when "00011010010000011" => rgb <= "101000";
					when "00011010010000100" => rgb <= "101000";
					when "00011010010000101" => rgb <= "101000";
					when "00011010010000110" => rgb <= "101000";
					when "00011010010000111" => rgb <= "101000";
					when "00011010010001000" => rgb <= "101000";
					when "00011010010001001" => rgb <= "101000";
					when "00011010010001010" => rgb <= "101000";
					when "00011010010001011" => rgb <= "101000";
					when "00011010010001100" => rgb <= "101000";
					when "00011010010001101" => rgb <= "101000";
					when "00011010010001110" => rgb <= "101000";
					when "00011010010001111" => rgb <= "101000";
					when "00011010010010000" => rgb <= "101000";
					when "00011010010010001" => rgb <= "101000";
					when "00011010010010010" => rgb <= "101000";
					when "00011010010010011" => rgb <= "101000";
					when "00011010010010100" => rgb <= "101000";
					when "00011010010010101" => rgb <= "101000";
					when "00011010010010110" => rgb <= "101000";
					when "00011010010010111" => rgb <= "101000";
					when "00011010010011000" => rgb <= "101000";
					when "00011010010011001" => rgb <= "101000";
					when "00011010010011010" => rgb <= "101000";
					when "00011010010011011" => rgb <= "101000";
					when "00011010010011100" => rgb <= "101000";
					when "00011010010011101" => rgb <= "101000";
					when "00011010010011110" => rgb <= "101000";
					when "00011010010011111" => rgb <= "101000";
					when "00011010010100000" => rgb <= "101000";
					when "00011010010100001" => rgb <= "101000";
					when "00011010010100010" => rgb <= "101000";
					when "00011010010100011" => rgb <= "101000";
					when "00011010010100100" => rgb <= "101000";
					when "00011010010100101" => rgb <= "101000";
					when "00011010010100110" => rgb <= "101000";
					when "00011010010100111" => rgb <= "101000";
					when "00011010010101000" => rgb <= "101000";
					when "00011010010101001" => rgb <= "101000";
					when "00011010010101010" => rgb <= "101000";
					when "00011010010101011" => rgb <= "101000";
					when "00011010010101100" => rgb <= "101000";
					when "00011010010101101" => rgb <= "101000";
					when "00011010010101110" => rgb <= "101000";
					when "00011010010101111" => rgb <= "101000";
					when "00011010010110000" => rgb <= "101000";
					when "00011010010110001" => rgb <= "101000";
					when "00011010010110010" => rgb <= "101000";
					when "00011010010110011" => rgb <= "101000";
					when "00011010010110100" => rgb <= "101000";
					when "00011010010110101" => rgb <= "101000";
					when "00011010010110110" => rgb <= "101000";
					when "00011010010110111" => rgb <= "101000";
					when "00011010010111000" => rgb <= "101000";
					when "00011010010111001" => rgb <= "101000";
					when "00011010010111010" => rgb <= "101000";
					when "00011010010111011" => rgb <= "101000";
					when "00011010010111100" => rgb <= "101000";
					when "00011010010111101" => rgb <= "101000";
					when "00011010010111110" => rgb <= "101000";
					when "00011010010111111" => rgb <= "101000";
					when "00011010011000000" => rgb <= "100100";
					when "00011010011000001" => rgb <= "000000";
					when "00011010011000010" => rgb <= "000000";
					when "00011010011000011" => rgb <= "000000";
					when "00011010011000100" => rgb <= "000000";
					when "00011010011000101" => rgb <= "000000";
					when "00011010011000110" => rgb <= "000000";
					when "00011010011000111" => rgb <= "000000";
					when "00011010011001000" => rgb <= "000000";
					when "00011010011001001" => rgb <= "000000";
					when "00011010011001010" => rgb <= "000000";
					when "00011010011001011" => rgb <= "000000";
					when "00011010011001100" => rgb <= "000000";
					when "00011010011001101" => rgb <= "000000";
					when "00011010011001110" => rgb <= "000000";
					when "00011010011001111" => rgb <= "000000";
					when "00011010011010000" => rgb <= "000000";
					when "00011010011010001" => rgb <= "000000";
					when "00011010011010010" => rgb <= "000000";
					when "00011010011010011" => rgb <= "000000";
					when "00011010011010100" => rgb <= "000000";
					when "00011010011010101" => rgb <= "000000";
					when "00011010011010110" => rgb <= "000000";
					when "00011010011010111" => rgb <= "000000";
					when "00011010011011000" => rgb <= "000000";
					when "00011010011011001" => rgb <= "000000";
					when "00011010011011010" => rgb <= "000000";
					when "00011010011011011" => rgb <= "000000";
					when "00011010011011100" => rgb <= "000000";
					when "00011010011011101" => rgb <= "000000";
					when "00011010011011110" => rgb <= "000000";
					when "00011010011011111" => rgb <= "000000";
					when "00011010011100000" => rgb <= "000000";
					when "00011010011100001" => rgb <= "000000";
					when "00011010011100010" => rgb <= "000000";
					when "00011010011100011" => rgb <= "000000";
					when "00011010011100100" => rgb <= "000000";
					when "00011010011100101" => rgb <= "000000";
					when "00011010011100110" => rgb <= "000000";
					when "00011010011100111" => rgb <= "000000";
					when "00011010011101000" => rgb <= "000000";
					when "00011010011101001" => rgb <= "000000";
					when "00011010011101010" => rgb <= "000000";
					when "00011010011101011" => rgb <= "000000";
					when "00011010011101100" => rgb <= "000000";
					when "00011010011101101" => rgb <= "000000";
					when "00011010011101110" => rgb <= "000000";
					when "00011010011101111" => rgb <= "000000";
					when "00011010011110000" => rgb <= "000000";
					when "00011010011110001" => rgb <= "000000";
					when "00011010011110010" => rgb <= "000000";
					when "00011010011110011" => rgb <= "000000";
					when "00011010011110100" => rgb <= "000000";
					when "00011010011110101" => rgb <= "000000";
					when "00011010011110110" => rgb <= "000000";
					when "00011010011110111" => rgb <= "000000";
					when "00011010011111000" => rgb <= "000000";
					when "00011010011111001" => rgb <= "000000";
					when "00011010011111010" => rgb <= "000000";
					when "00011010011111011" => rgb <= "000000";
					when "00011010011111100" => rgb <= "000000";
					when "00011010011111101" => rgb <= "000000";
					when "00011010011111110" => rgb <= "000000";
					when "00011010011111111" => rgb <= "000000";
					when "00011010100000000" => rgb <= "000000";
					when "00011010100000001" => rgb <= "000000";
					when "00011010100000010" => rgb <= "000000";
					when "00011010100000011" => rgb <= "000000";
					when "00011010100000100" => rgb <= "000000";
					when "00011010100000101" => rgb <= "000000";
					when "00011010100000110" => rgb <= "000000";
					when "00011010100000111" => rgb <= "000000";
					when "00011010100001000" => rgb <= "000000";
					when "00011010100001001" => rgb <= "000000";
					when "00011010100001010" => rgb <= "000000";
					when "00011010100001011" => rgb <= "000000";
					when "00011010100001100" => rgb <= "000000";
					when "00011010100001101" => rgb <= "000000";
					when "00011010100001110" => rgb <= "000000";
					when "00011010100001111" => rgb <= "000000";
					when "00011010100010000" => rgb <= "000000";
					when "00011010100010001" => rgb <= "000000";
					when "00011010100010010" => rgb <= "000000";
					when "00011010100010011" => rgb <= "000000";
					when "00011010100010100" => rgb <= "000000";
					when "00011010100010101" => rgb <= "000000";
					when "00011010100010110" => rgb <= "000000";
					when "00011010100010111" => rgb <= "000000";
					when "00011010100011000" => rgb <= "000000";
					when "00011010100011001" => rgb <= "000000";
					when "00011010100011010" => rgb <= "000000";
					when "00011010100011011" => rgb <= "000000";
					when "00011010100011100" => rgb <= "000000";
					when "00011010100011101" => rgb <= "000000";
					when "00011010100011110" => rgb <= "000000";
					when "00011010100011111" => rgb <= "000000";
					when "00011010100100000" => rgb <= "000000";
					when "00011010100100001" => rgb <= "000000";
					when "00011010100100010" => rgb <= "000000";
					when "00011010100100011" => rgb <= "000000";
					when "00011010100100100" => rgb <= "000000";
					when "00011010100100101" => rgb <= "000000";
					when "00011010100100110" => rgb <= "000000";
					when "00011010100100111" => rgb <= "000000";
					when "00011010100101000" => rgb <= "000000";
					when "00011010100101001" => rgb <= "000000";
					when "00011010100101010" => rgb <= "000000";
					when "00011010100101011" => rgb <= "000000";
					when "00011010100101100" => rgb <= "000000";
					when "00011010100101101" => rgb <= "000000";
					when "00011010100101110" => rgb <= "000000";
					when "00011010100101111" => rgb <= "000000";
					when "00011010100110000" => rgb <= "000000";
					when "00011010100110001" => rgb <= "000000";
					when "00011010100110010" => rgb <= "000000";
					when "00011010100110011" => rgb <= "000000";
					when "00011010100110100" => rgb <= "000000";
					when "00011010100110101" => rgb <= "000000";
					when "00011010100110110" => rgb <= "000000";
					when "00011010100110111" => rgb <= "000000";
					when "00011010100111000" => rgb <= "000000";
					when "00011010100111001" => rgb <= "000000";
					when "00011010100111010" => rgb <= "000000";
					when "00011010100111011" => rgb <= "000000";
					when "00011010100111100" => rgb <= "000000";
					when "00011010100111101" => rgb <= "000000";
					when "00011010100111110" => rgb <= "000000";
					when "00011010100111111" => rgb <= "000000";
					when "00011011000000000" => rgb <= "000000";
					when "00011011000000001" => rgb <= "000000";
					when "00011011000000010" => rgb <= "000000";
					when "00011011000000011" => rgb <= "000000";
					when "00011011000000100" => rgb <= "000000";
					when "00011011000000101" => rgb <= "000000";
					when "00011011000000110" => rgb <= "000000";
					when "00011011000000111" => rgb <= "000000";
					when "00011011000001000" => rgb <= "000000";
					when "00011011000001001" => rgb <= "000000";
					when "00011011000001010" => rgb <= "000000";
					when "00011011000001011" => rgb <= "000000";
					when "00011011000001100" => rgb <= "000000";
					when "00011011000001101" => rgb <= "000000";
					when "00011011000001110" => rgb <= "000000";
					when "00011011000001111" => rgb <= "000000";
					when "00011011000010000" => rgb <= "000000";
					when "00011011000010001" => rgb <= "000000";
					when "00011011000010010" => rgb <= "000000";
					when "00011011000010011" => rgb <= "000000";
					when "00011011000010100" => rgb <= "000000";
					when "00011011000010101" => rgb <= "000000";
					when "00011011000010110" => rgb <= "000000";
					when "00011011000010111" => rgb <= "000000";
					when "00011011000011000" => rgb <= "000000";
					when "00011011000011001" => rgb <= "000000";
					when "00011011000011010" => rgb <= "000000";
					when "00011011000011011" => rgb <= "000000";
					when "00011011000011100" => rgb <= "000000";
					when "00011011000011101" => rgb <= "000000";
					when "00011011000011110" => rgb <= "000000";
					when "00011011000011111" => rgb <= "000000";
					when "00011011000100000" => rgb <= "000000";
					when "00011011000100001" => rgb <= "000000";
					when "00011011000100010" => rgb <= "000000";
					when "00011011000100011" => rgb <= "000000";
					when "00011011000100100" => rgb <= "000000";
					when "00011011000100101" => rgb <= "000000";
					when "00011011000100110" => rgb <= "000000";
					when "00011011000100111" => rgb <= "000000";
					when "00011011000101000" => rgb <= "000000";
					when "00011011000101001" => rgb <= "000000";
					when "00011011000101010" => rgb <= "000000";
					when "00011011000101011" => rgb <= "000000";
					when "00011011000101100" => rgb <= "000000";
					when "00011011000101101" => rgb <= "000000";
					when "00011011000101110" => rgb <= "000000";
					when "00011011000101111" => rgb <= "000000";
					when "00011011000110000" => rgb <= "000000";
					when "00011011000110001" => rgb <= "000000";
					when "00011011000110010" => rgb <= "000000";
					when "00011011000110011" => rgb <= "000000";
					when "00011011000110100" => rgb <= "000000";
					when "00011011000110101" => rgb <= "000000";
					when "00011011000110110" => rgb <= "000000";
					when "00011011000110111" => rgb <= "000000";
					when "00011011000111000" => rgb <= "000000";
					when "00011011000111001" => rgb <= "000000";
					when "00011011000111010" => rgb <= "000000";
					when "00011011000111011" => rgb <= "000000";
					when "00011011000111100" => rgb <= "000000";
					when "00011011000111101" => rgb <= "000000";
					when "00011011000111110" => rgb <= "000000";
					when "00011011000111111" => rgb <= "000000";
					when "00011011001000000" => rgb <= "000000";
					when "00011011001000001" => rgb <= "000000";
					when "00011011001000010" => rgb <= "000000";
					when "00011011001000011" => rgb <= "000000";
					when "00011011001000100" => rgb <= "000000";
					when "00011011001000101" => rgb <= "000000";
					when "00011011001000110" => rgb <= "000000";
					when "00011011001000111" => rgb <= "000000";
					when "00011011001001000" => rgb <= "000000";
					when "00011011001001001" => rgb <= "000000";
					when "00011011001001010" => rgb <= "000000";
					when "00011011001001011" => rgb <= "000000";
					when "00011011001001100" => rgb <= "000000";
					when "00011011001001101" => rgb <= "000000";
					when "00011011001001110" => rgb <= "000000";
					when "00011011001001111" => rgb <= "000000";
					when "00011011001010000" => rgb <= "000000";
					when "00011011001010001" => rgb <= "000000";
					when "00011011001010010" => rgb <= "000000";
					when "00011011001010011" => rgb <= "000000";
					when "00011011001010100" => rgb <= "000000";
					when "00011011001010101" => rgb <= "000000";
					when "00011011001010110" => rgb <= "000000";
					when "00011011001010111" => rgb <= "000000";
					when "00011011001011000" => rgb <= "000000";
					when "00011011001011001" => rgb <= "000000";
					when "00011011001011010" => rgb <= "000000";
					when "00011011001011011" => rgb <= "000000";
					when "00011011001011100" => rgb <= "000000";
					when "00011011001011101" => rgb <= "000000";
					when "00011011001011110" => rgb <= "000000";
					when "00011011001011111" => rgb <= "000000";
					when "00011011001100000" => rgb <= "000000";
					when "00011011001100001" => rgb <= "000000";
					when "00011011001100010" => rgb <= "000000";
					when "00011011001100011" => rgb <= "000000";
					when "00011011001100100" => rgb <= "000000";
					when "00011011001100101" => rgb <= "000000";
					when "00011011001100110" => rgb <= "000000";
					when "00011011001100111" => rgb <= "000000";
					when "00011011001101000" => rgb <= "000000";
					when "00011011001101001" => rgb <= "000000";
					when "00011011001101010" => rgb <= "000000";
					when "00011011001101011" => rgb <= "000000";
					when "00011011001101100" => rgb <= "000000";
					when "00011011001101101" => rgb <= "000000";
					when "00011011001101110" => rgb <= "000000";
					when "00011011001101111" => rgb <= "000000";
					when "00011011001110000" => rgb <= "000000";
					when "00011011001110001" => rgb <= "000000";
					when "00011011001110010" => rgb <= "000000";
					when "00011011001110011" => rgb <= "000000";
					when "00011011001110100" => rgb <= "000000";
					when "00011011001110101" => rgb <= "000000";
					when "00011011001110110" => rgb <= "000000";
					when "00011011001110111" => rgb <= "000000";
					when "00011011001111000" => rgb <= "000000";
					when "00011011001111001" => rgb <= "000000";
					when "00011011001111010" => rgb <= "000000";
					when "00011011001111011" => rgb <= "000000";
					when "00011011001111100" => rgb <= "000000";
					when "00011011001111101" => rgb <= "101000";
					when "00011011001111110" => rgb <= "101000";
					when "00011011001111111" => rgb <= "101000";
					when "00011011010000000" => rgb <= "101000";
					when "00011011010000001" => rgb <= "101000";
					when "00011011010000010" => rgb <= "101000";
					when "00011011010000011" => rgb <= "101000";
					when "00011011010000100" => rgb <= "101000";
					when "00011011010000101" => rgb <= "101000";
					when "00011011010000110" => rgb <= "101000";
					when "00011011010000111" => rgb <= "101000";
					when "00011011010001000" => rgb <= "101000";
					when "00011011010001001" => rgb <= "101000";
					when "00011011010001010" => rgb <= "101000";
					when "00011011010001011" => rgb <= "101000";
					when "00011011010001100" => rgb <= "101000";
					when "00011011010001101" => rgb <= "101000";
					when "00011011010001110" => rgb <= "101000";
					when "00011011010001111" => rgb <= "101000";
					when "00011011010010000" => rgb <= "101000";
					when "00011011010010001" => rgb <= "101000";
					when "00011011010010010" => rgb <= "101000";
					when "00011011010010011" => rgb <= "101000";
					when "00011011010010100" => rgb <= "101000";
					when "00011011010010101" => rgb <= "101000";
					when "00011011010010110" => rgb <= "101000";
					when "00011011010010111" => rgb <= "101000";
					when "00011011010011000" => rgb <= "101000";
					when "00011011010011001" => rgb <= "101000";
					when "00011011010011010" => rgb <= "101000";
					when "00011011010011011" => rgb <= "101000";
					when "00011011010011100" => rgb <= "101000";
					when "00011011010011101" => rgb <= "101000";
					when "00011011010011110" => rgb <= "101000";
					when "00011011010011111" => rgb <= "101000";
					when "00011011010100000" => rgb <= "101000";
					when "00011011010100001" => rgb <= "101000";
					when "00011011010100010" => rgb <= "101000";
					when "00011011010100011" => rgb <= "101000";
					when "00011011010100100" => rgb <= "101000";
					when "00011011010100101" => rgb <= "101000";
					when "00011011010100110" => rgb <= "101000";
					when "00011011010100111" => rgb <= "101000";
					when "00011011010101000" => rgb <= "101000";
					when "00011011010101001" => rgb <= "101000";
					when "00011011010101010" => rgb <= "101000";
					when "00011011010101011" => rgb <= "101000";
					when "00011011010101100" => rgb <= "101000";
					when "00011011010101101" => rgb <= "101000";
					when "00011011010101110" => rgb <= "101000";
					when "00011011010101111" => rgb <= "101000";
					when "00011011010110000" => rgb <= "101000";
					when "00011011010110001" => rgb <= "101000";
					when "00011011010110010" => rgb <= "101000";
					when "00011011010110011" => rgb <= "101000";
					when "00011011010110100" => rgb <= "101000";
					when "00011011010110101" => rgb <= "101000";
					when "00011011010110110" => rgb <= "101000";
					when "00011011010110111" => rgb <= "101000";
					when "00011011010111000" => rgb <= "101000";
					when "00011011010111001" => rgb <= "101000";
					when "00011011010111010" => rgb <= "101000";
					when "00011011010111011" => rgb <= "101000";
					when "00011011010111100" => rgb <= "101000";
					when "00011011010111101" => rgb <= "101000";
					when "00011011010111110" => rgb <= "101000";
					when "00011011010111111" => rgb <= "101000";
					when "00011011011000000" => rgb <= "100100";
					when "00011011011000001" => rgb <= "000000";
					when "00011011011000010" => rgb <= "000000";
					when "00011011011000011" => rgb <= "000000";
					when "00011011011000100" => rgb <= "000000";
					when "00011011011000101" => rgb <= "000000";
					when "00011011011000110" => rgb <= "000000";
					when "00011011011000111" => rgb <= "000000";
					when "00011011011001000" => rgb <= "000000";
					when "00011011011001001" => rgb <= "000000";
					when "00011011011001010" => rgb <= "000000";
					when "00011011011001011" => rgb <= "000000";
					when "00011011011001100" => rgb <= "000000";
					when "00011011011001101" => rgb <= "000000";
					when "00011011011001110" => rgb <= "000000";
					when "00011011011001111" => rgb <= "000000";
					when "00011011011010000" => rgb <= "000000";
					when "00011011011010001" => rgb <= "000000";
					when "00011011011010010" => rgb <= "000000";
					when "00011011011010011" => rgb <= "000000";
					when "00011011011010100" => rgb <= "000000";
					when "00011011011010101" => rgb <= "000000";
					when "00011011011010110" => rgb <= "000000";
					when "00011011011010111" => rgb <= "000000";
					when "00011011011011000" => rgb <= "000000";
					when "00011011011011001" => rgb <= "000000";
					when "00011011011011010" => rgb <= "000000";
					when "00011011011011011" => rgb <= "000000";
					when "00011011011011100" => rgb <= "000000";
					when "00011011011011101" => rgb <= "000000";
					when "00011011011011110" => rgb <= "000000";
					when "00011011011011111" => rgb <= "000000";
					when "00011011011100000" => rgb <= "000000";
					when "00011011011100001" => rgb <= "000000";
					when "00011011011100010" => rgb <= "000000";
					when "00011011011100011" => rgb <= "000000";
					when "00011011011100100" => rgb <= "000000";
					when "00011011011100101" => rgb <= "000000";
					when "00011011011100110" => rgb <= "000000";
					when "00011011011100111" => rgb <= "000000";
					when "00011011011101000" => rgb <= "000000";
					when "00011011011101001" => rgb <= "000000";
					when "00011011011101010" => rgb <= "000000";
					when "00011011011101011" => rgb <= "000000";
					when "00011011011101100" => rgb <= "000000";
					when "00011011011101101" => rgb <= "000000";
					when "00011011011101110" => rgb <= "000000";
					when "00011011011101111" => rgb <= "000000";
					when "00011011011110000" => rgb <= "000000";
					when "00011011011110001" => rgb <= "000000";
					when "00011011011110010" => rgb <= "000000";
					when "00011011011110011" => rgb <= "000000";
					when "00011011011110100" => rgb <= "000000";
					when "00011011011110101" => rgb <= "000000";
					when "00011011011110110" => rgb <= "000000";
					when "00011011011110111" => rgb <= "000000";
					when "00011011011111000" => rgb <= "000000";
					when "00011011011111001" => rgb <= "000000";
					when "00011011011111010" => rgb <= "000000";
					when "00011011011111011" => rgb <= "000000";
					when "00011011011111100" => rgb <= "000000";
					when "00011011011111101" => rgb <= "000000";
					when "00011011011111110" => rgb <= "000000";
					when "00011011011111111" => rgb <= "000000";
					when "00011011100000000" => rgb <= "000000";
					when "00011011100000001" => rgb <= "000000";
					when "00011011100000010" => rgb <= "000000";
					when "00011011100000011" => rgb <= "000000";
					when "00011011100000100" => rgb <= "000000";
					when "00011011100000101" => rgb <= "000000";
					when "00011011100000110" => rgb <= "000000";
					when "00011011100000111" => rgb <= "000000";
					when "00011011100001000" => rgb <= "000000";
					when "00011011100001001" => rgb <= "000000";
					when "00011011100001010" => rgb <= "000000";
					when "00011011100001011" => rgb <= "000000";
					when "00011011100001100" => rgb <= "000000";
					when "00011011100001101" => rgb <= "000000";
					when "00011011100001110" => rgb <= "000000";
					when "00011011100001111" => rgb <= "000000";
					when "00011011100010000" => rgb <= "000000";
					when "00011011100010001" => rgb <= "000000";
					when "00011011100010010" => rgb <= "000000";
					when "00011011100010011" => rgb <= "000000";
					when "00011011100010100" => rgb <= "000000";
					when "00011011100010101" => rgb <= "000000";
					when "00011011100010110" => rgb <= "000000";
					when "00011011100010111" => rgb <= "000000";
					when "00011011100011000" => rgb <= "000000";
					when "00011011100011001" => rgb <= "000000";
					when "00011011100011010" => rgb <= "000000";
					when "00011011100011011" => rgb <= "000000";
					when "00011011100011100" => rgb <= "000000";
					when "00011011100011101" => rgb <= "000000";
					when "00011011100011110" => rgb <= "000000";
					when "00011011100011111" => rgb <= "000000";
					when "00011011100100000" => rgb <= "000000";
					when "00011011100100001" => rgb <= "000000";
					when "00011011100100010" => rgb <= "000000";
					when "00011011100100011" => rgb <= "000000";
					when "00011011100100100" => rgb <= "000000";
					when "00011011100100101" => rgb <= "000000";
					when "00011011100100110" => rgb <= "000000";
					when "00011011100100111" => rgb <= "000000";
					when "00011011100101000" => rgb <= "000000";
					when "00011011100101001" => rgb <= "000000";
					when "00011011100101010" => rgb <= "000000";
					when "00011011100101011" => rgb <= "000000";
					when "00011011100101100" => rgb <= "000000";
					when "00011011100101101" => rgb <= "000000";
					when "00011011100101110" => rgb <= "000000";
					when "00011011100101111" => rgb <= "000000";
					when "00011011100110000" => rgb <= "000000";
					when "00011011100110001" => rgb <= "000000";
					when "00011011100110010" => rgb <= "000000";
					when "00011011100110011" => rgb <= "000000";
					when "00011011100110100" => rgb <= "000000";
					when "00011011100110101" => rgb <= "000000";
					when "00011011100110110" => rgb <= "000000";
					when "00011011100110111" => rgb <= "000000";
					when "00011011100111000" => rgb <= "000000";
					when "00011011100111001" => rgb <= "000000";
					when "00011011100111010" => rgb <= "000000";
					when "00011011100111011" => rgb <= "000000";
					when "00011011100111100" => rgb <= "000000";
					when "00011011100111101" => rgb <= "000000";
					when "00011011100111110" => rgb <= "000000";
					when "00011011100111111" => rgb <= "000000";
					when "00011100000000000" => rgb <= "000000";
					when "00011100000000001" => rgb <= "000000";
					when "00011100000000010" => rgb <= "000000";
					when "00011100000000011" => rgb <= "000000";
					when "00011100000000100" => rgb <= "000000";
					when "00011100000000101" => rgb <= "000000";
					when "00011100000000110" => rgb <= "000000";
					when "00011100000000111" => rgb <= "000000";
					when "00011100000001000" => rgb <= "000000";
					when "00011100000001001" => rgb <= "000000";
					when "00011100000001010" => rgb <= "000000";
					when "00011100000001011" => rgb <= "000000";
					when "00011100000001100" => rgb <= "000000";
					when "00011100000001101" => rgb <= "000000";
					when "00011100000001110" => rgb <= "000000";
					when "00011100000001111" => rgb <= "000000";
					when "00011100000010000" => rgb <= "000000";
					when "00011100000010001" => rgb <= "000000";
					when "00011100000010010" => rgb <= "000000";
					when "00011100000010011" => rgb <= "000000";
					when "00011100000010100" => rgb <= "000000";
					when "00011100000010101" => rgb <= "000000";
					when "00011100000010110" => rgb <= "000000";
					when "00011100000010111" => rgb <= "000000";
					when "00011100000011000" => rgb <= "000000";
					when "00011100000011001" => rgb <= "000000";
					when "00011100000011010" => rgb <= "000000";
					when "00011100000011011" => rgb <= "000000";
					when "00011100000011100" => rgb <= "000000";
					when "00011100000011101" => rgb <= "000000";
					when "00011100000011110" => rgb <= "000000";
					when "00011100000011111" => rgb <= "000000";
					when "00011100000100000" => rgb <= "000000";
					when "00011100000100001" => rgb <= "000000";
					when "00011100000100010" => rgb <= "000000";
					when "00011100000100011" => rgb <= "000000";
					when "00011100000100100" => rgb <= "000000";
					when "00011100000100101" => rgb <= "000000";
					when "00011100000100110" => rgb <= "000000";
					when "00011100000100111" => rgb <= "000000";
					when "00011100000101000" => rgb <= "000000";
					when "00011100000101001" => rgb <= "000000";
					when "00011100000101010" => rgb <= "000000";
					when "00011100000101011" => rgb <= "000000";
					when "00011100000101100" => rgb <= "000000";
					when "00011100000101101" => rgb <= "000000";
					when "00011100000101110" => rgb <= "000000";
					when "00011100000101111" => rgb <= "000000";
					when "00011100000110000" => rgb <= "000000";
					when "00011100000110001" => rgb <= "000000";
					when "00011100000110010" => rgb <= "000000";
					when "00011100000110011" => rgb <= "000000";
					when "00011100000110100" => rgb <= "000000";
					when "00011100000110101" => rgb <= "000000";
					when "00011100000110110" => rgb <= "000000";
					when "00011100000110111" => rgb <= "000000";
					when "00011100000111000" => rgb <= "000000";
					when "00011100000111001" => rgb <= "000000";
					when "00011100000111010" => rgb <= "000000";
					when "00011100000111011" => rgb <= "000000";
					when "00011100000111100" => rgb <= "000000";
					when "00011100000111101" => rgb <= "000000";
					when "00011100000111110" => rgb <= "000000";
					when "00011100000111111" => rgb <= "000000";
					when "00011100001000000" => rgb <= "000000";
					when "00011100001000001" => rgb <= "000000";
					when "00011100001000010" => rgb <= "000000";
					when "00011100001000011" => rgb <= "000000";
					when "00011100001000100" => rgb <= "000000";
					when "00011100001000101" => rgb <= "000000";
					when "00011100001000110" => rgb <= "000000";
					when "00011100001000111" => rgb <= "000000";
					when "00011100001001000" => rgb <= "000000";
					when "00011100001001001" => rgb <= "000000";
					when "00011100001001010" => rgb <= "000000";
					when "00011100001001011" => rgb <= "000000";
					when "00011100001001100" => rgb <= "000000";
					when "00011100001001101" => rgb <= "000000";
					when "00011100001001110" => rgb <= "000000";
					when "00011100001001111" => rgb <= "000000";
					when "00011100001010000" => rgb <= "000000";
					when "00011100001010001" => rgb <= "000000";
					when "00011100001010010" => rgb <= "000000";
					when "00011100001010011" => rgb <= "000000";
					when "00011100001010100" => rgb <= "000000";
					when "00011100001010101" => rgb <= "000000";
					when "00011100001010110" => rgb <= "000000";
					when "00011100001010111" => rgb <= "000000";
					when "00011100001011000" => rgb <= "000000";
					when "00011100001011001" => rgb <= "000000";
					when "00011100001011010" => rgb <= "000000";
					when "00011100001011011" => rgb <= "000000";
					when "00011100001011100" => rgb <= "000000";
					when "00011100001011101" => rgb <= "000000";
					when "00011100001011110" => rgb <= "000000";
					when "00011100001011111" => rgb <= "000000";
					when "00011100001100000" => rgb <= "000000";
					when "00011100001100001" => rgb <= "000000";
					when "00011100001100010" => rgb <= "000000";
					when "00011100001100011" => rgb <= "000000";
					when "00011100001100100" => rgb <= "000000";
					when "00011100001100101" => rgb <= "000000";
					when "00011100001100110" => rgb <= "000000";
					when "00011100001100111" => rgb <= "000000";
					when "00011100001101000" => rgb <= "000000";
					when "00011100001101001" => rgb <= "000000";
					when "00011100001101010" => rgb <= "000000";
					when "00011100001101011" => rgb <= "000000";
					when "00011100001101100" => rgb <= "000000";
					when "00011100001101101" => rgb <= "000000";
					when "00011100001101110" => rgb <= "000000";
					when "00011100001101111" => rgb <= "000000";
					when "00011100001110000" => rgb <= "000000";
					when "00011100001110001" => rgb <= "000000";
					when "00011100001110010" => rgb <= "000000";
					when "00011100001110011" => rgb <= "000000";
					when "00011100001110100" => rgb <= "000000";
					when "00011100001110101" => rgb <= "000000";
					when "00011100001110110" => rgb <= "000000";
					when "00011100001110111" => rgb <= "000000";
					when "00011100001111000" => rgb <= "000000";
					when "00011100001111001" => rgb <= "000000";
					when "00011100001111010" => rgb <= "000000";
					when "00011100001111011" => rgb <= "000000";
					when "00011100001111100" => rgb <= "000000";
					when "00011100001111101" => rgb <= "101000";
					when "00011100001111110" => rgb <= "101000";
					when "00011100001111111" => rgb <= "101000";
					when "00011100010000000" => rgb <= "101000";
					when "00011100010000001" => rgb <= "101000";
					when "00011100010000010" => rgb <= "101000";
					when "00011100010000011" => rgb <= "101000";
					when "00011100010000100" => rgb <= "101000";
					when "00011100010000101" => rgb <= "101000";
					when "00011100010000110" => rgb <= "101000";
					when "00011100010000111" => rgb <= "101000";
					when "00011100010001000" => rgb <= "101001";
					when "00011100010001001" => rgb <= "101001";
					when "00011100010001010" => rgb <= "101001";
					when "00011100010001011" => rgb <= "101001";
					when "00011100010001100" => rgb <= "101001";
					when "00011100010001101" => rgb <= "101001";
					when "00011100010001110" => rgb <= "101001";
					when "00011100010001111" => rgb <= "101001";
					when "00011100010010000" => rgb <= "101001";
					when "00011100010010001" => rgb <= "101001";
					when "00011100010010010" => rgb <= "101001";
					when "00011100010010011" => rgb <= "101001";
					when "00011100010010100" => rgb <= "101001";
					when "00011100010010101" => rgb <= "101001";
					when "00011100010010110" => rgb <= "101001";
					when "00011100010010111" => rgb <= "101001";
					when "00011100010011000" => rgb <= "101001";
					when "00011100010011001" => rgb <= "101001";
					when "00011100010011010" => rgb <= "101001";
					when "00011100010011011" => rgb <= "101001";
					when "00011100010011100" => rgb <= "101001";
					when "00011100010011101" => rgb <= "101001";
					when "00011100010011110" => rgb <= "101001";
					when "00011100010011111" => rgb <= "101000";
					when "00011100010100000" => rgb <= "101000";
					when "00011100010100001" => rgb <= "101000";
					when "00011100010100010" => rgb <= "101000";
					when "00011100010100011" => rgb <= "101000";
					when "00011100010100100" => rgb <= "101000";
					when "00011100010100101" => rgb <= "101000";
					when "00011100010100110" => rgb <= "101000";
					when "00011100010100111" => rgb <= "101000";
					when "00011100010101000" => rgb <= "101000";
					when "00011100010101001" => rgb <= "101000";
					when "00011100010101010" => rgb <= "101000";
					when "00011100010101011" => rgb <= "101000";
					when "00011100010101100" => rgb <= "101000";
					when "00011100010101101" => rgb <= "101000";
					when "00011100010101110" => rgb <= "101000";
					when "00011100010101111" => rgb <= "101000";
					when "00011100010110000" => rgb <= "101000";
					when "00011100010110001" => rgb <= "101000";
					when "00011100010110010" => rgb <= "101000";
					when "00011100010110011" => rgb <= "101000";
					when "00011100010110100" => rgb <= "101000";
					when "00011100010110101" => rgb <= "101000";
					when "00011100010110110" => rgb <= "101000";
					when "00011100010110111" => rgb <= "101000";
					when "00011100010111000" => rgb <= "101000";
					when "00011100010111001" => rgb <= "101000";
					when "00011100010111010" => rgb <= "101000";
					when "00011100010111011" => rgb <= "101000";
					when "00011100010111100" => rgb <= "101000";
					when "00011100010111101" => rgb <= "101000";
					when "00011100010111110" => rgb <= "101000";
					when "00011100010111111" => rgb <= "101000";
					when "00011100011000000" => rgb <= "100100";
					when "00011100011000001" => rgb <= "000000";
					when "00011100011000010" => rgb <= "000000";
					when "00011100011000011" => rgb <= "000000";
					when "00011100011000100" => rgb <= "000000";
					when "00011100011000101" => rgb <= "000000";
					when "00011100011000110" => rgb <= "000000";
					when "00011100011000111" => rgb <= "000000";
					when "00011100011001000" => rgb <= "000000";
					when "00011100011001001" => rgb <= "000000";
					when "00011100011001010" => rgb <= "000000";
					when "00011100011001011" => rgb <= "000000";
					when "00011100011001100" => rgb <= "000000";
					when "00011100011001101" => rgb <= "000000";
					when "00011100011001110" => rgb <= "000000";
					when "00011100011001111" => rgb <= "000000";
					when "00011100011010000" => rgb <= "000000";
					when "00011100011010001" => rgb <= "000000";
					when "00011100011010010" => rgb <= "000000";
					when "00011100011010011" => rgb <= "000000";
					when "00011100011010100" => rgb <= "000000";
					when "00011100011010101" => rgb <= "000000";
					when "00011100011010110" => rgb <= "000000";
					when "00011100011010111" => rgb <= "000000";
					when "00011100011011000" => rgb <= "000000";
					when "00011100011011001" => rgb <= "000000";
					when "00011100011011010" => rgb <= "000000";
					when "00011100011011011" => rgb <= "000000";
					when "00011100011011100" => rgb <= "000000";
					when "00011100011011101" => rgb <= "000000";
					when "00011100011011110" => rgb <= "000000";
					when "00011100011011111" => rgb <= "000000";
					when "00011100011100000" => rgb <= "000000";
					when "00011100011100001" => rgb <= "000000";
					when "00011100011100010" => rgb <= "000000";
					when "00011100011100011" => rgb <= "000000";
					when "00011100011100100" => rgb <= "000000";
					when "00011100011100101" => rgb <= "000000";
					when "00011100011100110" => rgb <= "000000";
					when "00011100011100111" => rgb <= "000000";
					when "00011100011101000" => rgb <= "000000";
					when "00011100011101001" => rgb <= "000000";
					when "00011100011101010" => rgb <= "000000";
					when "00011100011101011" => rgb <= "000000";
					when "00011100011101100" => rgb <= "000000";
					when "00011100011101101" => rgb <= "000000";
					when "00011100011101110" => rgb <= "000000";
					when "00011100011101111" => rgb <= "000000";
					when "00011100011110000" => rgb <= "000000";
					when "00011100011110001" => rgb <= "000000";
					when "00011100011110010" => rgb <= "000000";
					when "00011100011110011" => rgb <= "000000";
					when "00011100011110100" => rgb <= "000000";
					when "00011100011110101" => rgb <= "000000";
					when "00011100011110110" => rgb <= "000000";
					when "00011100011110111" => rgb <= "000000";
					when "00011100011111000" => rgb <= "000000";
					when "00011100011111001" => rgb <= "000000";
					when "00011100011111010" => rgb <= "000000";
					when "00011100011111011" => rgb <= "000000";
					when "00011100011111100" => rgb <= "000000";
					when "00011100011111101" => rgb <= "000000";
					when "00011100011111110" => rgb <= "000000";
					when "00011100011111111" => rgb <= "000000";
					when "00011100100000000" => rgb <= "000000";
					when "00011100100000001" => rgb <= "000000";
					when "00011100100000010" => rgb <= "000000";
					when "00011100100000011" => rgb <= "000000";
					when "00011100100000100" => rgb <= "000000";
					when "00011100100000101" => rgb <= "000000";
					when "00011100100000110" => rgb <= "000000";
					when "00011100100000111" => rgb <= "000000";
					when "00011100100001000" => rgb <= "000000";
					when "00011100100001001" => rgb <= "000000";
					when "00011100100001010" => rgb <= "000000";
					when "00011100100001011" => rgb <= "000000";
					when "00011100100001100" => rgb <= "000000";
					when "00011100100001101" => rgb <= "000000";
					when "00011100100001110" => rgb <= "000000";
					when "00011100100001111" => rgb <= "000000";
					when "00011100100010000" => rgb <= "000000";
					when "00011100100010001" => rgb <= "000000";
					when "00011100100010010" => rgb <= "000000";
					when "00011100100010011" => rgb <= "000000";
					when "00011100100010100" => rgb <= "000000";
					when "00011100100010101" => rgb <= "000000";
					when "00011100100010110" => rgb <= "000000";
					when "00011100100010111" => rgb <= "000000";
					when "00011100100011000" => rgb <= "000000";
					when "00011100100011001" => rgb <= "000000";
					when "00011100100011010" => rgb <= "000000";
					when "00011100100011011" => rgb <= "000000";
					when "00011100100011100" => rgb <= "000000";
					when "00011100100011101" => rgb <= "000000";
					when "00011100100011110" => rgb <= "000000";
					when "00011100100011111" => rgb <= "000000";
					when "00011100100100000" => rgb <= "000000";
					when "00011100100100001" => rgb <= "000000";
					when "00011100100100010" => rgb <= "000000";
					when "00011100100100011" => rgb <= "000000";
					when "00011100100100100" => rgb <= "000000";
					when "00011100100100101" => rgb <= "000000";
					when "00011100100100110" => rgb <= "000000";
					when "00011100100100111" => rgb <= "000000";
					when "00011100100101000" => rgb <= "000000";
					when "00011100100101001" => rgb <= "000000";
					when "00011100100101010" => rgb <= "000000";
					when "00011100100101011" => rgb <= "000000";
					when "00011100100101100" => rgb <= "000000";
					when "00011100100101101" => rgb <= "000000";
					when "00011100100101110" => rgb <= "000000";
					when "00011100100101111" => rgb <= "000000";
					when "00011100100110000" => rgb <= "000000";
					when "00011100100110001" => rgb <= "000000";
					when "00011100100110010" => rgb <= "000000";
					when "00011100100110011" => rgb <= "000000";
					when "00011100100110100" => rgb <= "000000";
					when "00011100100110101" => rgb <= "000000";
					when "00011100100110110" => rgb <= "000000";
					when "00011100100110111" => rgb <= "000000";
					when "00011100100111000" => rgb <= "000000";
					when "00011100100111001" => rgb <= "000000";
					when "00011100100111010" => rgb <= "000000";
					when "00011100100111011" => rgb <= "000000";
					when "00011100100111100" => rgb <= "000000";
					when "00011100100111101" => rgb <= "000000";
					when "00011100100111110" => rgb <= "000000";
					when "00011100100111111" => rgb <= "000000";
					when "00011101000000000" => rgb <= "000000";
					when "00011101000000001" => rgb <= "000000";
					when "00011101000000010" => rgb <= "000000";
					when "00011101000000011" => rgb <= "000000";
					when "00011101000000100" => rgb <= "000000";
					when "00011101000000101" => rgb <= "000000";
					when "00011101000000110" => rgb <= "000000";
					when "00011101000000111" => rgb <= "000000";
					when "00011101000001000" => rgb <= "000000";
					when "00011101000001001" => rgb <= "000000";
					when "00011101000001010" => rgb <= "000000";
					when "00011101000001011" => rgb <= "000000";
					when "00011101000001100" => rgb <= "000000";
					when "00011101000001101" => rgb <= "000000";
					when "00011101000001110" => rgb <= "000000";
					when "00011101000001111" => rgb <= "000000";
					when "00011101000010000" => rgb <= "000000";
					when "00011101000010001" => rgb <= "000000";
					when "00011101000010010" => rgb <= "000000";
					when "00011101000010011" => rgb <= "000000";
					when "00011101000010100" => rgb <= "000000";
					when "00011101000010101" => rgb <= "000000";
					when "00011101000010110" => rgb <= "000000";
					when "00011101000010111" => rgb <= "000000";
					when "00011101000011000" => rgb <= "000000";
					when "00011101000011001" => rgb <= "000000";
					when "00011101000011010" => rgb <= "000000";
					when "00011101000011011" => rgb <= "000000";
					when "00011101000011100" => rgb <= "000000";
					when "00011101000011101" => rgb <= "000000";
					when "00011101000011110" => rgb <= "000000";
					when "00011101000011111" => rgb <= "000000";
					when "00011101000100000" => rgb <= "000000";
					when "00011101000100001" => rgb <= "000000";
					when "00011101000100010" => rgb <= "000000";
					when "00011101000100011" => rgb <= "000000";
					when "00011101000100100" => rgb <= "000000";
					when "00011101000100101" => rgb <= "000000";
					when "00011101000100110" => rgb <= "000000";
					when "00011101000100111" => rgb <= "000000";
					when "00011101000101000" => rgb <= "000000";
					when "00011101000101001" => rgb <= "000000";
					when "00011101000101010" => rgb <= "000000";
					when "00011101000101011" => rgb <= "000000";
					when "00011101000101100" => rgb <= "000000";
					when "00011101000101101" => rgb <= "000000";
					when "00011101000101110" => rgb <= "000000";
					when "00011101000101111" => rgb <= "000000";
					when "00011101000110000" => rgb <= "000000";
					when "00011101000110001" => rgb <= "000000";
					when "00011101000110010" => rgb <= "000000";
					when "00011101000110011" => rgb <= "000000";
					when "00011101000110100" => rgb <= "000000";
					when "00011101000110101" => rgb <= "000000";
					when "00011101000110110" => rgb <= "000000";
					when "00011101000110111" => rgb <= "000000";
					when "00011101000111000" => rgb <= "000000";
					when "00011101000111001" => rgb <= "000000";
					when "00011101000111010" => rgb <= "000000";
					when "00011101000111011" => rgb <= "000000";
					when "00011101000111100" => rgb <= "000000";
					when "00011101000111101" => rgb <= "000000";
					when "00011101000111110" => rgb <= "000000";
					when "00011101000111111" => rgb <= "000000";
					when "00011101001000000" => rgb <= "000000";
					when "00011101001000001" => rgb <= "000000";
					when "00011101001000010" => rgb <= "000000";
					when "00011101001000011" => rgb <= "000000";
					when "00011101001000100" => rgb <= "000000";
					when "00011101001000101" => rgb <= "000000";
					when "00011101001000110" => rgb <= "000000";
					when "00011101001000111" => rgb <= "000000";
					when "00011101001001000" => rgb <= "000000";
					when "00011101001001001" => rgb <= "000000";
					when "00011101001001010" => rgb <= "000000";
					when "00011101001001011" => rgb <= "000000";
					when "00011101001001100" => rgb <= "000000";
					when "00011101001001101" => rgb <= "000000";
					when "00011101001001110" => rgb <= "000000";
					when "00011101001001111" => rgb <= "000000";
					when "00011101001010000" => rgb <= "000000";
					when "00011101001010001" => rgb <= "000000";
					when "00011101001010010" => rgb <= "000000";
					when "00011101001010011" => rgb <= "000000";
					when "00011101001010100" => rgb <= "000000";
					when "00011101001010101" => rgb <= "000000";
					when "00011101001010110" => rgb <= "000000";
					when "00011101001010111" => rgb <= "000000";
					when "00011101001011000" => rgb <= "000000";
					when "00011101001011001" => rgb <= "000000";
					when "00011101001011010" => rgb <= "000000";
					when "00011101001011011" => rgb <= "000000";
					when "00011101001011100" => rgb <= "000000";
					when "00011101001011101" => rgb <= "000000";
					when "00011101001011110" => rgb <= "000000";
					when "00011101001011111" => rgb <= "000000";
					when "00011101001100000" => rgb <= "000000";
					when "00011101001100001" => rgb <= "000000";
					when "00011101001100010" => rgb <= "000000";
					when "00011101001100011" => rgb <= "000000";
					when "00011101001100100" => rgb <= "000000";
					when "00011101001100101" => rgb <= "000000";
					when "00011101001100110" => rgb <= "000000";
					when "00011101001100111" => rgb <= "000000";
					when "00011101001101000" => rgb <= "000000";
					when "00011101001101001" => rgb <= "000000";
					when "00011101001101010" => rgb <= "000000";
					when "00011101001101011" => rgb <= "000000";
					when "00011101001101100" => rgb <= "000000";
					when "00011101001101101" => rgb <= "000000";
					when "00011101001101110" => rgb <= "000000";
					when "00011101001101111" => rgb <= "000000";
					when "00011101001110000" => rgb <= "000000";
					when "00011101001110001" => rgb <= "000000";
					when "00011101001110010" => rgb <= "000000";
					when "00011101001110011" => rgb <= "000000";
					when "00011101001110100" => rgb <= "000000";
					when "00011101001110101" => rgb <= "000000";
					when "00011101001110110" => rgb <= "000000";
					when "00011101001110111" => rgb <= "000000";
					when "00011101001111000" => rgb <= "000000";
					when "00011101001111001" => rgb <= "000000";
					when "00011101001111010" => rgb <= "000000";
					when "00011101001111011" => rgb <= "000000";
					when "00011101001111100" => rgb <= "000000";
					when "00011101001111101" => rgb <= "101000";
					when "00011101001111110" => rgb <= "101000";
					when "00011101001111111" => rgb <= "101000";
					when "00011101010000000" => rgb <= "101000";
					when "00011101010000001" => rgb <= "101000";
					when "00011101010000010" => rgb <= "101000";
					when "00011101010000011" => rgb <= "101000";
					when "00011101010000100" => rgb <= "101000";
					when "00011101010000101" => rgb <= "101000";
					when "00011101010000110" => rgb <= "101000";
					when "00011101010000111" => rgb <= "101000";
					when "00011101010001000" => rgb <= "101001";
					when "00011101010001001" => rgb <= "111001";
					when "00011101010001010" => rgb <= "111001";
					when "00011101010001011" => rgb <= "111001";
					when "00011101010001100" => rgb <= "111001";
					when "00011101010001101" => rgb <= "111001";
					when "00011101010001110" => rgb <= "111001";
					when "00011101010001111" => rgb <= "111001";
					when "00011101010010000" => rgb <= "111001";
					when "00011101010010001" => rgb <= "111001";
					when "00011101010010010" => rgb <= "111001";
					when "00011101010010011" => rgb <= "111001";
					when "00011101010010100" => rgb <= "111001";
					when "00011101010010101" => rgb <= "111001";
					when "00011101010010110" => rgb <= "111001";
					when "00011101010010111" => rgb <= "111001";
					when "00011101010011000" => rgb <= "111001";
					when "00011101010011001" => rgb <= "111001";
					when "00011101010011010" => rgb <= "111001";
					when "00011101010011011" => rgb <= "111001";
					when "00011101010011100" => rgb <= "111001";
					when "00011101010011101" => rgb <= "111010";
					when "00011101010011110" => rgb <= "111001";
					when "00011101010011111" => rgb <= "101001";
					when "00011101010100000" => rgb <= "101000";
					when "00011101010100001" => rgb <= "101000";
					when "00011101010100010" => rgb <= "101000";
					when "00011101010100011" => rgb <= "101000";
					when "00011101010100100" => rgb <= "101000";
					when "00011101010100101" => rgb <= "101000";
					when "00011101010100110" => rgb <= "101000";
					when "00011101010100111" => rgb <= "101000";
					when "00011101010101000" => rgb <= "101000";
					when "00011101010101001" => rgb <= "101000";
					when "00011101010101010" => rgb <= "101000";
					when "00011101010101011" => rgb <= "101000";
					when "00011101010101100" => rgb <= "101000";
					when "00011101010101101" => rgb <= "101000";
					when "00011101010101110" => rgb <= "101000";
					when "00011101010101111" => rgb <= "101000";
					when "00011101010110000" => rgb <= "101000";
					when "00011101010110001" => rgb <= "101000";
					when "00011101010110010" => rgb <= "101000";
					when "00011101010110011" => rgb <= "101000";
					when "00011101010110100" => rgb <= "101000";
					when "00011101010110101" => rgb <= "101000";
					when "00011101010110110" => rgb <= "101000";
					when "00011101010110111" => rgb <= "101000";
					when "00011101010111000" => rgb <= "101000";
					when "00011101010111001" => rgb <= "101000";
					when "00011101010111010" => rgb <= "101000";
					when "00011101010111011" => rgb <= "101000";
					when "00011101010111100" => rgb <= "101000";
					when "00011101010111101" => rgb <= "101000";
					when "00011101010111110" => rgb <= "101000";
					when "00011101010111111" => rgb <= "101000";
					when "00011101011000000" => rgb <= "100100";
					when "00011101011000001" => rgb <= "000000";
					when "00011101011000010" => rgb <= "000000";
					when "00011101011000011" => rgb <= "000000";
					when "00011101011000100" => rgb <= "000000";
					when "00011101011000101" => rgb <= "000000";
					when "00011101011000110" => rgb <= "000000";
					when "00011101011000111" => rgb <= "000000";
					when "00011101011001000" => rgb <= "000000";
					when "00011101011001001" => rgb <= "000000";
					when "00011101011001010" => rgb <= "000000";
					when "00011101011001011" => rgb <= "000000";
					when "00011101011001100" => rgb <= "000000";
					when "00011101011001101" => rgb <= "000000";
					when "00011101011001110" => rgb <= "000000";
					when "00011101011001111" => rgb <= "000000";
					when "00011101011010000" => rgb <= "000000";
					when "00011101011010001" => rgb <= "000000";
					when "00011101011010010" => rgb <= "000000";
					when "00011101011010011" => rgb <= "000000";
					when "00011101011010100" => rgb <= "000000";
					when "00011101011010101" => rgb <= "000000";
					when "00011101011010110" => rgb <= "000000";
					when "00011101011010111" => rgb <= "000000";
					when "00011101011011000" => rgb <= "000000";
					when "00011101011011001" => rgb <= "000000";
					when "00011101011011010" => rgb <= "000000";
					when "00011101011011011" => rgb <= "000000";
					when "00011101011011100" => rgb <= "000000";
					when "00011101011011101" => rgb <= "000000";
					when "00011101011011110" => rgb <= "000000";
					when "00011101011011111" => rgb <= "000000";
					when "00011101011100000" => rgb <= "000000";
					when "00011101011100001" => rgb <= "000000";
					when "00011101011100010" => rgb <= "000000";
					when "00011101011100011" => rgb <= "000000";
					when "00011101011100100" => rgb <= "000000";
					when "00011101011100101" => rgb <= "000000";
					when "00011101011100110" => rgb <= "000000";
					when "00011101011100111" => rgb <= "000000";
					when "00011101011101000" => rgb <= "000000";
					when "00011101011101001" => rgb <= "000000";
					when "00011101011101010" => rgb <= "000000";
					when "00011101011101011" => rgb <= "000000";
					when "00011101011101100" => rgb <= "000000";
					when "00011101011101101" => rgb <= "000000";
					when "00011101011101110" => rgb <= "000000";
					when "00011101011101111" => rgb <= "000000";
					when "00011101011110000" => rgb <= "000000";
					when "00011101011110001" => rgb <= "000000";
					when "00011101011110010" => rgb <= "000000";
					when "00011101011110011" => rgb <= "000000";
					when "00011101011110100" => rgb <= "000000";
					when "00011101011110101" => rgb <= "000000";
					when "00011101011110110" => rgb <= "000000";
					when "00011101011110111" => rgb <= "000000";
					when "00011101011111000" => rgb <= "000000";
					when "00011101011111001" => rgb <= "000000";
					when "00011101011111010" => rgb <= "000000";
					when "00011101011111011" => rgb <= "000000";
					when "00011101011111100" => rgb <= "000000";
					when "00011101011111101" => rgb <= "000000";
					when "00011101011111110" => rgb <= "000000";
					when "00011101011111111" => rgb <= "000000";
					when "00011101100000000" => rgb <= "000000";
					when "00011101100000001" => rgb <= "000000";
					when "00011101100000010" => rgb <= "000000";
					when "00011101100000011" => rgb <= "000000";
					when "00011101100000100" => rgb <= "000000";
					when "00011101100000101" => rgb <= "000000";
					when "00011101100000110" => rgb <= "000000";
					when "00011101100000111" => rgb <= "000000";
					when "00011101100001000" => rgb <= "000000";
					when "00011101100001001" => rgb <= "000000";
					when "00011101100001010" => rgb <= "000000";
					when "00011101100001011" => rgb <= "000000";
					when "00011101100001100" => rgb <= "000000";
					when "00011101100001101" => rgb <= "000000";
					when "00011101100001110" => rgb <= "000000";
					when "00011101100001111" => rgb <= "000000";
					when "00011101100010000" => rgb <= "000000";
					when "00011101100010001" => rgb <= "000000";
					when "00011101100010010" => rgb <= "000000";
					when "00011101100010011" => rgb <= "000000";
					when "00011101100010100" => rgb <= "000000";
					when "00011101100010101" => rgb <= "000000";
					when "00011101100010110" => rgb <= "000000";
					when "00011101100010111" => rgb <= "000000";
					when "00011101100011000" => rgb <= "000000";
					when "00011101100011001" => rgb <= "000000";
					when "00011101100011010" => rgb <= "000000";
					when "00011101100011011" => rgb <= "000000";
					when "00011101100011100" => rgb <= "000000";
					when "00011101100011101" => rgb <= "000000";
					when "00011101100011110" => rgb <= "000000";
					when "00011101100011111" => rgb <= "000000";
					when "00011101100100000" => rgb <= "000000";
					when "00011101100100001" => rgb <= "000000";
					when "00011101100100010" => rgb <= "000000";
					when "00011101100100011" => rgb <= "000000";
					when "00011101100100100" => rgb <= "000000";
					when "00011101100100101" => rgb <= "000000";
					when "00011101100100110" => rgb <= "000000";
					when "00011101100100111" => rgb <= "000000";
					when "00011101100101000" => rgb <= "000000";
					when "00011101100101001" => rgb <= "000000";
					when "00011101100101010" => rgb <= "000000";
					when "00011101100101011" => rgb <= "000000";
					when "00011101100101100" => rgb <= "000000";
					when "00011101100101101" => rgb <= "000000";
					when "00011101100101110" => rgb <= "000000";
					when "00011101100101111" => rgb <= "000000";
					when "00011101100110000" => rgb <= "000000";
					when "00011101100110001" => rgb <= "000000";
					when "00011101100110010" => rgb <= "000000";
					when "00011101100110011" => rgb <= "000000";
					when "00011101100110100" => rgb <= "000000";
					when "00011101100110101" => rgb <= "000000";
					when "00011101100110110" => rgb <= "000000";
					when "00011101100110111" => rgb <= "000000";
					when "00011101100111000" => rgb <= "000000";
					when "00011101100111001" => rgb <= "000000";
					when "00011101100111010" => rgb <= "000000";
					when "00011101100111011" => rgb <= "000000";
					when "00011101100111100" => rgb <= "000000";
					when "00011101100111101" => rgb <= "000000";
					when "00011101100111110" => rgb <= "000000";
					when "00011101100111111" => rgb <= "000000";
					when "00011110000000000" => rgb <= "000000";
					when "00011110000000001" => rgb <= "000000";
					when "00011110000000010" => rgb <= "000000";
					when "00011110000000011" => rgb <= "000000";
					when "00011110000000100" => rgb <= "000000";
					when "00011110000000101" => rgb <= "000000";
					when "00011110000000110" => rgb <= "000000";
					when "00011110000000111" => rgb <= "000000";
					when "00011110000001000" => rgb <= "000000";
					when "00011110000001001" => rgb <= "000000";
					when "00011110000001010" => rgb <= "000000";
					when "00011110000001011" => rgb <= "000000";
					when "00011110000001100" => rgb <= "000000";
					when "00011110000001101" => rgb <= "000000";
					when "00011110000001110" => rgb <= "000000";
					when "00011110000001111" => rgb <= "000000";
					when "00011110000010000" => rgb <= "000000";
					when "00011110000010001" => rgb <= "000000";
					when "00011110000010010" => rgb <= "000000";
					when "00011110000010011" => rgb <= "000000";
					when "00011110000010100" => rgb <= "000000";
					when "00011110000010101" => rgb <= "000000";
					when "00011110000010110" => rgb <= "000000";
					when "00011110000010111" => rgb <= "000000";
					when "00011110000011000" => rgb <= "000000";
					when "00011110000011001" => rgb <= "000000";
					when "00011110000011010" => rgb <= "000000";
					when "00011110000011011" => rgb <= "000000";
					when "00011110000011100" => rgb <= "000000";
					when "00011110000011101" => rgb <= "000000";
					when "00011110000011110" => rgb <= "000000";
					when "00011110000011111" => rgb <= "000000";
					when "00011110000100000" => rgb <= "000000";
					when "00011110000100001" => rgb <= "000000";
					when "00011110000100010" => rgb <= "000000";
					when "00011110000100011" => rgb <= "000000";
					when "00011110000100100" => rgb <= "000000";
					when "00011110000100101" => rgb <= "000000";
					when "00011110000100110" => rgb <= "000000";
					when "00011110000100111" => rgb <= "000000";
					when "00011110000101000" => rgb <= "000000";
					when "00011110000101001" => rgb <= "000000";
					when "00011110000101010" => rgb <= "000000";
					when "00011110000101011" => rgb <= "000000";
					when "00011110000101100" => rgb <= "000000";
					when "00011110000101101" => rgb <= "000000";
					when "00011110000101110" => rgb <= "000000";
					when "00011110000101111" => rgb <= "000000";
					when "00011110000110000" => rgb <= "000000";
					when "00011110000110001" => rgb <= "000000";
					when "00011110000110010" => rgb <= "000000";
					when "00011110000110011" => rgb <= "000000";
					when "00011110000110100" => rgb <= "000000";
					when "00011110000110101" => rgb <= "000000";
					when "00011110000110110" => rgb <= "000000";
					when "00011110000110111" => rgb <= "000000";
					when "00011110000111000" => rgb <= "000000";
					when "00011110000111001" => rgb <= "000000";
					when "00011110000111010" => rgb <= "000000";
					when "00011110000111011" => rgb <= "000000";
					when "00011110000111100" => rgb <= "000000";
					when "00011110000111101" => rgb <= "000000";
					when "00011110000111110" => rgb <= "000000";
					when "00011110000111111" => rgb <= "000000";
					when "00011110001000000" => rgb <= "000000";
					when "00011110001000001" => rgb <= "000000";
					when "00011110001000010" => rgb <= "000000";
					when "00011110001000011" => rgb <= "000000";
					when "00011110001000100" => rgb <= "000000";
					when "00011110001000101" => rgb <= "000000";
					when "00011110001000110" => rgb <= "000000";
					when "00011110001000111" => rgb <= "000000";
					when "00011110001001000" => rgb <= "000000";
					when "00011110001001001" => rgb <= "000000";
					when "00011110001001010" => rgb <= "000000";
					when "00011110001001011" => rgb <= "000000";
					when "00011110001001100" => rgb <= "000000";
					when "00011110001001101" => rgb <= "000000";
					when "00011110001001110" => rgb <= "000000";
					when "00011110001001111" => rgb <= "000000";
					when "00011110001010000" => rgb <= "000000";
					when "00011110001010001" => rgb <= "000000";
					when "00011110001010010" => rgb <= "000000";
					when "00011110001010011" => rgb <= "000000";
					when "00011110001010100" => rgb <= "000000";
					when "00011110001010101" => rgb <= "000000";
					when "00011110001010110" => rgb <= "000000";
					when "00011110001010111" => rgb <= "000000";
					when "00011110001011000" => rgb <= "000000";
					when "00011110001011001" => rgb <= "000000";
					when "00011110001011010" => rgb <= "000000";
					when "00011110001011011" => rgb <= "000000";
					when "00011110001011100" => rgb <= "000000";
					when "00011110001011101" => rgb <= "000000";
					when "00011110001011110" => rgb <= "000000";
					when "00011110001011111" => rgb <= "000000";
					when "00011110001100000" => rgb <= "000000";
					when "00011110001100001" => rgb <= "000000";
					when "00011110001100010" => rgb <= "000000";
					when "00011110001100011" => rgb <= "000000";
					when "00011110001100100" => rgb <= "000000";
					when "00011110001100101" => rgb <= "000000";
					when "00011110001100110" => rgb <= "000000";
					when "00011110001100111" => rgb <= "000000";
					when "00011110001101000" => rgb <= "000000";
					when "00011110001101001" => rgb <= "000000";
					when "00011110001101010" => rgb <= "000000";
					when "00011110001101011" => rgb <= "000000";
					when "00011110001101100" => rgb <= "000000";
					when "00011110001101101" => rgb <= "000000";
					when "00011110001101110" => rgb <= "000000";
					when "00011110001101111" => rgb <= "000000";
					when "00011110001110000" => rgb <= "000000";
					when "00011110001110001" => rgb <= "000000";
					when "00011110001110010" => rgb <= "000000";
					when "00011110001110011" => rgb <= "000000";
					when "00011110001110100" => rgb <= "000000";
					when "00011110001110101" => rgb <= "000000";
					when "00011110001110110" => rgb <= "000000";
					when "00011110001110111" => rgb <= "000000";
					when "00011110001111000" => rgb <= "000000";
					when "00011110001111001" => rgb <= "000000";
					when "00011110001111010" => rgb <= "000000";
					when "00011110001111011" => rgb <= "000000";
					when "00011110001111100" => rgb <= "000000";
					when "00011110001111101" => rgb <= "101000";
					when "00011110001111110" => rgb <= "101000";
					when "00011110001111111" => rgb <= "101000";
					when "00011110010000000" => rgb <= "101000";
					when "00011110010000001" => rgb <= "101000";
					when "00011110010000010" => rgb <= "101000";
					when "00011110010000011" => rgb <= "101000";
					when "00011110010000100" => rgb <= "101000";
					when "00011110010000101" => rgb <= "101000";
					when "00011110010000110" => rgb <= "101000";
					when "00011110010000111" => rgb <= "101000";
					when "00011110010001000" => rgb <= "101001";
					when "00011110010001001" => rgb <= "101001";
					when "00011110010001010" => rgb <= "111001";
					when "00011110010001011" => rgb <= "101001";
					when "00011110010001100" => rgb <= "101001";
					when "00011110010001101" => rgb <= "111001";
					when "00011110010001110" => rgb <= "101001";
					when "00011110010001111" => rgb <= "111001";
					when "00011110010010000" => rgb <= "101001";
					when "00011110010010001" => rgb <= "101001";
					when "00011110010010010" => rgb <= "101001";
					when "00011110010010011" => rgb <= "101001";
					when "00011110010010100" => rgb <= "101001";
					when "00011110010010101" => rgb <= "101001";
					when "00011110010010110" => rgb <= "101001";
					when "00011110010010111" => rgb <= "101001";
					when "00011110010011000" => rgb <= "101001";
					when "00011110010011001" => rgb <= "101001";
					when "00011110010011010" => rgb <= "111001";
					when "00011110010011011" => rgb <= "111001";
					when "00011110010011100" => rgb <= "101001";
					when "00011110010011101" => rgb <= "111001";
					when "00011110010011110" => rgb <= "111001";
					when "00011110010011111" => rgb <= "101000";
					when "00011110010100000" => rgb <= "101000";
					when "00011110010100001" => rgb <= "101000";
					when "00011110010100010" => rgb <= "101000";
					when "00011110010100011" => rgb <= "101000";
					when "00011110010100100" => rgb <= "101000";
					when "00011110010100101" => rgb <= "101000";
					when "00011110010100110" => rgb <= "101000";
					when "00011110010100111" => rgb <= "101000";
					when "00011110010101000" => rgb <= "101000";
					when "00011110010101001" => rgb <= "101000";
					when "00011110010101010" => rgb <= "101000";
					when "00011110010101011" => rgb <= "101000";
					when "00011110010101100" => rgb <= "101000";
					when "00011110010101101" => rgb <= "101000";
					when "00011110010101110" => rgb <= "101000";
					when "00011110010101111" => rgb <= "101000";
					when "00011110010110000" => rgb <= "101000";
					when "00011110010110001" => rgb <= "101000";
					when "00011110010110010" => rgb <= "101000";
					when "00011110010110011" => rgb <= "101000";
					when "00011110010110100" => rgb <= "101000";
					when "00011110010110101" => rgb <= "101000";
					when "00011110010110110" => rgb <= "101000";
					when "00011110010110111" => rgb <= "101000";
					when "00011110010111000" => rgb <= "101000";
					when "00011110010111001" => rgb <= "101000";
					when "00011110010111010" => rgb <= "101000";
					when "00011110010111011" => rgb <= "101000";
					when "00011110010111100" => rgb <= "101000";
					when "00011110010111101" => rgb <= "101000";
					when "00011110010111110" => rgb <= "101000";
					when "00011110010111111" => rgb <= "101000";
					when "00011110011000000" => rgb <= "100100";
					when "00011110011000001" => rgb <= "000000";
					when "00011110011000010" => rgb <= "000000";
					when "00011110011000011" => rgb <= "000000";
					when "00011110011000100" => rgb <= "000000";
					when "00011110011000101" => rgb <= "000000";
					when "00011110011000110" => rgb <= "000000";
					when "00011110011000111" => rgb <= "000000";
					when "00011110011001000" => rgb <= "000000";
					when "00011110011001001" => rgb <= "000000";
					when "00011110011001010" => rgb <= "000000";
					when "00011110011001011" => rgb <= "000000";
					when "00011110011001100" => rgb <= "000000";
					when "00011110011001101" => rgb <= "000000";
					when "00011110011001110" => rgb <= "000000";
					when "00011110011001111" => rgb <= "000000";
					when "00011110011010000" => rgb <= "000000";
					when "00011110011010001" => rgb <= "000000";
					when "00011110011010010" => rgb <= "000000";
					when "00011110011010011" => rgb <= "000000";
					when "00011110011010100" => rgb <= "000000";
					when "00011110011010101" => rgb <= "000000";
					when "00011110011010110" => rgb <= "000000";
					when "00011110011010111" => rgb <= "000000";
					when "00011110011011000" => rgb <= "000000";
					when "00011110011011001" => rgb <= "000000";
					when "00011110011011010" => rgb <= "000000";
					when "00011110011011011" => rgb <= "000000";
					when "00011110011011100" => rgb <= "000000";
					when "00011110011011101" => rgb <= "000000";
					when "00011110011011110" => rgb <= "000000";
					when "00011110011011111" => rgb <= "000000";
					when "00011110011100000" => rgb <= "000000";
					when "00011110011100001" => rgb <= "000000";
					when "00011110011100010" => rgb <= "000000";
					when "00011110011100011" => rgb <= "000000";
					when "00011110011100100" => rgb <= "000000";
					when "00011110011100101" => rgb <= "000000";
					when "00011110011100110" => rgb <= "000000";
					when "00011110011100111" => rgb <= "000000";
					when "00011110011101000" => rgb <= "000000";
					when "00011110011101001" => rgb <= "000000";
					when "00011110011101010" => rgb <= "000000";
					when "00011110011101011" => rgb <= "000000";
					when "00011110011101100" => rgb <= "000000";
					when "00011110011101101" => rgb <= "000000";
					when "00011110011101110" => rgb <= "000000";
					when "00011110011101111" => rgb <= "000000";
					when "00011110011110000" => rgb <= "000000";
					when "00011110011110001" => rgb <= "000000";
					when "00011110011110010" => rgb <= "000000";
					when "00011110011110011" => rgb <= "000000";
					when "00011110011110100" => rgb <= "000000";
					when "00011110011110101" => rgb <= "000000";
					when "00011110011110110" => rgb <= "000000";
					when "00011110011110111" => rgb <= "000000";
					when "00011110011111000" => rgb <= "000000";
					when "00011110011111001" => rgb <= "000000";
					when "00011110011111010" => rgb <= "000000";
					when "00011110011111011" => rgb <= "000000";
					when "00011110011111100" => rgb <= "000000";
					when "00011110011111101" => rgb <= "000000";
					when "00011110011111110" => rgb <= "000000";
					when "00011110011111111" => rgb <= "000000";
					when "00011110100000000" => rgb <= "000000";
					when "00011110100000001" => rgb <= "000000";
					when "00011110100000010" => rgb <= "000000";
					when "00011110100000011" => rgb <= "000000";
					when "00011110100000100" => rgb <= "000000";
					when "00011110100000101" => rgb <= "000000";
					when "00011110100000110" => rgb <= "000000";
					when "00011110100000111" => rgb <= "000000";
					when "00011110100001000" => rgb <= "000000";
					when "00011110100001001" => rgb <= "000000";
					when "00011110100001010" => rgb <= "000000";
					when "00011110100001011" => rgb <= "000000";
					when "00011110100001100" => rgb <= "000000";
					when "00011110100001101" => rgb <= "000000";
					when "00011110100001110" => rgb <= "000000";
					when "00011110100001111" => rgb <= "000000";
					when "00011110100010000" => rgb <= "000000";
					when "00011110100010001" => rgb <= "000000";
					when "00011110100010010" => rgb <= "000000";
					when "00011110100010011" => rgb <= "000000";
					when "00011110100010100" => rgb <= "000000";
					when "00011110100010101" => rgb <= "000000";
					when "00011110100010110" => rgb <= "000000";
					when "00011110100010111" => rgb <= "000000";
					when "00011110100011000" => rgb <= "000000";
					when "00011110100011001" => rgb <= "000000";
					when "00011110100011010" => rgb <= "000000";
					when "00011110100011011" => rgb <= "000000";
					when "00011110100011100" => rgb <= "000000";
					when "00011110100011101" => rgb <= "000000";
					when "00011110100011110" => rgb <= "000000";
					when "00011110100011111" => rgb <= "000000";
					when "00011110100100000" => rgb <= "000000";
					when "00011110100100001" => rgb <= "000000";
					when "00011110100100010" => rgb <= "000000";
					when "00011110100100011" => rgb <= "000000";
					when "00011110100100100" => rgb <= "000000";
					when "00011110100100101" => rgb <= "000000";
					when "00011110100100110" => rgb <= "000000";
					when "00011110100100111" => rgb <= "000000";
					when "00011110100101000" => rgb <= "000000";
					when "00011110100101001" => rgb <= "000000";
					when "00011110100101010" => rgb <= "000000";
					when "00011110100101011" => rgb <= "000000";
					when "00011110100101100" => rgb <= "000000";
					when "00011110100101101" => rgb <= "000000";
					when "00011110100101110" => rgb <= "000000";
					when "00011110100101111" => rgb <= "000000";
					when "00011110100110000" => rgb <= "000000";
					when "00011110100110001" => rgb <= "000000";
					when "00011110100110010" => rgb <= "000000";
					when "00011110100110011" => rgb <= "000000";
					when "00011110100110100" => rgb <= "000000";
					when "00011110100110101" => rgb <= "000000";
					when "00011110100110110" => rgb <= "000000";
					when "00011110100110111" => rgb <= "000000";
					when "00011110100111000" => rgb <= "000000";
					when "00011110100111001" => rgb <= "000000";
					when "00011110100111010" => rgb <= "000000";
					when "00011110100111011" => rgb <= "000000";
					when "00011110100111100" => rgb <= "000000";
					when "00011110100111101" => rgb <= "000000";
					when "00011110100111110" => rgb <= "000000";
					when "00011110100111111" => rgb <= "000000";
					when "00011111000000000" => rgb <= "000000";
					when "00011111000000001" => rgb <= "000000";
					when "00011111000000010" => rgb <= "000000";
					when "00011111000000011" => rgb <= "000000";
					when "00011111000000100" => rgb <= "000000";
					when "00011111000000101" => rgb <= "000000";
					when "00011111000000110" => rgb <= "000000";
					when "00011111000000111" => rgb <= "000000";
					when "00011111000001000" => rgb <= "000000";
					when "00011111000001001" => rgb <= "000000";
					when "00011111000001010" => rgb <= "000000";
					when "00011111000001011" => rgb <= "000000";
					when "00011111000001100" => rgb <= "000000";
					when "00011111000001101" => rgb <= "000000";
					when "00011111000001110" => rgb <= "000000";
					when "00011111000001111" => rgb <= "000000";
					when "00011111000010000" => rgb <= "000000";
					when "00011111000010001" => rgb <= "000000";
					when "00011111000010010" => rgb <= "000000";
					when "00011111000010011" => rgb <= "000000";
					when "00011111000010100" => rgb <= "000000";
					when "00011111000010101" => rgb <= "000000";
					when "00011111000010110" => rgb <= "000000";
					when "00011111000010111" => rgb <= "000000";
					when "00011111000011000" => rgb <= "000000";
					when "00011111000011001" => rgb <= "000000";
					when "00011111000011010" => rgb <= "000000";
					when "00011111000011011" => rgb <= "000000";
					when "00011111000011100" => rgb <= "000000";
					when "00011111000011101" => rgb <= "000000";
					when "00011111000011110" => rgb <= "000000";
					when "00011111000011111" => rgb <= "000000";
					when "00011111000100000" => rgb <= "000000";
					when "00011111000100001" => rgb <= "000000";
					when "00011111000100010" => rgb <= "000000";
					when "00011111000100011" => rgb <= "000000";
					when "00011111000100100" => rgb <= "000000";
					when "00011111000100101" => rgb <= "000000";
					when "00011111000100110" => rgb <= "000000";
					when "00011111000100111" => rgb <= "000000";
					when "00011111000101000" => rgb <= "000000";
					when "00011111000101001" => rgb <= "000000";
					when "00011111000101010" => rgb <= "000000";
					when "00011111000101011" => rgb <= "000000";
					when "00011111000101100" => rgb <= "000000";
					when "00011111000101101" => rgb <= "000000";
					when "00011111000101110" => rgb <= "000000";
					when "00011111000101111" => rgb <= "000000";
					when "00011111000110000" => rgb <= "000000";
					when "00011111000110001" => rgb <= "000000";
					when "00011111000110010" => rgb <= "000000";
					when "00011111000110011" => rgb <= "000000";
					when "00011111000110100" => rgb <= "000000";
					when "00011111000110101" => rgb <= "000000";
					when "00011111000110110" => rgb <= "000000";
					when "00011111000110111" => rgb <= "000000";
					when "00011111000111000" => rgb <= "000000";
					when "00011111000111001" => rgb <= "000000";
					when "00011111000111010" => rgb <= "000000";
					when "00011111000111011" => rgb <= "000000";
					when "00011111000111100" => rgb <= "000000";
					when "00011111000111101" => rgb <= "000000";
					when "00011111000111110" => rgb <= "000000";
					when "00011111000111111" => rgb <= "000000";
					when "00011111001000000" => rgb <= "000000";
					when "00011111001000001" => rgb <= "000000";
					when "00011111001000010" => rgb <= "000000";
					when "00011111001000011" => rgb <= "000000";
					when "00011111001000100" => rgb <= "000000";
					when "00011111001000101" => rgb <= "000000";
					when "00011111001000110" => rgb <= "000000";
					when "00011111001000111" => rgb <= "000000";
					when "00011111001001000" => rgb <= "000000";
					when "00011111001001001" => rgb <= "000000";
					when "00011111001001010" => rgb <= "000000";
					when "00011111001001011" => rgb <= "000000";
					when "00011111001001100" => rgb <= "000000";
					when "00011111001001101" => rgb <= "000000";
					when "00011111001001110" => rgb <= "000000";
					when "00011111001001111" => rgb <= "000000";
					when "00011111001010000" => rgb <= "000000";
					when "00011111001010001" => rgb <= "000000";
					when "00011111001010010" => rgb <= "000000";
					when "00011111001010011" => rgb <= "000000";
					when "00011111001010100" => rgb <= "000000";
					when "00011111001010101" => rgb <= "000000";
					when "00011111001010110" => rgb <= "000000";
					when "00011111001010111" => rgb <= "000000";
					when "00011111001011000" => rgb <= "000000";
					when "00011111001011001" => rgb <= "000000";
					when "00011111001011010" => rgb <= "000000";
					when "00011111001011011" => rgb <= "000000";
					when "00011111001011100" => rgb <= "000000";
					when "00011111001011101" => rgb <= "000000";
					when "00011111001011110" => rgb <= "000000";
					when "00011111001011111" => rgb <= "000000";
					when "00011111001100000" => rgb <= "000000";
					when "00011111001100001" => rgb <= "000000";
					when "00011111001100010" => rgb <= "000000";
					when "00011111001100011" => rgb <= "000000";
					when "00011111001100100" => rgb <= "000000";
					when "00011111001100101" => rgb <= "000000";
					when "00011111001100110" => rgb <= "000000";
					when "00011111001100111" => rgb <= "000000";
					when "00011111001101000" => rgb <= "000000";
					when "00011111001101001" => rgb <= "000000";
					when "00011111001101010" => rgb <= "000000";
					when "00011111001101011" => rgb <= "000000";
					when "00011111001101100" => rgb <= "000000";
					when "00011111001101101" => rgb <= "000000";
					when "00011111001101110" => rgb <= "000000";
					when "00011111001101111" => rgb <= "000000";
					when "00011111001110000" => rgb <= "000000";
					when "00011111001110001" => rgb <= "000000";
					when "00011111001110010" => rgb <= "000000";
					when "00011111001110011" => rgb <= "000000";
					when "00011111001110100" => rgb <= "000000";
					when "00011111001110101" => rgb <= "000000";
					when "00011111001110110" => rgb <= "000000";
					when "00011111001110111" => rgb <= "000000";
					when "00011111001111000" => rgb <= "000000";
					when "00011111001111001" => rgb <= "000000";
					when "00011111001111010" => rgb <= "000000";
					when "00011111001111011" => rgb <= "000000";
					when "00011111001111100" => rgb <= "000000";
					when "00011111001111101" => rgb <= "101000";
					when "00011111001111110" => rgb <= "101000";
					when "00011111001111111" => rgb <= "101000";
					when "00011111010000000" => rgb <= "101000";
					when "00011111010000001" => rgb <= "101000";
					when "00011111010000010" => rgb <= "101000";
					when "00011111010000011" => rgb <= "101000";
					when "00011111010000100" => rgb <= "101000";
					when "00011111010000101" => rgb <= "101000";
					when "00011111010000110" => rgb <= "101000";
					when "00011111010000111" => rgb <= "101000";
					when "00011111010001000" => rgb <= "101001";
					when "00011111010001001" => rgb <= "101001";
					when "00011111010001010" => rgb <= "111001";
					when "00011111010001011" => rgb <= "101010";
					when "00011111010001100" => rgb <= "101001";
					when "00011111010001101" => rgb <= "111001";
					when "00011111010001110" => rgb <= "111001";
					when "00011111010001111" => rgb <= "111010";
					when "00011111010010000" => rgb <= "101001";
					when "00011111010010001" => rgb <= "101001";
					when "00011111010010010" => rgb <= "101001";
					when "00011111010010011" => rgb <= "101001";
					when "00011111010010100" => rgb <= "101001";
					when "00011111010010101" => rgb <= "101001";
					when "00011111010010110" => rgb <= "101001";
					when "00011111010010111" => rgb <= "101001";
					when "00011111010011000" => rgb <= "101001";
					when "00011111010011001" => rgb <= "101001";
					when "00011111010011010" => rgb <= "111001";
					when "00011111010011011" => rgb <= "111001";
					when "00011111010011100" => rgb <= "101001";
					when "00011111010011101" => rgb <= "111010";
					when "00011111010011110" => rgb <= "111001";
					when "00011111010011111" => rgb <= "101000";
					when "00011111010100000" => rgb <= "101000";
					when "00011111010100001" => rgb <= "101000";
					when "00011111010100010" => rgb <= "101000";
					when "00011111010100011" => rgb <= "101000";
					when "00011111010100100" => rgb <= "101000";
					when "00011111010100101" => rgb <= "101000";
					when "00011111010100110" => rgb <= "101000";
					when "00011111010100111" => rgb <= "101000";
					when "00011111010101000" => rgb <= "101000";
					when "00011111010101001" => rgb <= "101000";
					when "00011111010101010" => rgb <= "101000";
					when "00011111010101011" => rgb <= "101000";
					when "00011111010101100" => rgb <= "101000";
					when "00011111010101101" => rgb <= "101000";
					when "00011111010101110" => rgb <= "101000";
					when "00011111010101111" => rgb <= "101000";
					when "00011111010110000" => rgb <= "101000";
					when "00011111010110001" => rgb <= "101000";
					when "00011111010110010" => rgb <= "101000";
					when "00011111010110011" => rgb <= "101000";
					when "00011111010110100" => rgb <= "101000";
					when "00011111010110101" => rgb <= "101000";
					when "00011111010110110" => rgb <= "101000";
					when "00011111010110111" => rgb <= "101000";
					when "00011111010111000" => rgb <= "101000";
					when "00011111010111001" => rgb <= "101000";
					when "00011111010111010" => rgb <= "101000";
					when "00011111010111011" => rgb <= "101000";
					when "00011111010111100" => rgb <= "101000";
					when "00011111010111101" => rgb <= "101000";
					when "00011111010111110" => rgb <= "101000";
					when "00011111010111111" => rgb <= "101000";
					when "00011111011000000" => rgb <= "100100";
					when "00011111011000001" => rgb <= "000000";
					when "00011111011000010" => rgb <= "000000";
					when "00011111011000011" => rgb <= "000000";
					when "00011111011000100" => rgb <= "000000";
					when "00011111011000101" => rgb <= "000000";
					when "00011111011000110" => rgb <= "000000";
					when "00011111011000111" => rgb <= "000000";
					when "00011111011001000" => rgb <= "000000";
					when "00011111011001001" => rgb <= "000000";
					when "00011111011001010" => rgb <= "000000";
					when "00011111011001011" => rgb <= "000000";
					when "00011111011001100" => rgb <= "000000";
					when "00011111011001101" => rgb <= "000000";
					when "00011111011001110" => rgb <= "000000";
					when "00011111011001111" => rgb <= "000000";
					when "00011111011010000" => rgb <= "000000";
					when "00011111011010001" => rgb <= "000000";
					when "00011111011010010" => rgb <= "000000";
					when "00011111011010011" => rgb <= "000000";
					when "00011111011010100" => rgb <= "000000";
					when "00011111011010101" => rgb <= "000000";
					when "00011111011010110" => rgb <= "000000";
					when "00011111011010111" => rgb <= "000000";
					when "00011111011011000" => rgb <= "000000";
					when "00011111011011001" => rgb <= "000000";
					when "00011111011011010" => rgb <= "000000";
					when "00011111011011011" => rgb <= "000000";
					when "00011111011011100" => rgb <= "000000";
					when "00011111011011101" => rgb <= "000000";
					when "00011111011011110" => rgb <= "000000";
					when "00011111011011111" => rgb <= "000000";
					when "00011111011100000" => rgb <= "000000";
					when "00011111011100001" => rgb <= "000000";
					when "00011111011100010" => rgb <= "000000";
					when "00011111011100011" => rgb <= "000000";
					when "00011111011100100" => rgb <= "000000";
					when "00011111011100101" => rgb <= "000000";
					when "00011111011100110" => rgb <= "000000";
					when "00011111011100111" => rgb <= "000000";
					when "00011111011101000" => rgb <= "000000";
					when "00011111011101001" => rgb <= "000000";
					when "00011111011101010" => rgb <= "000000";
					when "00011111011101011" => rgb <= "000000";
					when "00011111011101100" => rgb <= "000000";
					when "00011111011101101" => rgb <= "000000";
					when "00011111011101110" => rgb <= "000000";
					when "00011111011101111" => rgb <= "000000";
					when "00011111011110000" => rgb <= "000000";
					when "00011111011110001" => rgb <= "000000";
					when "00011111011110010" => rgb <= "000000";
					when "00011111011110011" => rgb <= "000000";
					when "00011111011110100" => rgb <= "000000";
					when "00011111011110101" => rgb <= "000000";
					when "00011111011110110" => rgb <= "000000";
					when "00011111011110111" => rgb <= "000000";
					when "00011111011111000" => rgb <= "000000";
					when "00011111011111001" => rgb <= "000000";
					when "00011111011111010" => rgb <= "000000";
					when "00011111011111011" => rgb <= "000000";
					when "00011111011111100" => rgb <= "000000";
					when "00011111011111101" => rgb <= "000000";
					when "00011111011111110" => rgb <= "000000";
					when "00011111011111111" => rgb <= "000000";
					when "00011111100000000" => rgb <= "000000";
					when "00011111100000001" => rgb <= "000000";
					when "00011111100000010" => rgb <= "000000";
					when "00011111100000011" => rgb <= "000000";
					when "00011111100000100" => rgb <= "000000";
					when "00011111100000101" => rgb <= "000000";
					when "00011111100000110" => rgb <= "000000";
					when "00011111100000111" => rgb <= "000000";
					when "00011111100001000" => rgb <= "000000";
					when "00011111100001001" => rgb <= "000000";
					when "00011111100001010" => rgb <= "000000";
					when "00011111100001011" => rgb <= "000000";
					when "00011111100001100" => rgb <= "000000";
					when "00011111100001101" => rgb <= "000000";
					when "00011111100001110" => rgb <= "000000";
					when "00011111100001111" => rgb <= "000000";
					when "00011111100010000" => rgb <= "000000";
					when "00011111100010001" => rgb <= "000000";
					when "00011111100010010" => rgb <= "000000";
					when "00011111100010011" => rgb <= "000000";
					when "00011111100010100" => rgb <= "000000";
					when "00011111100010101" => rgb <= "000000";
					when "00011111100010110" => rgb <= "000000";
					when "00011111100010111" => rgb <= "000000";
					when "00011111100011000" => rgb <= "000000";
					when "00011111100011001" => rgb <= "000000";
					when "00011111100011010" => rgb <= "000000";
					when "00011111100011011" => rgb <= "000000";
					when "00011111100011100" => rgb <= "000000";
					when "00011111100011101" => rgb <= "000000";
					when "00011111100011110" => rgb <= "000000";
					when "00011111100011111" => rgb <= "000000";
					when "00011111100100000" => rgb <= "000000";
					when "00011111100100001" => rgb <= "000000";
					when "00011111100100010" => rgb <= "000000";
					when "00011111100100011" => rgb <= "000000";
					when "00011111100100100" => rgb <= "000000";
					when "00011111100100101" => rgb <= "000000";
					when "00011111100100110" => rgb <= "000000";
					when "00011111100100111" => rgb <= "000000";
					when "00011111100101000" => rgb <= "000000";
					when "00011111100101001" => rgb <= "000000";
					when "00011111100101010" => rgb <= "000000";
					when "00011111100101011" => rgb <= "000000";
					when "00011111100101100" => rgb <= "000000";
					when "00011111100101101" => rgb <= "000000";
					when "00011111100101110" => rgb <= "000000";
					when "00011111100101111" => rgb <= "000000";
					when "00011111100110000" => rgb <= "000000";
					when "00011111100110001" => rgb <= "000000";
					when "00011111100110010" => rgb <= "000000";
					when "00011111100110011" => rgb <= "000000";
					when "00011111100110100" => rgb <= "000000";
					when "00011111100110101" => rgb <= "000000";
					when "00011111100110110" => rgb <= "000000";
					when "00011111100110111" => rgb <= "000000";
					when "00011111100111000" => rgb <= "000000";
					when "00011111100111001" => rgb <= "000000";
					when "00011111100111010" => rgb <= "000000";
					when "00011111100111011" => rgb <= "000000";
					when "00011111100111100" => rgb <= "000000";
					when "00011111100111101" => rgb <= "000000";
					when "00011111100111110" => rgb <= "000000";
					when "00011111100111111" => rgb <= "000000";
					when "00100000000000000" => rgb <= "000000";
					when "00100000000000001" => rgb <= "000000";
					when "00100000000000010" => rgb <= "000000";
					when "00100000000000011" => rgb <= "000000";
					when "00100000000000100" => rgb <= "000000";
					when "00100000000000101" => rgb <= "000000";
					when "00100000000000110" => rgb <= "000000";
					when "00100000000000111" => rgb <= "000000";
					when "00100000000001000" => rgb <= "000000";
					when "00100000000001001" => rgb <= "000000";
					when "00100000000001010" => rgb <= "000000";
					when "00100000000001011" => rgb <= "000000";
					when "00100000000001100" => rgb <= "000000";
					when "00100000000001101" => rgb <= "000000";
					when "00100000000001110" => rgb <= "000000";
					when "00100000000001111" => rgb <= "000000";
					when "00100000000010000" => rgb <= "000000";
					when "00100000000010001" => rgb <= "000000";
					when "00100000000010010" => rgb <= "000000";
					when "00100000000010011" => rgb <= "000000";
					when "00100000000010100" => rgb <= "000000";
					when "00100000000010101" => rgb <= "000000";
					when "00100000000010110" => rgb <= "000000";
					when "00100000000010111" => rgb <= "000000";
					when "00100000000011000" => rgb <= "000000";
					when "00100000000011001" => rgb <= "000000";
					when "00100000000011010" => rgb <= "000000";
					when "00100000000011011" => rgb <= "000000";
					when "00100000000011100" => rgb <= "000000";
					when "00100000000011101" => rgb <= "000000";
					when "00100000000011110" => rgb <= "000000";
					when "00100000000011111" => rgb <= "000000";
					when "00100000000100000" => rgb <= "000000";
					when "00100000000100001" => rgb <= "000000";
					when "00100000000100010" => rgb <= "000000";
					when "00100000000100011" => rgb <= "000000";
					when "00100000000100100" => rgb <= "000000";
					when "00100000000100101" => rgb <= "000000";
					when "00100000000100110" => rgb <= "000000";
					when "00100000000100111" => rgb <= "000000";
					when "00100000000101000" => rgb <= "000000";
					when "00100000000101001" => rgb <= "000000";
					when "00100000000101010" => rgb <= "000000";
					when "00100000000101011" => rgb <= "000000";
					when "00100000000101100" => rgb <= "000000";
					when "00100000000101101" => rgb <= "000000";
					when "00100000000101110" => rgb <= "000000";
					when "00100000000101111" => rgb <= "000000";
					when "00100000000110000" => rgb <= "000000";
					when "00100000000110001" => rgb <= "000000";
					when "00100000000110010" => rgb <= "000000";
					when "00100000000110011" => rgb <= "000000";
					when "00100000000110100" => rgb <= "000000";
					when "00100000000110101" => rgb <= "000000";
					when "00100000000110110" => rgb <= "000000";
					when "00100000000110111" => rgb <= "000000";
					when "00100000000111000" => rgb <= "000000";
					when "00100000000111001" => rgb <= "000000";
					when "00100000000111010" => rgb <= "000000";
					when "00100000000111011" => rgb <= "000000";
					when "00100000000111100" => rgb <= "000000";
					when "00100000000111101" => rgb <= "000000";
					when "00100000000111110" => rgb <= "000000";
					when "00100000000111111" => rgb <= "000000";
					when "00100000001000000" => rgb <= "000000";
					when "00100000001000001" => rgb <= "000000";
					when "00100000001000010" => rgb <= "000000";
					when "00100000001000011" => rgb <= "000000";
					when "00100000001000100" => rgb <= "000000";
					when "00100000001000101" => rgb <= "000000";
					when "00100000001000110" => rgb <= "000000";
					when "00100000001000111" => rgb <= "000000";
					when "00100000001001000" => rgb <= "000000";
					when "00100000001001001" => rgb <= "000000";
					when "00100000001001010" => rgb <= "000000";
					when "00100000001001011" => rgb <= "000000";
					when "00100000001001100" => rgb <= "000000";
					when "00100000001001101" => rgb <= "000000";
					when "00100000001001110" => rgb <= "000000";
					when "00100000001001111" => rgb <= "000000";
					when "00100000001010000" => rgb <= "000000";
					when "00100000001010001" => rgb <= "000000";
					when "00100000001010010" => rgb <= "000000";
					when "00100000001010011" => rgb <= "000000";
					when "00100000001010100" => rgb <= "000000";
					when "00100000001010101" => rgb <= "000000";
					when "00100000001010110" => rgb <= "000000";
					when "00100000001010111" => rgb <= "000000";
					when "00100000001011000" => rgb <= "000000";
					when "00100000001011001" => rgb <= "000000";
					when "00100000001011010" => rgb <= "000000";
					when "00100000001011011" => rgb <= "000000";
					when "00100000001011100" => rgb <= "000000";
					when "00100000001011101" => rgb <= "000000";
					when "00100000001011110" => rgb <= "000000";
					when "00100000001011111" => rgb <= "000000";
					when "00100000001100000" => rgb <= "000000";
					when "00100000001100001" => rgb <= "000000";
					when "00100000001100010" => rgb <= "000000";
					when "00100000001100011" => rgb <= "000000";
					when "00100000001100100" => rgb <= "000000";
					when "00100000001100101" => rgb <= "000000";
					when "00100000001100110" => rgb <= "000000";
					when "00100000001100111" => rgb <= "000000";
					when "00100000001101000" => rgb <= "000000";
					when "00100000001101001" => rgb <= "000000";
					when "00100000001101010" => rgb <= "000000";
					when "00100000001101011" => rgb <= "000000";
					when "00100000001101100" => rgb <= "000000";
					when "00100000001101101" => rgb <= "000000";
					when "00100000001101110" => rgb <= "000000";
					when "00100000001101111" => rgb <= "000000";
					when "00100000001110000" => rgb <= "000000";
					when "00100000001110001" => rgb <= "000000";
					when "00100000001110010" => rgb <= "000000";
					when "00100000001110011" => rgb <= "000000";
					when "00100000001110100" => rgb <= "000000";
					when "00100000001110101" => rgb <= "000000";
					when "00100000001110110" => rgb <= "000000";
					when "00100000001110111" => rgb <= "000000";
					when "00100000001111000" => rgb <= "000000";
					when "00100000001111001" => rgb <= "000000";
					when "00100000001111010" => rgb <= "000000";
					when "00100000001111011" => rgb <= "000000";
					when "00100000001111100" => rgb <= "000000";
					when "00100000001111101" => rgb <= "101000";
					when "00100000001111110" => rgb <= "101000";
					when "00100000001111111" => rgb <= "101000";
					when "00100000010000000" => rgb <= "101000";
					when "00100000010000001" => rgb <= "101000";
					when "00100000010000010" => rgb <= "101000";
					when "00100000010000011" => rgb <= "101000";
					when "00100000010000100" => rgb <= "101000";
					when "00100000010000101" => rgb <= "101000";
					when "00100000010000110" => rgb <= "101000";
					when "00100000010000111" => rgb <= "101000";
					when "00100000010001000" => rgb <= "101001";
					when "00100000010001001" => rgb <= "111001";
					when "00100000010001010" => rgb <= "101001";
					when "00100000010001011" => rgb <= "101001";
					when "00100000010001100" => rgb <= "111001";
					when "00100000010001101" => rgb <= "111001";
					when "00100000010001110" => rgb <= "111001";
					when "00100000010001111" => rgb <= "101001";
					when "00100000010010000" => rgb <= "111001";
					when "00100000010010001" => rgb <= "111001";
					when "00100000010010010" => rgb <= "111001";
					when "00100000010010011" => rgb <= "111001";
					when "00100000010010100" => rgb <= "111001";
					when "00100000010010101" => rgb <= "111001";
					when "00100000010010110" => rgb <= "111001";
					when "00100000010010111" => rgb <= "111001";
					when "00100000010011000" => rgb <= "111001";
					when "00100000010011001" => rgb <= "101001";
					when "00100000010011010" => rgb <= "101001";
					when "00100000010011011" => rgb <= "111001";
					when "00100000010011100" => rgb <= "111001";
					when "00100000010011101" => rgb <= "101001";
					when "00100000010011110" => rgb <= "111001";
					when "00100000010011111" => rgb <= "101000";
					when "00100000010100000" => rgb <= "101000";
					when "00100000010100001" => rgb <= "101000";
					when "00100000010100010" => rgb <= "101000";
					when "00100000010100011" => rgb <= "101000";
					when "00100000010100100" => rgb <= "101000";
					when "00100000010100101" => rgb <= "101000";
					when "00100000010100110" => rgb <= "101000";
					when "00100000010100111" => rgb <= "101000";
					when "00100000010101000" => rgb <= "101000";
					when "00100000010101001" => rgb <= "101000";
					when "00100000010101010" => rgb <= "101000";
					when "00100000010101011" => rgb <= "101000";
					when "00100000010101100" => rgb <= "101000";
					when "00100000010101101" => rgb <= "101000";
					when "00100000010101110" => rgb <= "101000";
					when "00100000010101111" => rgb <= "101000";
					when "00100000010110000" => rgb <= "101000";
					when "00100000010110001" => rgb <= "101000";
					when "00100000010110010" => rgb <= "101000";
					when "00100000010110011" => rgb <= "101000";
					when "00100000010110100" => rgb <= "101000";
					when "00100000010110101" => rgb <= "101000";
					when "00100000010110110" => rgb <= "101000";
					when "00100000010110111" => rgb <= "101000";
					when "00100000010111000" => rgb <= "101000";
					when "00100000010111001" => rgb <= "101000";
					when "00100000010111010" => rgb <= "101000";
					when "00100000010111011" => rgb <= "101000";
					when "00100000010111100" => rgb <= "101000";
					when "00100000010111101" => rgb <= "101000";
					when "00100000010111110" => rgb <= "101000";
					when "00100000010111111" => rgb <= "101000";
					when "00100000011000000" => rgb <= "100100";
					when "00100000011000001" => rgb <= "000000";
					when "00100000011000010" => rgb <= "000000";
					when "00100000011000011" => rgb <= "000000";
					when "00100000011000100" => rgb <= "000000";
					when "00100000011000101" => rgb <= "000000";
					when "00100000011000110" => rgb <= "000000";
					when "00100000011000111" => rgb <= "000000";
					when "00100000011001000" => rgb <= "000000";
					when "00100000011001001" => rgb <= "000000";
					when "00100000011001010" => rgb <= "000000";
					when "00100000011001011" => rgb <= "000000";
					when "00100000011001100" => rgb <= "000000";
					when "00100000011001101" => rgb <= "000000";
					when "00100000011001110" => rgb <= "000000";
					when "00100000011001111" => rgb <= "000000";
					when "00100000011010000" => rgb <= "000000";
					when "00100000011010001" => rgb <= "000000";
					when "00100000011010010" => rgb <= "000000";
					when "00100000011010011" => rgb <= "000000";
					when "00100000011010100" => rgb <= "000000";
					when "00100000011010101" => rgb <= "000000";
					when "00100000011010110" => rgb <= "000000";
					when "00100000011010111" => rgb <= "000000";
					when "00100000011011000" => rgb <= "000000";
					when "00100000011011001" => rgb <= "000000";
					when "00100000011011010" => rgb <= "000000";
					when "00100000011011011" => rgb <= "000000";
					when "00100000011011100" => rgb <= "000000";
					when "00100000011011101" => rgb <= "000000";
					when "00100000011011110" => rgb <= "000000";
					when "00100000011011111" => rgb <= "000000";
					when "00100000011100000" => rgb <= "000000";
					when "00100000011100001" => rgb <= "000000";
					when "00100000011100010" => rgb <= "000000";
					when "00100000011100011" => rgb <= "000000";
					when "00100000011100100" => rgb <= "000000";
					when "00100000011100101" => rgb <= "000000";
					when "00100000011100110" => rgb <= "000000";
					when "00100000011100111" => rgb <= "000000";
					when "00100000011101000" => rgb <= "000000";
					when "00100000011101001" => rgb <= "000000";
					when "00100000011101010" => rgb <= "000000";
					when "00100000011101011" => rgb <= "000000";
					when "00100000011101100" => rgb <= "000000";
					when "00100000011101101" => rgb <= "000000";
					when "00100000011101110" => rgb <= "000000";
					when "00100000011101111" => rgb <= "000000";
					when "00100000011110000" => rgb <= "000000";
					when "00100000011110001" => rgb <= "000000";
					when "00100000011110010" => rgb <= "000000";
					when "00100000011110011" => rgb <= "000000";
					when "00100000011110100" => rgb <= "000000";
					when "00100000011110101" => rgb <= "000000";
					when "00100000011110110" => rgb <= "000000";
					when "00100000011110111" => rgb <= "000000";
					when "00100000011111000" => rgb <= "000000";
					when "00100000011111001" => rgb <= "000000";
					when "00100000011111010" => rgb <= "000000";
					when "00100000011111011" => rgb <= "000000";
					when "00100000011111100" => rgb <= "000000";
					when "00100000011111101" => rgb <= "000000";
					when "00100000011111110" => rgb <= "000000";
					when "00100000011111111" => rgb <= "000000";
					when "00100000100000000" => rgb <= "000000";
					when "00100000100000001" => rgb <= "000000";
					when "00100000100000010" => rgb <= "000000";
					when "00100000100000011" => rgb <= "000000";
					when "00100000100000100" => rgb <= "000000";
					when "00100000100000101" => rgb <= "000000";
					when "00100000100000110" => rgb <= "000000";
					when "00100000100000111" => rgb <= "000000";
					when "00100000100001000" => rgb <= "000000";
					when "00100000100001001" => rgb <= "000000";
					when "00100000100001010" => rgb <= "000000";
					when "00100000100001011" => rgb <= "000000";
					when "00100000100001100" => rgb <= "000000";
					when "00100000100001101" => rgb <= "000000";
					when "00100000100001110" => rgb <= "000000";
					when "00100000100001111" => rgb <= "000000";
					when "00100000100010000" => rgb <= "000000";
					when "00100000100010001" => rgb <= "000000";
					when "00100000100010010" => rgb <= "000000";
					when "00100000100010011" => rgb <= "000000";
					when "00100000100010100" => rgb <= "000000";
					when "00100000100010101" => rgb <= "000000";
					when "00100000100010110" => rgb <= "000000";
					when "00100000100010111" => rgb <= "000000";
					when "00100000100011000" => rgb <= "000000";
					when "00100000100011001" => rgb <= "000000";
					when "00100000100011010" => rgb <= "000000";
					when "00100000100011011" => rgb <= "000000";
					when "00100000100011100" => rgb <= "000000";
					when "00100000100011101" => rgb <= "000000";
					when "00100000100011110" => rgb <= "000000";
					when "00100000100011111" => rgb <= "000000";
					when "00100000100100000" => rgb <= "000000";
					when "00100000100100001" => rgb <= "000000";
					when "00100000100100010" => rgb <= "000000";
					when "00100000100100011" => rgb <= "000000";
					when "00100000100100100" => rgb <= "000000";
					when "00100000100100101" => rgb <= "000000";
					when "00100000100100110" => rgb <= "000000";
					when "00100000100100111" => rgb <= "000000";
					when "00100000100101000" => rgb <= "000000";
					when "00100000100101001" => rgb <= "000000";
					when "00100000100101010" => rgb <= "000000";
					when "00100000100101011" => rgb <= "000000";
					when "00100000100101100" => rgb <= "000000";
					when "00100000100101101" => rgb <= "000000";
					when "00100000100101110" => rgb <= "000000";
					when "00100000100101111" => rgb <= "000000";
					when "00100000100110000" => rgb <= "000000";
					when "00100000100110001" => rgb <= "000000";
					when "00100000100110010" => rgb <= "000000";
					when "00100000100110011" => rgb <= "000000";
					when "00100000100110100" => rgb <= "000000";
					when "00100000100110101" => rgb <= "000000";
					when "00100000100110110" => rgb <= "000000";
					when "00100000100110111" => rgb <= "000000";
					when "00100000100111000" => rgb <= "000000";
					when "00100000100111001" => rgb <= "000000";
					when "00100000100111010" => rgb <= "000000";
					when "00100000100111011" => rgb <= "000000";
					when "00100000100111100" => rgb <= "000000";
					when "00100000100111101" => rgb <= "000000";
					when "00100000100111110" => rgb <= "000000";
					when "00100000100111111" => rgb <= "000000";
					when "00100001000000000" => rgb <= "000000";
					when "00100001000000001" => rgb <= "000000";
					when "00100001000000010" => rgb <= "000000";
					when "00100001000000011" => rgb <= "000000";
					when "00100001000000100" => rgb <= "000000";
					when "00100001000000101" => rgb <= "000000";
					when "00100001000000110" => rgb <= "000000";
					when "00100001000000111" => rgb <= "000000";
					when "00100001000001000" => rgb <= "000000";
					when "00100001000001001" => rgb <= "000000";
					when "00100001000001010" => rgb <= "000000";
					when "00100001000001011" => rgb <= "000000";
					when "00100001000001100" => rgb <= "000000";
					when "00100001000001101" => rgb <= "000000";
					when "00100001000001110" => rgb <= "000000";
					when "00100001000001111" => rgb <= "000000";
					when "00100001000010000" => rgb <= "000000";
					when "00100001000010001" => rgb <= "000000";
					when "00100001000010010" => rgb <= "000000";
					when "00100001000010011" => rgb <= "000000";
					when "00100001000010100" => rgb <= "000000";
					when "00100001000010101" => rgb <= "000000";
					when "00100001000010110" => rgb <= "000000";
					when "00100001000010111" => rgb <= "000000";
					when "00100001000011000" => rgb <= "000000";
					when "00100001000011001" => rgb <= "000000";
					when "00100001000011010" => rgb <= "000000";
					when "00100001000011011" => rgb <= "000000";
					when "00100001000011100" => rgb <= "000000";
					when "00100001000011101" => rgb <= "000000";
					when "00100001000011110" => rgb <= "000000";
					when "00100001000011111" => rgb <= "000000";
					when "00100001000100000" => rgb <= "000000";
					when "00100001000100001" => rgb <= "000000";
					when "00100001000100010" => rgb <= "000000";
					when "00100001000100011" => rgb <= "000000";
					when "00100001000100100" => rgb <= "000000";
					when "00100001000100101" => rgb <= "000000";
					when "00100001000100110" => rgb <= "000000";
					when "00100001000100111" => rgb <= "000000";
					when "00100001000101000" => rgb <= "000000";
					when "00100001000101001" => rgb <= "000000";
					when "00100001000101010" => rgb <= "000000";
					when "00100001000101011" => rgb <= "000000";
					when "00100001000101100" => rgb <= "000000";
					when "00100001000101101" => rgb <= "000000";
					when "00100001000101110" => rgb <= "000000";
					when "00100001000101111" => rgb <= "000000";
					when "00100001000110000" => rgb <= "000000";
					when "00100001000110001" => rgb <= "000000";
					when "00100001000110010" => rgb <= "000000";
					when "00100001000110011" => rgb <= "000000";
					when "00100001000110100" => rgb <= "000000";
					when "00100001000110101" => rgb <= "000000";
					when "00100001000110110" => rgb <= "000000";
					when "00100001000110111" => rgb <= "000000";
					when "00100001000111000" => rgb <= "000000";
					when "00100001000111001" => rgb <= "000000";
					when "00100001000111010" => rgb <= "000000";
					when "00100001000111011" => rgb <= "000000";
					when "00100001000111100" => rgb <= "000000";
					when "00100001000111101" => rgb <= "000000";
					when "00100001000111110" => rgb <= "000000";
					when "00100001000111111" => rgb <= "000000";
					when "00100001001000000" => rgb <= "000000";
					when "00100001001000001" => rgb <= "000000";
					when "00100001001000010" => rgb <= "000000";
					when "00100001001000011" => rgb <= "000000";
					when "00100001001000100" => rgb <= "000000";
					when "00100001001000101" => rgb <= "000000";
					when "00100001001000110" => rgb <= "000000";
					when "00100001001000111" => rgb <= "000000";
					when "00100001001001000" => rgb <= "000000";
					when "00100001001001001" => rgb <= "000000";
					when "00100001001001010" => rgb <= "000000";
					when "00100001001001011" => rgb <= "000000";
					when "00100001001001100" => rgb <= "000000";
					when "00100001001001101" => rgb <= "000000";
					when "00100001001001110" => rgb <= "000000";
					when "00100001001001111" => rgb <= "000000";
					when "00100001001010000" => rgb <= "000000";
					when "00100001001010001" => rgb <= "000000";
					when "00100001001010010" => rgb <= "000000";
					when "00100001001010011" => rgb <= "000000";
					when "00100001001010100" => rgb <= "000000";
					when "00100001001010101" => rgb <= "000000";
					when "00100001001010110" => rgb <= "000000";
					when "00100001001010111" => rgb <= "000000";
					when "00100001001011000" => rgb <= "000000";
					when "00100001001011001" => rgb <= "000000";
					when "00100001001011010" => rgb <= "000000";
					when "00100001001011011" => rgb <= "000000";
					when "00100001001011100" => rgb <= "000000";
					when "00100001001011101" => rgb <= "000000";
					when "00100001001011110" => rgb <= "000000";
					when "00100001001011111" => rgb <= "000000";
					when "00100001001100000" => rgb <= "000000";
					when "00100001001100001" => rgb <= "000000";
					when "00100001001100010" => rgb <= "000000";
					when "00100001001100011" => rgb <= "000000";
					when "00100001001100100" => rgb <= "000000";
					when "00100001001100101" => rgb <= "000000";
					when "00100001001100110" => rgb <= "000000";
					when "00100001001100111" => rgb <= "000000";
					when "00100001001101000" => rgb <= "000000";
					when "00100001001101001" => rgb <= "000000";
					when "00100001001101010" => rgb <= "000000";
					when "00100001001101011" => rgb <= "000000";
					when "00100001001101100" => rgb <= "000000";
					when "00100001001101101" => rgb <= "000000";
					when "00100001001101110" => rgb <= "000000";
					when "00100001001101111" => rgb <= "000000";
					when "00100001001110000" => rgb <= "000000";
					when "00100001001110001" => rgb <= "000000";
					when "00100001001110010" => rgb <= "000000";
					when "00100001001110011" => rgb <= "000000";
					when "00100001001110100" => rgb <= "000000";
					when "00100001001110101" => rgb <= "000000";
					when "00100001001110110" => rgb <= "000000";
					when "00100001001110111" => rgb <= "000000";
					when "00100001001111000" => rgb <= "000000";
					when "00100001001111001" => rgb <= "000000";
					when "00100001001111010" => rgb <= "000000";
					when "00100001001111011" => rgb <= "000000";
					when "00100001001111100" => rgb <= "000000";
					when "00100001001111101" => rgb <= "101000";
					when "00100001001111110" => rgb <= "101000";
					when "00100001001111111" => rgb <= "101000";
					when "00100001010000000" => rgb <= "101000";
					when "00100001010000001" => rgb <= "101000";
					when "00100001010000010" => rgb <= "101000";
					when "00100001010000011" => rgb <= "101000";
					when "00100001010000100" => rgb <= "101000";
					when "00100001010000101" => rgb <= "101000";
					when "00100001010000110" => rgb <= "101000";
					when "00100001010000111" => rgb <= "101000";
					when "00100001010001000" => rgb <= "101001";
					when "00100001010001001" => rgb <= "111001";
					when "00100001010001010" => rgb <= "101001";
					when "00100001010001011" => rgb <= "101001";
					when "00100001010001100" => rgb <= "111001";
					when "00100001010001101" => rgb <= "111001";
					when "00100001010001110" => rgb <= "111001";
					when "00100001010001111" => rgb <= "101001";
					when "00100001010010000" => rgb <= "101001";
					when "00100001010010001" => rgb <= "101001";
					when "00100001010010010" => rgb <= "101001";
					when "00100001010010011" => rgb <= "111001";
					when "00100001010010100" => rgb <= "111001";
					when "00100001010010101" => rgb <= "111001";
					when "00100001010010110" => rgb <= "111001";
					when "00100001010010111" => rgb <= "111001";
					when "00100001010011000" => rgb <= "111001";
					when "00100001010011001" => rgb <= "101001";
					when "00100001010011010" => rgb <= "101001";
					when "00100001010011011" => rgb <= "111001";
					when "00100001010011100" => rgb <= "111001";
					when "00100001010011101" => rgb <= "101001";
					when "00100001010011110" => rgb <= "111001";
					when "00100001010011111" => rgb <= "101000";
					when "00100001010100000" => rgb <= "101000";
					when "00100001010100001" => rgb <= "101000";
					when "00100001010100010" => rgb <= "101000";
					when "00100001010100011" => rgb <= "101000";
					when "00100001010100100" => rgb <= "101000";
					when "00100001010100101" => rgb <= "101000";
					when "00100001010100110" => rgb <= "101000";
					when "00100001010100111" => rgb <= "101000";
					when "00100001010101000" => rgb <= "101000";
					when "00100001010101001" => rgb <= "101000";
					when "00100001010101010" => rgb <= "101000";
					when "00100001010101011" => rgb <= "101000";
					when "00100001010101100" => rgb <= "101000";
					when "00100001010101101" => rgb <= "101000";
					when "00100001010101110" => rgb <= "101000";
					when "00100001010101111" => rgb <= "101000";
					when "00100001010110000" => rgb <= "101000";
					when "00100001010110001" => rgb <= "101000";
					when "00100001010110010" => rgb <= "101000";
					when "00100001010110011" => rgb <= "101000";
					when "00100001010110100" => rgb <= "101000";
					when "00100001010110101" => rgb <= "101000";
					when "00100001010110110" => rgb <= "101000";
					when "00100001010110111" => rgb <= "101000";
					when "00100001010111000" => rgb <= "101000";
					when "00100001010111001" => rgb <= "101000";
					when "00100001010111010" => rgb <= "101000";
					when "00100001010111011" => rgb <= "101000";
					when "00100001010111100" => rgb <= "101000";
					when "00100001010111101" => rgb <= "101000";
					when "00100001010111110" => rgb <= "101000";
					when "00100001010111111" => rgb <= "101000";
					when "00100001011000000" => rgb <= "100100";
					when "00100001011000001" => rgb <= "000000";
					when "00100001011000010" => rgb <= "000000";
					when "00100001011000011" => rgb <= "000000";
					when "00100001011000100" => rgb <= "000000";
					when "00100001011000101" => rgb <= "000000";
					when "00100001011000110" => rgb <= "000000";
					when "00100001011000111" => rgb <= "000000";
					when "00100001011001000" => rgb <= "000000";
					when "00100001011001001" => rgb <= "000000";
					when "00100001011001010" => rgb <= "000000";
					when "00100001011001011" => rgb <= "000000";
					when "00100001011001100" => rgb <= "000000";
					when "00100001011001101" => rgb <= "000000";
					when "00100001011001110" => rgb <= "000000";
					when "00100001011001111" => rgb <= "000000";
					when "00100001011010000" => rgb <= "000000";
					when "00100001011010001" => rgb <= "000000";
					when "00100001011010010" => rgb <= "000000";
					when "00100001011010011" => rgb <= "000000";
					when "00100001011010100" => rgb <= "000000";
					when "00100001011010101" => rgb <= "000000";
					when "00100001011010110" => rgb <= "000000";
					when "00100001011010111" => rgb <= "000000";
					when "00100001011011000" => rgb <= "000000";
					when "00100001011011001" => rgb <= "000000";
					when "00100001011011010" => rgb <= "000000";
					when "00100001011011011" => rgb <= "000000";
					when "00100001011011100" => rgb <= "000000";
					when "00100001011011101" => rgb <= "000000";
					when "00100001011011110" => rgb <= "000000";
					when "00100001011011111" => rgb <= "000000";
					when "00100001011100000" => rgb <= "000000";
					when "00100001011100001" => rgb <= "000000";
					when "00100001011100010" => rgb <= "000000";
					when "00100001011100011" => rgb <= "000000";
					when "00100001011100100" => rgb <= "000000";
					when "00100001011100101" => rgb <= "000000";
					when "00100001011100110" => rgb <= "000000";
					when "00100001011100111" => rgb <= "000000";
					when "00100001011101000" => rgb <= "000000";
					when "00100001011101001" => rgb <= "000000";
					when "00100001011101010" => rgb <= "000000";
					when "00100001011101011" => rgb <= "000000";
					when "00100001011101100" => rgb <= "000000";
					when "00100001011101101" => rgb <= "000000";
					when "00100001011101110" => rgb <= "000000";
					when "00100001011101111" => rgb <= "000000";
					when "00100001011110000" => rgb <= "000000";
					when "00100001011110001" => rgb <= "000000";
					when "00100001011110010" => rgb <= "000000";
					when "00100001011110011" => rgb <= "000000";
					when "00100001011110100" => rgb <= "000000";
					when "00100001011110101" => rgb <= "000000";
					when "00100001011110110" => rgb <= "000000";
					when "00100001011110111" => rgb <= "000000";
					when "00100001011111000" => rgb <= "000000";
					when "00100001011111001" => rgb <= "000000";
					when "00100001011111010" => rgb <= "000000";
					when "00100001011111011" => rgb <= "000000";
					when "00100001011111100" => rgb <= "000000";
					when "00100001011111101" => rgb <= "000000";
					when "00100001011111110" => rgb <= "000000";
					when "00100001011111111" => rgb <= "000000";
					when "00100001100000000" => rgb <= "000000";
					when "00100001100000001" => rgb <= "000000";
					when "00100001100000010" => rgb <= "000000";
					when "00100001100000011" => rgb <= "000000";
					when "00100001100000100" => rgb <= "000000";
					when "00100001100000101" => rgb <= "000000";
					when "00100001100000110" => rgb <= "000000";
					when "00100001100000111" => rgb <= "000000";
					when "00100001100001000" => rgb <= "000000";
					when "00100001100001001" => rgb <= "000000";
					when "00100001100001010" => rgb <= "000000";
					when "00100001100001011" => rgb <= "000000";
					when "00100001100001100" => rgb <= "000000";
					when "00100001100001101" => rgb <= "000000";
					when "00100001100001110" => rgb <= "000000";
					when "00100001100001111" => rgb <= "000000";
					when "00100001100010000" => rgb <= "000000";
					when "00100001100010001" => rgb <= "000000";
					when "00100001100010010" => rgb <= "000000";
					when "00100001100010011" => rgb <= "000000";
					when "00100001100010100" => rgb <= "000000";
					when "00100001100010101" => rgb <= "000000";
					when "00100001100010110" => rgb <= "000000";
					when "00100001100010111" => rgb <= "000000";
					when "00100001100011000" => rgb <= "000000";
					when "00100001100011001" => rgb <= "000000";
					when "00100001100011010" => rgb <= "000000";
					when "00100001100011011" => rgb <= "000000";
					when "00100001100011100" => rgb <= "000000";
					when "00100001100011101" => rgb <= "000000";
					when "00100001100011110" => rgb <= "000000";
					when "00100001100011111" => rgb <= "000000";
					when "00100001100100000" => rgb <= "000000";
					when "00100001100100001" => rgb <= "000000";
					when "00100001100100010" => rgb <= "000000";
					when "00100001100100011" => rgb <= "000000";
					when "00100001100100100" => rgb <= "000000";
					when "00100001100100101" => rgb <= "000000";
					when "00100001100100110" => rgb <= "000000";
					when "00100001100100111" => rgb <= "000000";
					when "00100001100101000" => rgb <= "000000";
					when "00100001100101001" => rgb <= "000000";
					when "00100001100101010" => rgb <= "000000";
					when "00100001100101011" => rgb <= "000000";
					when "00100001100101100" => rgb <= "000000";
					when "00100001100101101" => rgb <= "000000";
					when "00100001100101110" => rgb <= "000000";
					when "00100001100101111" => rgb <= "000000";
					when "00100001100110000" => rgb <= "000000";
					when "00100001100110001" => rgb <= "000000";
					when "00100001100110010" => rgb <= "000000";
					when "00100001100110011" => rgb <= "000000";
					when "00100001100110100" => rgb <= "000000";
					when "00100001100110101" => rgb <= "000000";
					when "00100001100110110" => rgb <= "000000";
					when "00100001100110111" => rgb <= "000000";
					when "00100001100111000" => rgb <= "000000";
					when "00100001100111001" => rgb <= "000000";
					when "00100001100111010" => rgb <= "000000";
					when "00100001100111011" => rgb <= "000000";
					when "00100001100111100" => rgb <= "000000";
					when "00100001100111101" => rgb <= "000000";
					when "00100001100111110" => rgb <= "000000";
					when "00100001100111111" => rgb <= "000000";
					when "00100010000000000" => rgb <= "000000";
					when "00100010000000001" => rgb <= "000000";
					when "00100010000000010" => rgb <= "000000";
					when "00100010000000011" => rgb <= "000000";
					when "00100010000000100" => rgb <= "000000";
					when "00100010000000101" => rgb <= "000000";
					when "00100010000000110" => rgb <= "000000";
					when "00100010000000111" => rgb <= "000000";
					when "00100010000001000" => rgb <= "000000";
					when "00100010000001001" => rgb <= "000000";
					when "00100010000001010" => rgb <= "000000";
					when "00100010000001011" => rgb <= "000000";
					when "00100010000001100" => rgb <= "000000";
					when "00100010000001101" => rgb <= "000000";
					when "00100010000001110" => rgb <= "000000";
					when "00100010000001111" => rgb <= "000000";
					when "00100010000010000" => rgb <= "000000";
					when "00100010000010001" => rgb <= "000000";
					when "00100010000010010" => rgb <= "000000";
					when "00100010000010011" => rgb <= "000000";
					when "00100010000010100" => rgb <= "000000";
					when "00100010000010101" => rgb <= "000000";
					when "00100010000010110" => rgb <= "000000";
					when "00100010000010111" => rgb <= "000000";
					when "00100010000011000" => rgb <= "000000";
					when "00100010000011001" => rgb <= "000000";
					when "00100010000011010" => rgb <= "000000";
					when "00100010000011011" => rgb <= "000000";
					when "00100010000011100" => rgb <= "000000";
					when "00100010000011101" => rgb <= "000000";
					when "00100010000011110" => rgb <= "000000";
					when "00100010000011111" => rgb <= "000000";
					when "00100010000100000" => rgb <= "000000";
					when "00100010000100001" => rgb <= "000000";
					when "00100010000100010" => rgb <= "000000";
					when "00100010000100011" => rgb <= "000000";
					when "00100010000100100" => rgb <= "000000";
					when "00100010000100101" => rgb <= "000000";
					when "00100010000100110" => rgb <= "000000";
					when "00100010000100111" => rgb <= "000000";
					when "00100010000101000" => rgb <= "000000";
					when "00100010000101001" => rgb <= "000000";
					when "00100010000101010" => rgb <= "000000";
					when "00100010000101011" => rgb <= "000000";
					when "00100010000101100" => rgb <= "000000";
					when "00100010000101101" => rgb <= "000000";
					when "00100010000101110" => rgb <= "000000";
					when "00100010000101111" => rgb <= "000000";
					when "00100010000110000" => rgb <= "000000";
					when "00100010000110001" => rgb <= "000000";
					when "00100010000110010" => rgb <= "000000";
					when "00100010000110011" => rgb <= "000000";
					when "00100010000110100" => rgb <= "000000";
					when "00100010000110101" => rgb <= "000000";
					when "00100010000110110" => rgb <= "000000";
					when "00100010000110111" => rgb <= "000000";
					when "00100010000111000" => rgb <= "000000";
					when "00100010000111001" => rgb <= "000000";
					when "00100010000111010" => rgb <= "000000";
					when "00100010000111011" => rgb <= "000000";
					when "00100010000111100" => rgb <= "000000";
					when "00100010000111101" => rgb <= "000000";
					when "00100010000111110" => rgb <= "000000";
					when "00100010000111111" => rgb <= "000000";
					when "00100010001000000" => rgb <= "000000";
					when "00100010001000001" => rgb <= "000000";
					when "00100010001000010" => rgb <= "000000";
					when "00100010001000011" => rgb <= "000000";
					when "00100010001000100" => rgb <= "000000";
					when "00100010001000101" => rgb <= "000000";
					when "00100010001000110" => rgb <= "000000";
					when "00100010001000111" => rgb <= "000000";
					when "00100010001001000" => rgb <= "000000";
					when "00100010001001001" => rgb <= "000000";
					when "00100010001001010" => rgb <= "000000";
					when "00100010001001011" => rgb <= "000000";
					when "00100010001001100" => rgb <= "000000";
					when "00100010001001101" => rgb <= "000000";
					when "00100010001001110" => rgb <= "000000";
					when "00100010001001111" => rgb <= "000000";
					when "00100010001010000" => rgb <= "000000";
					when "00100010001010001" => rgb <= "000000";
					when "00100010001010010" => rgb <= "000000";
					when "00100010001010011" => rgb <= "000000";
					when "00100010001010100" => rgb <= "000000";
					when "00100010001010101" => rgb <= "000000";
					when "00100010001010110" => rgb <= "000000";
					when "00100010001010111" => rgb <= "000000";
					when "00100010001011000" => rgb <= "000000";
					when "00100010001011001" => rgb <= "000000";
					when "00100010001011010" => rgb <= "000000";
					when "00100010001011011" => rgb <= "000000";
					when "00100010001011100" => rgb <= "000000";
					when "00100010001011101" => rgb <= "000000";
					when "00100010001011110" => rgb <= "000000";
					when "00100010001011111" => rgb <= "000000";
					when "00100010001100000" => rgb <= "000000";
					when "00100010001100001" => rgb <= "000000";
					when "00100010001100010" => rgb <= "000000";
					when "00100010001100011" => rgb <= "000000";
					when "00100010001100100" => rgb <= "000000";
					when "00100010001100101" => rgb <= "000000";
					when "00100010001100110" => rgb <= "000000";
					when "00100010001100111" => rgb <= "000000";
					when "00100010001101000" => rgb <= "000000";
					when "00100010001101001" => rgb <= "000000";
					when "00100010001101010" => rgb <= "000000";
					when "00100010001101011" => rgb <= "000000";
					when "00100010001101100" => rgb <= "000000";
					when "00100010001101101" => rgb <= "000000";
					when "00100010001101110" => rgb <= "000000";
					when "00100010001101111" => rgb <= "000000";
					when "00100010001110000" => rgb <= "000000";
					when "00100010001110001" => rgb <= "000000";
					when "00100010001110010" => rgb <= "000000";
					when "00100010001110011" => rgb <= "000000";
					when "00100010001110100" => rgb <= "000000";
					when "00100010001110101" => rgb <= "000000";
					when "00100010001110110" => rgb <= "000000";
					when "00100010001110111" => rgb <= "000000";
					when "00100010001111000" => rgb <= "000000";
					when "00100010001111001" => rgb <= "000000";
					when "00100010001111010" => rgb <= "000000";
					when "00100010001111011" => rgb <= "000000";
					when "00100010001111100" => rgb <= "000000";
					when "00100010001111101" => rgb <= "101000";
					when "00100010001111110" => rgb <= "101000";
					when "00100010001111111" => rgb <= "101000";
					when "00100010010000000" => rgb <= "101000";
					when "00100010010000001" => rgb <= "101000";
					when "00100010010000010" => rgb <= "101000";
					when "00100010010000011" => rgb <= "101000";
					when "00100010010000100" => rgb <= "101000";
					when "00100010010000101" => rgb <= "101000";
					when "00100010010000110" => rgb <= "101000";
					when "00100010010000111" => rgb <= "101000";
					when "00100010010001000" => rgb <= "101001";
					when "00100010010001001" => rgb <= "111001";
					when "00100010010001010" => rgb <= "101001";
					when "00100010010001011" => rgb <= "101001";
					when "00100010010001100" => rgb <= "111001";
					when "00100010010001101" => rgb <= "111001";
					when "00100010010001110" => rgb <= "111001";
					when "00100010010001111" => rgb <= "101001";
					when "00100010010010000" => rgb <= "111001";
					when "00100010010010001" => rgb <= "111001";
					when "00100010010010010" => rgb <= "111001";
					when "00100010010010011" => rgb <= "111001";
					when "00100010010010100" => rgb <= "111001";
					when "00100010010010101" => rgb <= "111001";
					when "00100010010010110" => rgb <= "111001";
					when "00100010010010111" => rgb <= "111001";
					when "00100010010011000" => rgb <= "111001";
					when "00100010010011001" => rgb <= "101001";
					when "00100010010011010" => rgb <= "101001";
					when "00100010010011011" => rgb <= "111001";
					when "00100010010011100" => rgb <= "111001";
					when "00100010010011101" => rgb <= "101001";
					when "00100010010011110" => rgb <= "111001";
					when "00100010010011111" => rgb <= "101000";
					when "00100010010100000" => rgb <= "101000";
					when "00100010010100001" => rgb <= "101000";
					when "00100010010100010" => rgb <= "101000";
					when "00100010010100011" => rgb <= "101000";
					when "00100010010100100" => rgb <= "101000";
					when "00100010010100101" => rgb <= "101000";
					when "00100010010100110" => rgb <= "101000";
					when "00100010010100111" => rgb <= "101000";
					when "00100010010101000" => rgb <= "101000";
					when "00100010010101001" => rgb <= "101000";
					when "00100010010101010" => rgb <= "101000";
					when "00100010010101011" => rgb <= "101000";
					when "00100010010101100" => rgb <= "101000";
					when "00100010010101101" => rgb <= "101000";
					when "00100010010101110" => rgb <= "101000";
					when "00100010010101111" => rgb <= "101000";
					when "00100010010110000" => rgb <= "101000";
					when "00100010010110001" => rgb <= "101000";
					when "00100010010110010" => rgb <= "101000";
					when "00100010010110011" => rgb <= "101000";
					when "00100010010110100" => rgb <= "101000";
					when "00100010010110101" => rgb <= "101000";
					when "00100010010110110" => rgb <= "101000";
					when "00100010010110111" => rgb <= "101000";
					when "00100010010111000" => rgb <= "101000";
					when "00100010010111001" => rgb <= "101000";
					when "00100010010111010" => rgb <= "101000";
					when "00100010010111011" => rgb <= "101000";
					when "00100010010111100" => rgb <= "101000";
					when "00100010010111101" => rgb <= "101000";
					when "00100010010111110" => rgb <= "101000";
					when "00100010010111111" => rgb <= "101000";
					when "00100010011000000" => rgb <= "100100";
					when "00100010011000001" => rgb <= "000000";
					when "00100010011000010" => rgb <= "000000";
					when "00100010011000011" => rgb <= "000000";
					when "00100010011000100" => rgb <= "000000";
					when "00100010011000101" => rgb <= "000000";
					when "00100010011000110" => rgb <= "000000";
					when "00100010011000111" => rgb <= "000000";
					when "00100010011001000" => rgb <= "000000";
					when "00100010011001001" => rgb <= "000000";
					when "00100010011001010" => rgb <= "000000";
					when "00100010011001011" => rgb <= "000000";
					when "00100010011001100" => rgb <= "000000";
					when "00100010011001101" => rgb <= "000000";
					when "00100010011001110" => rgb <= "000000";
					when "00100010011001111" => rgb <= "000000";
					when "00100010011010000" => rgb <= "000000";
					when "00100010011010001" => rgb <= "000000";
					when "00100010011010010" => rgb <= "000000";
					when "00100010011010011" => rgb <= "000000";
					when "00100010011010100" => rgb <= "000000";
					when "00100010011010101" => rgb <= "000000";
					when "00100010011010110" => rgb <= "000000";
					when "00100010011010111" => rgb <= "000000";
					when "00100010011011000" => rgb <= "000000";
					when "00100010011011001" => rgb <= "000000";
					when "00100010011011010" => rgb <= "000000";
					when "00100010011011011" => rgb <= "000000";
					when "00100010011011100" => rgb <= "000000";
					when "00100010011011101" => rgb <= "000000";
					when "00100010011011110" => rgb <= "000000";
					when "00100010011011111" => rgb <= "000000";
					when "00100010011100000" => rgb <= "000000";
					when "00100010011100001" => rgb <= "000000";
					when "00100010011100010" => rgb <= "000000";
					when "00100010011100011" => rgb <= "000000";
					when "00100010011100100" => rgb <= "000000";
					when "00100010011100101" => rgb <= "000000";
					when "00100010011100110" => rgb <= "000000";
					when "00100010011100111" => rgb <= "000000";
					when "00100010011101000" => rgb <= "000000";
					when "00100010011101001" => rgb <= "000000";
					when "00100010011101010" => rgb <= "000000";
					when "00100010011101011" => rgb <= "000000";
					when "00100010011101100" => rgb <= "000000";
					when "00100010011101101" => rgb <= "000000";
					when "00100010011101110" => rgb <= "000000";
					when "00100010011101111" => rgb <= "000000";
					when "00100010011110000" => rgb <= "000000";
					when "00100010011110001" => rgb <= "000000";
					when "00100010011110010" => rgb <= "000000";
					when "00100010011110011" => rgb <= "000000";
					when "00100010011110100" => rgb <= "000000";
					when "00100010011110101" => rgb <= "000000";
					when "00100010011110110" => rgb <= "000000";
					when "00100010011110111" => rgb <= "000000";
					when "00100010011111000" => rgb <= "000000";
					when "00100010011111001" => rgb <= "000000";
					when "00100010011111010" => rgb <= "000000";
					when "00100010011111011" => rgb <= "000000";
					when "00100010011111100" => rgb <= "000000";
					when "00100010011111101" => rgb <= "000000";
					when "00100010011111110" => rgb <= "000000";
					when "00100010011111111" => rgb <= "000000";
					when "00100010100000000" => rgb <= "000000";
					when "00100010100000001" => rgb <= "000000";
					when "00100010100000010" => rgb <= "000000";
					when "00100010100000011" => rgb <= "000000";
					when "00100010100000100" => rgb <= "000000";
					when "00100010100000101" => rgb <= "000000";
					when "00100010100000110" => rgb <= "000000";
					when "00100010100000111" => rgb <= "000000";
					when "00100010100001000" => rgb <= "000000";
					when "00100010100001001" => rgb <= "000000";
					when "00100010100001010" => rgb <= "000000";
					when "00100010100001011" => rgb <= "000000";
					when "00100010100001100" => rgb <= "000000";
					when "00100010100001101" => rgb <= "000000";
					when "00100010100001110" => rgb <= "000000";
					when "00100010100001111" => rgb <= "000000";
					when "00100010100010000" => rgb <= "000000";
					when "00100010100010001" => rgb <= "000000";
					when "00100010100010010" => rgb <= "000000";
					when "00100010100010011" => rgb <= "000000";
					when "00100010100010100" => rgb <= "000000";
					when "00100010100010101" => rgb <= "000000";
					when "00100010100010110" => rgb <= "000000";
					when "00100010100010111" => rgb <= "000000";
					when "00100010100011000" => rgb <= "000000";
					when "00100010100011001" => rgb <= "000000";
					when "00100010100011010" => rgb <= "000000";
					when "00100010100011011" => rgb <= "000000";
					when "00100010100011100" => rgb <= "000000";
					when "00100010100011101" => rgb <= "000000";
					when "00100010100011110" => rgb <= "000000";
					when "00100010100011111" => rgb <= "000000";
					when "00100010100100000" => rgb <= "000000";
					when "00100010100100001" => rgb <= "000000";
					when "00100010100100010" => rgb <= "000000";
					when "00100010100100011" => rgb <= "000000";
					when "00100010100100100" => rgb <= "000000";
					when "00100010100100101" => rgb <= "000000";
					when "00100010100100110" => rgb <= "000000";
					when "00100010100100111" => rgb <= "000000";
					when "00100010100101000" => rgb <= "000000";
					when "00100010100101001" => rgb <= "000000";
					when "00100010100101010" => rgb <= "000000";
					when "00100010100101011" => rgb <= "000000";
					when "00100010100101100" => rgb <= "000000";
					when "00100010100101101" => rgb <= "000000";
					when "00100010100101110" => rgb <= "000000";
					when "00100010100101111" => rgb <= "000000";
					when "00100010100110000" => rgb <= "000000";
					when "00100010100110001" => rgb <= "000000";
					when "00100010100110010" => rgb <= "000000";
					when "00100010100110011" => rgb <= "000000";
					when "00100010100110100" => rgb <= "000000";
					when "00100010100110101" => rgb <= "000000";
					when "00100010100110110" => rgb <= "000000";
					when "00100010100110111" => rgb <= "000000";
					when "00100010100111000" => rgb <= "000000";
					when "00100010100111001" => rgb <= "000000";
					when "00100010100111010" => rgb <= "000000";
					when "00100010100111011" => rgb <= "000000";
					when "00100010100111100" => rgb <= "000000";
					when "00100010100111101" => rgb <= "000000";
					when "00100010100111110" => rgb <= "000000";
					when "00100010100111111" => rgb <= "000000";
					when "00100011000000000" => rgb <= "000000";
					when "00100011000000001" => rgb <= "000000";
					when "00100011000000010" => rgb <= "000000";
					when "00100011000000011" => rgb <= "000000";
					when "00100011000000100" => rgb <= "000000";
					when "00100011000000101" => rgb <= "000000";
					when "00100011000000110" => rgb <= "000000";
					when "00100011000000111" => rgb <= "000000";
					when "00100011000001000" => rgb <= "000000";
					when "00100011000001001" => rgb <= "000000";
					when "00100011000001010" => rgb <= "000000";
					when "00100011000001011" => rgb <= "000000";
					when "00100011000001100" => rgb <= "000000";
					when "00100011000001101" => rgb <= "000000";
					when "00100011000001110" => rgb <= "000000";
					when "00100011000001111" => rgb <= "000000";
					when "00100011000010000" => rgb <= "000000";
					when "00100011000010001" => rgb <= "000000";
					when "00100011000010010" => rgb <= "000000";
					when "00100011000010011" => rgb <= "000000";
					when "00100011000010100" => rgb <= "000000";
					when "00100011000010101" => rgb <= "000000";
					when "00100011000010110" => rgb <= "000000";
					when "00100011000010111" => rgb <= "000000";
					when "00100011000011000" => rgb <= "000000";
					when "00100011000011001" => rgb <= "000000";
					when "00100011000011010" => rgb <= "000000";
					when "00100011000011011" => rgb <= "000000";
					when "00100011000011100" => rgb <= "000000";
					when "00100011000011101" => rgb <= "000000";
					when "00100011000011110" => rgb <= "000000";
					when "00100011000011111" => rgb <= "000000";
					when "00100011000100000" => rgb <= "000000";
					when "00100011000100001" => rgb <= "000000";
					when "00100011000100010" => rgb <= "000000";
					when "00100011000100011" => rgb <= "000000";
					when "00100011000100100" => rgb <= "000000";
					when "00100011000100101" => rgb <= "000000";
					when "00100011000100110" => rgb <= "000000";
					when "00100011000100111" => rgb <= "000000";
					when "00100011000101000" => rgb <= "000000";
					when "00100011000101001" => rgb <= "000000";
					when "00100011000101010" => rgb <= "000000";
					when "00100011000101011" => rgb <= "000000";
					when "00100011000101100" => rgb <= "000000";
					when "00100011000101101" => rgb <= "000000";
					when "00100011000101110" => rgb <= "000000";
					when "00100011000101111" => rgb <= "000000";
					when "00100011000110000" => rgb <= "000000";
					when "00100011000110001" => rgb <= "000000";
					when "00100011000110010" => rgb <= "000000";
					when "00100011000110011" => rgb <= "000000";
					when "00100011000110100" => rgb <= "000000";
					when "00100011000110101" => rgb <= "000000";
					when "00100011000110110" => rgb <= "000000";
					when "00100011000110111" => rgb <= "000000";
					when "00100011000111000" => rgb <= "000000";
					when "00100011000111001" => rgb <= "000000";
					when "00100011000111010" => rgb <= "000000";
					when "00100011000111011" => rgb <= "000000";
					when "00100011000111100" => rgb <= "000000";
					when "00100011000111101" => rgb <= "000000";
					when "00100011000111110" => rgb <= "000000";
					when "00100011000111111" => rgb <= "000000";
					when "00100011001000000" => rgb <= "000000";
					when "00100011001000001" => rgb <= "000000";
					when "00100011001000010" => rgb <= "000000";
					when "00100011001000011" => rgb <= "000000";
					when "00100011001000100" => rgb <= "000000";
					when "00100011001000101" => rgb <= "000000";
					when "00100011001000110" => rgb <= "000000";
					when "00100011001000111" => rgb <= "000000";
					when "00100011001001000" => rgb <= "000000";
					when "00100011001001001" => rgb <= "000000";
					when "00100011001001010" => rgb <= "000000";
					when "00100011001001011" => rgb <= "000000";
					when "00100011001001100" => rgb <= "000000";
					when "00100011001001101" => rgb <= "000000";
					when "00100011001001110" => rgb <= "000000";
					when "00100011001001111" => rgb <= "000000";
					when "00100011001010000" => rgb <= "000000";
					when "00100011001010001" => rgb <= "000000";
					when "00100011001010010" => rgb <= "000000";
					when "00100011001010011" => rgb <= "000000";
					when "00100011001010100" => rgb <= "000000";
					when "00100011001010101" => rgb <= "000000";
					when "00100011001010110" => rgb <= "000000";
					when "00100011001010111" => rgb <= "000000";
					when "00100011001011000" => rgb <= "000000";
					when "00100011001011001" => rgb <= "000000";
					when "00100011001011010" => rgb <= "000000";
					when "00100011001011011" => rgb <= "000000";
					when "00100011001011100" => rgb <= "000000";
					when "00100011001011101" => rgb <= "000000";
					when "00100011001011110" => rgb <= "000000";
					when "00100011001011111" => rgb <= "000000";
					when "00100011001100000" => rgb <= "000000";
					when "00100011001100001" => rgb <= "000000";
					when "00100011001100010" => rgb <= "000000";
					when "00100011001100011" => rgb <= "000000";
					when "00100011001100100" => rgb <= "000000";
					when "00100011001100101" => rgb <= "000000";
					when "00100011001100110" => rgb <= "000000";
					when "00100011001100111" => rgb <= "000000";
					when "00100011001101000" => rgb <= "000000";
					when "00100011001101001" => rgb <= "000000";
					when "00100011001101010" => rgb <= "000000";
					when "00100011001101011" => rgb <= "000000";
					when "00100011001101100" => rgb <= "000000";
					when "00100011001101101" => rgb <= "000000";
					when "00100011001101110" => rgb <= "000000";
					when "00100011001101111" => rgb <= "000000";
					when "00100011001110000" => rgb <= "000000";
					when "00100011001110001" => rgb <= "000000";
					when "00100011001110010" => rgb <= "000000";
					when "00100011001110011" => rgb <= "000000";
					when "00100011001110100" => rgb <= "000000";
					when "00100011001110101" => rgb <= "000000";
					when "00100011001110110" => rgb <= "000000";
					when "00100011001110111" => rgb <= "000000";
					when "00100011001111000" => rgb <= "000000";
					when "00100011001111001" => rgb <= "000000";
					when "00100011001111010" => rgb <= "000000";
					when "00100011001111011" => rgb <= "000000";
					when "00100011001111100" => rgb <= "000000";
					when "00100011001111101" => rgb <= "101000";
					when "00100011001111110" => rgb <= "101000";
					when "00100011001111111" => rgb <= "101000";
					when "00100011010000000" => rgb <= "101000";
					when "00100011010000001" => rgb <= "101000";
					when "00100011010000010" => rgb <= "101000";
					when "00100011010000011" => rgb <= "101000";
					when "00100011010000100" => rgb <= "101000";
					when "00100011010000101" => rgb <= "101000";
					when "00100011010000110" => rgb <= "101000";
					when "00100011010000111" => rgb <= "101000";
					when "00100011010001000" => rgb <= "101001";
					when "00100011010001001" => rgb <= "111001";
					when "00100011010001010" => rgb <= "101001";
					when "00100011010001011" => rgb <= "101001";
					when "00100011010001100" => rgb <= "111001";
					when "00100011010001101" => rgb <= "111001";
					when "00100011010001110" => rgb <= "111001";
					when "00100011010001111" => rgb <= "101001";
					when "00100011010010000" => rgb <= "111001";
					when "00100011010010001" => rgb <= "111001";
					when "00100011010010010" => rgb <= "111001";
					when "00100011010010011" => rgb <= "111001";
					when "00100011010010100" => rgb <= "111001";
					when "00100011010010101" => rgb <= "111001";
					when "00100011010010110" => rgb <= "111001";
					when "00100011010010111" => rgb <= "111001";
					when "00100011010011000" => rgb <= "111001";
					when "00100011010011001" => rgb <= "101001";
					when "00100011010011010" => rgb <= "111001";
					when "00100011010011011" => rgb <= "111001";
					when "00100011010011100" => rgb <= "111001";
					when "00100011010011101" => rgb <= "101001";
					when "00100011010011110" => rgb <= "111001";
					when "00100011010011111" => rgb <= "101000";
					when "00100011010100000" => rgb <= "101000";
					when "00100011010100001" => rgb <= "101000";
					when "00100011010100010" => rgb <= "101000";
					when "00100011010100011" => rgb <= "101000";
					when "00100011010100100" => rgb <= "101000";
					when "00100011010100101" => rgb <= "101000";
					when "00100011010100110" => rgb <= "101000";
					when "00100011010100111" => rgb <= "101000";
					when "00100011010101000" => rgb <= "101000";
					when "00100011010101001" => rgb <= "101000";
					when "00100011010101010" => rgb <= "101000";
					when "00100011010101011" => rgb <= "101000";
					when "00100011010101100" => rgb <= "101000";
					when "00100011010101101" => rgb <= "101000";
					when "00100011010101110" => rgb <= "101000";
					when "00100011010101111" => rgb <= "101000";
					when "00100011010110000" => rgb <= "101000";
					when "00100011010110001" => rgb <= "101000";
					when "00100011010110010" => rgb <= "101000";
					when "00100011010110011" => rgb <= "101000";
					when "00100011010110100" => rgb <= "101000";
					when "00100011010110101" => rgb <= "101000";
					when "00100011010110110" => rgb <= "101000";
					when "00100011010110111" => rgb <= "101000";
					when "00100011010111000" => rgb <= "101000";
					when "00100011010111001" => rgb <= "101000";
					when "00100011010111010" => rgb <= "101000";
					when "00100011010111011" => rgb <= "101000";
					when "00100011010111100" => rgb <= "101000";
					when "00100011010111101" => rgb <= "101000";
					when "00100011010111110" => rgb <= "101000";
					when "00100011010111111" => rgb <= "101000";
					when "00100011011000000" => rgb <= "100100";
					when "00100011011000001" => rgb <= "000000";
					when "00100011011000010" => rgb <= "000000";
					when "00100011011000011" => rgb <= "000000";
					when "00100011011000100" => rgb <= "000000";
					when "00100011011000101" => rgb <= "000000";
					when "00100011011000110" => rgb <= "000000";
					when "00100011011000111" => rgb <= "000000";
					when "00100011011001000" => rgb <= "000000";
					when "00100011011001001" => rgb <= "000000";
					when "00100011011001010" => rgb <= "000000";
					when "00100011011001011" => rgb <= "000000";
					when "00100011011001100" => rgb <= "000000";
					when "00100011011001101" => rgb <= "000000";
					when "00100011011001110" => rgb <= "000000";
					when "00100011011001111" => rgb <= "000000";
					when "00100011011010000" => rgb <= "000000";
					when "00100011011010001" => rgb <= "000000";
					when "00100011011010010" => rgb <= "000000";
					when "00100011011010011" => rgb <= "000000";
					when "00100011011010100" => rgb <= "000000";
					when "00100011011010101" => rgb <= "000000";
					when "00100011011010110" => rgb <= "000000";
					when "00100011011010111" => rgb <= "000000";
					when "00100011011011000" => rgb <= "000000";
					when "00100011011011001" => rgb <= "000000";
					when "00100011011011010" => rgb <= "000000";
					when "00100011011011011" => rgb <= "000000";
					when "00100011011011100" => rgb <= "000000";
					when "00100011011011101" => rgb <= "000000";
					when "00100011011011110" => rgb <= "000000";
					when "00100011011011111" => rgb <= "000000";
					when "00100011011100000" => rgb <= "000000";
					when "00100011011100001" => rgb <= "000000";
					when "00100011011100010" => rgb <= "000000";
					when "00100011011100011" => rgb <= "000000";
					when "00100011011100100" => rgb <= "000000";
					when "00100011011100101" => rgb <= "000000";
					when "00100011011100110" => rgb <= "000000";
					when "00100011011100111" => rgb <= "000000";
					when "00100011011101000" => rgb <= "000000";
					when "00100011011101001" => rgb <= "000000";
					when "00100011011101010" => rgb <= "000000";
					when "00100011011101011" => rgb <= "000000";
					when "00100011011101100" => rgb <= "000000";
					when "00100011011101101" => rgb <= "000000";
					when "00100011011101110" => rgb <= "000000";
					when "00100011011101111" => rgb <= "000000";
					when "00100011011110000" => rgb <= "000000";
					when "00100011011110001" => rgb <= "000000";
					when "00100011011110010" => rgb <= "000000";
					when "00100011011110011" => rgb <= "000000";
					when "00100011011110100" => rgb <= "000000";
					when "00100011011110101" => rgb <= "000000";
					when "00100011011110110" => rgb <= "000000";
					when "00100011011110111" => rgb <= "000000";
					when "00100011011111000" => rgb <= "000000";
					when "00100011011111001" => rgb <= "000000";
					when "00100011011111010" => rgb <= "000000";
					when "00100011011111011" => rgb <= "000000";
					when "00100011011111100" => rgb <= "000000";
					when "00100011011111101" => rgb <= "000000";
					when "00100011011111110" => rgb <= "000000";
					when "00100011011111111" => rgb <= "000000";
					when "00100011100000000" => rgb <= "000000";
					when "00100011100000001" => rgb <= "000000";
					when "00100011100000010" => rgb <= "000000";
					when "00100011100000011" => rgb <= "000000";
					when "00100011100000100" => rgb <= "000000";
					when "00100011100000101" => rgb <= "000000";
					when "00100011100000110" => rgb <= "000000";
					when "00100011100000111" => rgb <= "000000";
					when "00100011100001000" => rgb <= "000000";
					when "00100011100001001" => rgb <= "000000";
					when "00100011100001010" => rgb <= "000000";
					when "00100011100001011" => rgb <= "000000";
					when "00100011100001100" => rgb <= "000000";
					when "00100011100001101" => rgb <= "000000";
					when "00100011100001110" => rgb <= "000000";
					when "00100011100001111" => rgb <= "000000";
					when "00100011100010000" => rgb <= "000000";
					when "00100011100010001" => rgb <= "000000";
					when "00100011100010010" => rgb <= "000000";
					when "00100011100010011" => rgb <= "000000";
					when "00100011100010100" => rgb <= "000000";
					when "00100011100010101" => rgb <= "000000";
					when "00100011100010110" => rgb <= "000000";
					when "00100011100010111" => rgb <= "000000";
					when "00100011100011000" => rgb <= "000000";
					when "00100011100011001" => rgb <= "000000";
					when "00100011100011010" => rgb <= "000000";
					when "00100011100011011" => rgb <= "000000";
					when "00100011100011100" => rgb <= "000000";
					when "00100011100011101" => rgb <= "000000";
					when "00100011100011110" => rgb <= "000000";
					when "00100011100011111" => rgb <= "000000";
					when "00100011100100000" => rgb <= "000000";
					when "00100011100100001" => rgb <= "000000";
					when "00100011100100010" => rgb <= "000000";
					when "00100011100100011" => rgb <= "000000";
					when "00100011100100100" => rgb <= "000000";
					when "00100011100100101" => rgb <= "000000";
					when "00100011100100110" => rgb <= "000000";
					when "00100011100100111" => rgb <= "000000";
					when "00100011100101000" => rgb <= "000000";
					when "00100011100101001" => rgb <= "000000";
					when "00100011100101010" => rgb <= "000000";
					when "00100011100101011" => rgb <= "000000";
					when "00100011100101100" => rgb <= "000000";
					when "00100011100101101" => rgb <= "000000";
					when "00100011100101110" => rgb <= "000000";
					when "00100011100101111" => rgb <= "000000";
					when "00100011100110000" => rgb <= "000000";
					when "00100011100110001" => rgb <= "000000";
					when "00100011100110010" => rgb <= "000000";
					when "00100011100110011" => rgb <= "000000";
					when "00100011100110100" => rgb <= "000000";
					when "00100011100110101" => rgb <= "000000";
					when "00100011100110110" => rgb <= "000000";
					when "00100011100110111" => rgb <= "000000";
					when "00100011100111000" => rgb <= "000000";
					when "00100011100111001" => rgb <= "000000";
					when "00100011100111010" => rgb <= "000000";
					when "00100011100111011" => rgb <= "000000";
					when "00100011100111100" => rgb <= "000000";
					when "00100011100111101" => rgb <= "000000";
					when "00100011100111110" => rgb <= "000000";
					when "00100011100111111" => rgb <= "000000";
					when "00100100000000000" => rgb <= "000000";
					when "00100100000000001" => rgb <= "000000";
					when "00100100000000010" => rgb <= "000000";
					when "00100100000000011" => rgb <= "000000";
					when "00100100000000100" => rgb <= "000000";
					when "00100100000000101" => rgb <= "000000";
					when "00100100000000110" => rgb <= "000000";
					when "00100100000000111" => rgb <= "000000";
					when "00100100000001000" => rgb <= "000000";
					when "00100100000001001" => rgb <= "000000";
					when "00100100000001010" => rgb <= "000000";
					when "00100100000001011" => rgb <= "000000";
					when "00100100000001100" => rgb <= "000000";
					when "00100100000001101" => rgb <= "000000";
					when "00100100000001110" => rgb <= "000000";
					when "00100100000001111" => rgb <= "000000";
					when "00100100000010000" => rgb <= "000000";
					when "00100100000010001" => rgb <= "000000";
					when "00100100000010010" => rgb <= "000000";
					when "00100100000010011" => rgb <= "000000";
					when "00100100000010100" => rgb <= "000000";
					when "00100100000010101" => rgb <= "000000";
					when "00100100000010110" => rgb <= "000000";
					when "00100100000010111" => rgb <= "000000";
					when "00100100000011000" => rgb <= "000000";
					when "00100100000011001" => rgb <= "000000";
					when "00100100000011010" => rgb <= "000000";
					when "00100100000011011" => rgb <= "000000";
					when "00100100000011100" => rgb <= "000000";
					when "00100100000011101" => rgb <= "000000";
					when "00100100000011110" => rgb <= "000000";
					when "00100100000011111" => rgb <= "000000";
					when "00100100000100000" => rgb <= "000000";
					when "00100100000100001" => rgb <= "000000";
					when "00100100000100010" => rgb <= "000000";
					when "00100100000100011" => rgb <= "000000";
					when "00100100000100100" => rgb <= "000000";
					when "00100100000100101" => rgb <= "000000";
					when "00100100000100110" => rgb <= "000000";
					when "00100100000100111" => rgb <= "000000";
					when "00100100000101000" => rgb <= "000000";
					when "00100100000101001" => rgb <= "000000";
					when "00100100000101010" => rgb <= "000000";
					when "00100100000101011" => rgb <= "000000";
					when "00100100000101100" => rgb <= "000000";
					when "00100100000101101" => rgb <= "000000";
					when "00100100000101110" => rgb <= "000000";
					when "00100100000101111" => rgb <= "000000";
					when "00100100000110000" => rgb <= "000000";
					when "00100100000110001" => rgb <= "000000";
					when "00100100000110010" => rgb <= "000000";
					when "00100100000110011" => rgb <= "000000";
					when "00100100000110100" => rgb <= "000000";
					when "00100100000110101" => rgb <= "000000";
					when "00100100000110110" => rgb <= "000000";
					when "00100100000110111" => rgb <= "000000";
					when "00100100000111000" => rgb <= "000000";
					when "00100100000111001" => rgb <= "000000";
					when "00100100000111010" => rgb <= "000000";
					when "00100100000111011" => rgb <= "000000";
					when "00100100000111100" => rgb <= "000000";
					when "00100100000111101" => rgb <= "000000";
					when "00100100000111110" => rgb <= "000000";
					when "00100100000111111" => rgb <= "000000";
					when "00100100001000000" => rgb <= "000000";
					when "00100100001000001" => rgb <= "000000";
					when "00100100001000010" => rgb <= "000000";
					when "00100100001000011" => rgb <= "000000";
					when "00100100001000100" => rgb <= "000000";
					when "00100100001000101" => rgb <= "000000";
					when "00100100001000110" => rgb <= "000000";
					when "00100100001000111" => rgb <= "000000";
					when "00100100001001000" => rgb <= "000000";
					when "00100100001001001" => rgb <= "000000";
					when "00100100001001010" => rgb <= "000000";
					when "00100100001001011" => rgb <= "000000";
					when "00100100001001100" => rgb <= "000000";
					when "00100100001001101" => rgb <= "000000";
					when "00100100001001110" => rgb <= "000000";
					when "00100100001001111" => rgb <= "000000";
					when "00100100001010000" => rgb <= "000000";
					when "00100100001010001" => rgb <= "000000";
					when "00100100001010010" => rgb <= "000000";
					when "00100100001010011" => rgb <= "000000";
					when "00100100001010100" => rgb <= "000000";
					when "00100100001010101" => rgb <= "000000";
					when "00100100001010110" => rgb <= "000000";
					when "00100100001010111" => rgb <= "000000";
					when "00100100001011000" => rgb <= "000000";
					when "00100100001011001" => rgb <= "000000";
					when "00100100001011010" => rgb <= "000000";
					when "00100100001011011" => rgb <= "000000";
					when "00100100001011100" => rgb <= "000000";
					when "00100100001011101" => rgb <= "000000";
					when "00100100001011110" => rgb <= "000000";
					when "00100100001011111" => rgb <= "000000";
					when "00100100001100000" => rgb <= "000000";
					when "00100100001100001" => rgb <= "000000";
					when "00100100001100010" => rgb <= "000000";
					when "00100100001100011" => rgb <= "000000";
					when "00100100001100100" => rgb <= "000000";
					when "00100100001100101" => rgb <= "000000";
					when "00100100001100110" => rgb <= "000000";
					when "00100100001100111" => rgb <= "000000";
					when "00100100001101000" => rgb <= "000000";
					when "00100100001101001" => rgb <= "000000";
					when "00100100001101010" => rgb <= "000000";
					when "00100100001101011" => rgb <= "000000";
					when "00100100001101100" => rgb <= "000000";
					when "00100100001101101" => rgb <= "000000";
					when "00100100001101110" => rgb <= "000000";
					when "00100100001101111" => rgb <= "000000";
					when "00100100001110000" => rgb <= "000000";
					when "00100100001110001" => rgb <= "000000";
					when "00100100001110010" => rgb <= "000000";
					when "00100100001110011" => rgb <= "000000";
					when "00100100001110100" => rgb <= "000000";
					when "00100100001110101" => rgb <= "000000";
					when "00100100001110110" => rgb <= "000000";
					when "00100100001110111" => rgb <= "000000";
					when "00100100001111000" => rgb <= "000000";
					when "00100100001111001" => rgb <= "000000";
					when "00100100001111010" => rgb <= "000000";
					when "00100100001111011" => rgb <= "000000";
					when "00100100001111100" => rgb <= "000000";
					when "00100100001111101" => rgb <= "101000";
					when "00100100001111110" => rgb <= "101000";
					when "00100100001111111" => rgb <= "101000";
					when "00100100010000000" => rgb <= "101000";
					when "00100100010000001" => rgb <= "101000";
					when "00100100010000010" => rgb <= "101000";
					when "00100100010000011" => rgb <= "101000";
					when "00100100010000100" => rgb <= "101000";
					when "00100100010000101" => rgb <= "101000";
					when "00100100010000110" => rgb <= "101000";
					when "00100100010000111" => rgb <= "101000";
					when "00100100010001000" => rgb <= "101001";
					when "00100100010001001" => rgb <= "111001";
					when "00100100010001010" => rgb <= "101001";
					when "00100100010001011" => rgb <= "101001";
					when "00100100010001100" => rgb <= "111001";
					when "00100100010001101" => rgb <= "111001";
					when "00100100010001110" => rgb <= "111001";
					when "00100100010001111" => rgb <= "101001";
					when "00100100010010000" => rgb <= "101001";
					when "00100100010010001" => rgb <= "101001";
					when "00100100010010010" => rgb <= "101001";
					when "00100100010010011" => rgb <= "101001";
					when "00100100010010100" => rgb <= "101001";
					when "00100100010010101" => rgb <= "101001";
					when "00100100010010110" => rgb <= "101001";
					when "00100100010010111" => rgb <= "101001";
					when "00100100010011000" => rgb <= "111001";
					when "00100100010011001" => rgb <= "101001";
					when "00100100010011010" => rgb <= "101001";
					when "00100100010011011" => rgb <= "111001";
					when "00100100010011100" => rgb <= "111001";
					when "00100100010011101" => rgb <= "101001";
					when "00100100010011110" => rgb <= "101001";
					when "00100100010011111" => rgb <= "101000";
					when "00100100010100000" => rgb <= "101000";
					when "00100100010100001" => rgb <= "101000";
					when "00100100010100010" => rgb <= "101000";
					when "00100100010100011" => rgb <= "101000";
					when "00100100010100100" => rgb <= "101000";
					when "00100100010100101" => rgb <= "101000";
					when "00100100010100110" => rgb <= "101000";
					when "00100100010100111" => rgb <= "101000";
					when "00100100010101000" => rgb <= "101000";
					when "00100100010101001" => rgb <= "101000";
					when "00100100010101010" => rgb <= "101000";
					when "00100100010101011" => rgb <= "101000";
					when "00100100010101100" => rgb <= "101000";
					when "00100100010101101" => rgb <= "101000";
					when "00100100010101110" => rgb <= "101000";
					when "00100100010101111" => rgb <= "101000";
					when "00100100010110000" => rgb <= "101000";
					when "00100100010110001" => rgb <= "101000";
					when "00100100010110010" => rgb <= "101000";
					when "00100100010110011" => rgb <= "101000";
					when "00100100010110100" => rgb <= "101000";
					when "00100100010110101" => rgb <= "101000";
					when "00100100010110110" => rgb <= "101000";
					when "00100100010110111" => rgb <= "101000";
					when "00100100010111000" => rgb <= "101000";
					when "00100100010111001" => rgb <= "101000";
					when "00100100010111010" => rgb <= "101000";
					when "00100100010111011" => rgb <= "101000";
					when "00100100010111100" => rgb <= "101000";
					when "00100100010111101" => rgb <= "101000";
					when "00100100010111110" => rgb <= "101000";
					when "00100100010111111" => rgb <= "101000";
					when "00100100011000000" => rgb <= "100100";
					when "00100100011000001" => rgb <= "000000";
					when "00100100011000010" => rgb <= "000000";
					when "00100100011000011" => rgb <= "000000";
					when "00100100011000100" => rgb <= "000000";
					when "00100100011000101" => rgb <= "000000";
					when "00100100011000110" => rgb <= "000000";
					when "00100100011000111" => rgb <= "000000";
					when "00100100011001000" => rgb <= "000000";
					when "00100100011001001" => rgb <= "000000";
					when "00100100011001010" => rgb <= "000000";
					when "00100100011001011" => rgb <= "000000";
					when "00100100011001100" => rgb <= "000000";
					when "00100100011001101" => rgb <= "000000";
					when "00100100011001110" => rgb <= "000000";
					when "00100100011001111" => rgb <= "000000";
					when "00100100011010000" => rgb <= "000000";
					when "00100100011010001" => rgb <= "000000";
					when "00100100011010010" => rgb <= "000000";
					when "00100100011010011" => rgb <= "000000";
					when "00100100011010100" => rgb <= "000000";
					when "00100100011010101" => rgb <= "000000";
					when "00100100011010110" => rgb <= "000000";
					when "00100100011010111" => rgb <= "000000";
					when "00100100011011000" => rgb <= "000000";
					when "00100100011011001" => rgb <= "000000";
					when "00100100011011010" => rgb <= "000000";
					when "00100100011011011" => rgb <= "000000";
					when "00100100011011100" => rgb <= "000000";
					when "00100100011011101" => rgb <= "000000";
					when "00100100011011110" => rgb <= "000000";
					when "00100100011011111" => rgb <= "000000";
					when "00100100011100000" => rgb <= "000000";
					when "00100100011100001" => rgb <= "000000";
					when "00100100011100010" => rgb <= "000000";
					when "00100100011100011" => rgb <= "000000";
					when "00100100011100100" => rgb <= "000000";
					when "00100100011100101" => rgb <= "000000";
					when "00100100011100110" => rgb <= "000000";
					when "00100100011100111" => rgb <= "000000";
					when "00100100011101000" => rgb <= "000000";
					when "00100100011101001" => rgb <= "000000";
					when "00100100011101010" => rgb <= "000000";
					when "00100100011101011" => rgb <= "000000";
					when "00100100011101100" => rgb <= "000000";
					when "00100100011101101" => rgb <= "000000";
					when "00100100011101110" => rgb <= "000000";
					when "00100100011101111" => rgb <= "000000";
					when "00100100011110000" => rgb <= "000000";
					when "00100100011110001" => rgb <= "000000";
					when "00100100011110010" => rgb <= "000000";
					when "00100100011110011" => rgb <= "000000";
					when "00100100011110100" => rgb <= "000000";
					when "00100100011110101" => rgb <= "000000";
					when "00100100011110110" => rgb <= "000000";
					when "00100100011110111" => rgb <= "000000";
					when "00100100011111000" => rgb <= "000000";
					when "00100100011111001" => rgb <= "000000";
					when "00100100011111010" => rgb <= "000000";
					when "00100100011111011" => rgb <= "000000";
					when "00100100011111100" => rgb <= "000000";
					when "00100100011111101" => rgb <= "000000";
					when "00100100011111110" => rgb <= "000000";
					when "00100100011111111" => rgb <= "000000";
					when "00100100100000000" => rgb <= "000000";
					when "00100100100000001" => rgb <= "000000";
					when "00100100100000010" => rgb <= "000000";
					when "00100100100000011" => rgb <= "000000";
					when "00100100100000100" => rgb <= "000000";
					when "00100100100000101" => rgb <= "000000";
					when "00100100100000110" => rgb <= "000000";
					when "00100100100000111" => rgb <= "000000";
					when "00100100100001000" => rgb <= "000000";
					when "00100100100001001" => rgb <= "000000";
					when "00100100100001010" => rgb <= "000000";
					when "00100100100001011" => rgb <= "000000";
					when "00100100100001100" => rgb <= "000000";
					when "00100100100001101" => rgb <= "000000";
					when "00100100100001110" => rgb <= "000000";
					when "00100100100001111" => rgb <= "000000";
					when "00100100100010000" => rgb <= "000000";
					when "00100100100010001" => rgb <= "000000";
					when "00100100100010010" => rgb <= "000000";
					when "00100100100010011" => rgb <= "000000";
					when "00100100100010100" => rgb <= "000000";
					when "00100100100010101" => rgb <= "000000";
					when "00100100100010110" => rgb <= "000000";
					when "00100100100010111" => rgb <= "000000";
					when "00100100100011000" => rgb <= "000000";
					when "00100100100011001" => rgb <= "000000";
					when "00100100100011010" => rgb <= "000000";
					when "00100100100011011" => rgb <= "000000";
					when "00100100100011100" => rgb <= "000000";
					when "00100100100011101" => rgb <= "000000";
					when "00100100100011110" => rgb <= "000000";
					when "00100100100011111" => rgb <= "000000";
					when "00100100100100000" => rgb <= "000000";
					when "00100100100100001" => rgb <= "000000";
					when "00100100100100010" => rgb <= "000000";
					when "00100100100100011" => rgb <= "000000";
					when "00100100100100100" => rgb <= "000000";
					when "00100100100100101" => rgb <= "000000";
					when "00100100100100110" => rgb <= "000000";
					when "00100100100100111" => rgb <= "000000";
					when "00100100100101000" => rgb <= "000000";
					when "00100100100101001" => rgb <= "000000";
					when "00100100100101010" => rgb <= "000000";
					when "00100100100101011" => rgb <= "000000";
					when "00100100100101100" => rgb <= "000000";
					when "00100100100101101" => rgb <= "000000";
					when "00100100100101110" => rgb <= "000000";
					when "00100100100101111" => rgb <= "000000";
					when "00100100100110000" => rgb <= "000000";
					when "00100100100110001" => rgb <= "000000";
					when "00100100100110010" => rgb <= "000000";
					when "00100100100110011" => rgb <= "000000";
					when "00100100100110100" => rgb <= "000000";
					when "00100100100110101" => rgb <= "000000";
					when "00100100100110110" => rgb <= "000000";
					when "00100100100110111" => rgb <= "000000";
					when "00100100100111000" => rgb <= "000000";
					when "00100100100111001" => rgb <= "000000";
					when "00100100100111010" => rgb <= "000000";
					when "00100100100111011" => rgb <= "000000";
					when "00100100100111100" => rgb <= "000000";
					when "00100100100111101" => rgb <= "000000";
					when "00100100100111110" => rgb <= "000000";
					when "00100100100111111" => rgb <= "000000";
					when "00100101000000000" => rgb <= "000000";
					when "00100101000000001" => rgb <= "000000";
					when "00100101000000010" => rgb <= "000000";
					when "00100101000000011" => rgb <= "000000";
					when "00100101000000100" => rgb <= "000000";
					when "00100101000000101" => rgb <= "000000";
					when "00100101000000110" => rgb <= "000000";
					when "00100101000000111" => rgb <= "000000";
					when "00100101000001000" => rgb <= "000000";
					when "00100101000001001" => rgb <= "000000";
					when "00100101000001010" => rgb <= "000000";
					when "00100101000001011" => rgb <= "000000";
					when "00100101000001100" => rgb <= "000000";
					when "00100101000001101" => rgb <= "000000";
					when "00100101000001110" => rgb <= "000000";
					when "00100101000001111" => rgb <= "000000";
					when "00100101000010000" => rgb <= "000000";
					when "00100101000010001" => rgb <= "000000";
					when "00100101000010010" => rgb <= "000000";
					when "00100101000010011" => rgb <= "000000";
					when "00100101000010100" => rgb <= "000000";
					when "00100101000010101" => rgb <= "000000";
					when "00100101000010110" => rgb <= "000000";
					when "00100101000010111" => rgb <= "000000";
					when "00100101000011000" => rgb <= "000000";
					when "00100101000011001" => rgb <= "000000";
					when "00100101000011010" => rgb <= "000000";
					when "00100101000011011" => rgb <= "000000";
					when "00100101000011100" => rgb <= "000000";
					when "00100101000011101" => rgb <= "000000";
					when "00100101000011110" => rgb <= "000000";
					when "00100101000011111" => rgb <= "000000";
					when "00100101000100000" => rgb <= "000000";
					when "00100101000100001" => rgb <= "000000";
					when "00100101000100010" => rgb <= "000000";
					when "00100101000100011" => rgb <= "000000";
					when "00100101000100100" => rgb <= "000000";
					when "00100101000100101" => rgb <= "000000";
					when "00100101000100110" => rgb <= "000000";
					when "00100101000100111" => rgb <= "000000";
					when "00100101000101000" => rgb <= "000000";
					when "00100101000101001" => rgb <= "000000";
					when "00100101000101010" => rgb <= "000000";
					when "00100101000101011" => rgb <= "000000";
					when "00100101000101100" => rgb <= "000000";
					when "00100101000101101" => rgb <= "000000";
					when "00100101000101110" => rgb <= "000000";
					when "00100101000101111" => rgb <= "000000";
					when "00100101000110000" => rgb <= "000000";
					when "00100101000110001" => rgb <= "000000";
					when "00100101000110010" => rgb <= "000000";
					when "00100101000110011" => rgb <= "000000";
					when "00100101000110100" => rgb <= "000000";
					when "00100101000110101" => rgb <= "000000";
					when "00100101000110110" => rgb <= "000000";
					when "00100101000110111" => rgb <= "000000";
					when "00100101000111000" => rgb <= "000000";
					when "00100101000111001" => rgb <= "000000";
					when "00100101000111010" => rgb <= "000000";
					when "00100101000111011" => rgb <= "000000";
					when "00100101000111100" => rgb <= "000000";
					when "00100101000111101" => rgb <= "000000";
					when "00100101000111110" => rgb <= "000000";
					when "00100101000111111" => rgb <= "000000";
					when "00100101001000000" => rgb <= "000000";
					when "00100101001000001" => rgb <= "000000";
					when "00100101001000010" => rgb <= "000000";
					when "00100101001000011" => rgb <= "000000";
					when "00100101001000100" => rgb <= "000000";
					when "00100101001000101" => rgb <= "000000";
					when "00100101001000110" => rgb <= "000000";
					when "00100101001000111" => rgb <= "000000";
					when "00100101001001000" => rgb <= "000000";
					when "00100101001001001" => rgb <= "000000";
					when "00100101001001010" => rgb <= "000000";
					when "00100101001001011" => rgb <= "000000";
					when "00100101001001100" => rgb <= "000000";
					when "00100101001001101" => rgb <= "000000";
					when "00100101001001110" => rgb <= "000000";
					when "00100101001001111" => rgb <= "000000";
					when "00100101001010000" => rgb <= "000000";
					when "00100101001010001" => rgb <= "000000";
					when "00100101001010010" => rgb <= "000000";
					when "00100101001010011" => rgb <= "000000";
					when "00100101001010100" => rgb <= "000000";
					when "00100101001010101" => rgb <= "000000";
					when "00100101001010110" => rgb <= "000000";
					when "00100101001010111" => rgb <= "000000";
					when "00100101001011000" => rgb <= "000000";
					when "00100101001011001" => rgb <= "000000";
					when "00100101001011010" => rgb <= "000000";
					when "00100101001011011" => rgb <= "000000";
					when "00100101001011100" => rgb <= "000000";
					when "00100101001011101" => rgb <= "000000";
					when "00100101001011110" => rgb <= "000000";
					when "00100101001011111" => rgb <= "000000";
					when "00100101001100000" => rgb <= "000000";
					when "00100101001100001" => rgb <= "000000";
					when "00100101001100010" => rgb <= "000000";
					when "00100101001100011" => rgb <= "000000";
					when "00100101001100100" => rgb <= "000000";
					when "00100101001100101" => rgb <= "000000";
					when "00100101001100110" => rgb <= "000000";
					when "00100101001100111" => rgb <= "000000";
					when "00100101001101000" => rgb <= "000000";
					when "00100101001101001" => rgb <= "000000";
					when "00100101001101010" => rgb <= "000000";
					when "00100101001101011" => rgb <= "000000";
					when "00100101001101100" => rgb <= "000000";
					when "00100101001101101" => rgb <= "000000";
					when "00100101001101110" => rgb <= "000000";
					when "00100101001101111" => rgb <= "000000";
					when "00100101001110000" => rgb <= "000000";
					when "00100101001110001" => rgb <= "000000";
					when "00100101001110010" => rgb <= "000000";
					when "00100101001110011" => rgb <= "000000";
					when "00100101001110100" => rgb <= "000000";
					when "00100101001110101" => rgb <= "000000";
					when "00100101001110110" => rgb <= "000000";
					when "00100101001110111" => rgb <= "000000";
					when "00100101001111000" => rgb <= "000000";
					when "00100101001111001" => rgb <= "000000";
					when "00100101001111010" => rgb <= "000000";
					when "00100101001111011" => rgb <= "000000";
					when "00100101001111100" => rgb <= "000000";
					when "00100101001111101" => rgb <= "101000";
					when "00100101001111110" => rgb <= "101000";
					when "00100101001111111" => rgb <= "101000";
					when "00100101010000000" => rgb <= "101000";
					when "00100101010000001" => rgb <= "101000";
					when "00100101010000010" => rgb <= "101000";
					when "00100101010000011" => rgb <= "101000";
					when "00100101010000100" => rgb <= "101000";
					when "00100101010000101" => rgb <= "101000";
					when "00100101010000110" => rgb <= "101000";
					when "00100101010000111" => rgb <= "101000";
					when "00100101010001000" => rgb <= "101001";
					when "00100101010001001" => rgb <= "111001";
					when "00100101010001010" => rgb <= "101001";
					when "00100101010001011" => rgb <= "101001";
					when "00100101010001100" => rgb <= "111001";
					when "00100101010001101" => rgb <= "111001";
					when "00100101010001110" => rgb <= "111001";
					when "00100101010001111" => rgb <= "101001";
					when "00100101010010000" => rgb <= "101001";
					when "00100101010010001" => rgb <= "101001";
					when "00100101010010010" => rgb <= "111001";
					when "00100101010010011" => rgb <= "111001";
					when "00100101010010100" => rgb <= "111001";
					when "00100101010010101" => rgb <= "111001";
					when "00100101010010110" => rgb <= "111001";
					when "00100101010010111" => rgb <= "111001";
					when "00100101010011000" => rgb <= "111001";
					when "00100101010011001" => rgb <= "101001";
					when "00100101010011010" => rgb <= "101001";
					when "00100101010011011" => rgb <= "111001";
					when "00100101010011100" => rgb <= "111001";
					when "00100101010011101" => rgb <= "101001";
					when "00100101010011110" => rgb <= "111001";
					when "00100101010011111" => rgb <= "101000";
					when "00100101010100000" => rgb <= "101000";
					when "00100101010100001" => rgb <= "101000";
					when "00100101010100010" => rgb <= "101000";
					when "00100101010100011" => rgb <= "101000";
					when "00100101010100100" => rgb <= "101000";
					when "00100101010100101" => rgb <= "101000";
					when "00100101010100110" => rgb <= "101000";
					when "00100101010100111" => rgb <= "101000";
					when "00100101010101000" => rgb <= "101000";
					when "00100101010101001" => rgb <= "101000";
					when "00100101010101010" => rgb <= "101000";
					when "00100101010101011" => rgb <= "101000";
					when "00100101010101100" => rgb <= "101000";
					when "00100101010101101" => rgb <= "101000";
					when "00100101010101110" => rgb <= "101000";
					when "00100101010101111" => rgb <= "101000";
					when "00100101010110000" => rgb <= "101000";
					when "00100101010110001" => rgb <= "101000";
					when "00100101010110010" => rgb <= "101000";
					when "00100101010110011" => rgb <= "101000";
					when "00100101010110100" => rgb <= "101000";
					when "00100101010110101" => rgb <= "101000";
					when "00100101010110110" => rgb <= "101000";
					when "00100101010110111" => rgb <= "101000";
					when "00100101010111000" => rgb <= "101000";
					when "00100101010111001" => rgb <= "101000";
					when "00100101010111010" => rgb <= "101000";
					when "00100101010111011" => rgb <= "101000";
					when "00100101010111100" => rgb <= "101000";
					when "00100101010111101" => rgb <= "101000";
					when "00100101010111110" => rgb <= "101000";
					when "00100101010111111" => rgb <= "101000";
					when "00100101011000000" => rgb <= "100100";
					when "00100101011000001" => rgb <= "000000";
					when "00100101011000010" => rgb <= "000000";
					when "00100101011000011" => rgb <= "000000";
					when "00100101011000100" => rgb <= "000000";
					when "00100101011000101" => rgb <= "000000";
					when "00100101011000110" => rgb <= "000000";
					when "00100101011000111" => rgb <= "000000";
					when "00100101011001000" => rgb <= "000000";
					when "00100101011001001" => rgb <= "000000";
					when "00100101011001010" => rgb <= "000000";
					when "00100101011001011" => rgb <= "000000";
					when "00100101011001100" => rgb <= "000000";
					when "00100101011001101" => rgb <= "000000";
					when "00100101011001110" => rgb <= "000000";
					when "00100101011001111" => rgb <= "000000";
					when "00100101011010000" => rgb <= "000000";
					when "00100101011010001" => rgb <= "000000";
					when "00100101011010010" => rgb <= "000000";
					when "00100101011010011" => rgb <= "000000";
					when "00100101011010100" => rgb <= "000000";
					when "00100101011010101" => rgb <= "000000";
					when "00100101011010110" => rgb <= "000000";
					when "00100101011010111" => rgb <= "000000";
					when "00100101011011000" => rgb <= "000000";
					when "00100101011011001" => rgb <= "000000";
					when "00100101011011010" => rgb <= "000000";
					when "00100101011011011" => rgb <= "000000";
					when "00100101011011100" => rgb <= "000000";
					when "00100101011011101" => rgb <= "000000";
					when "00100101011011110" => rgb <= "000000";
					when "00100101011011111" => rgb <= "000000";
					when "00100101011100000" => rgb <= "000000";
					when "00100101011100001" => rgb <= "000000";
					when "00100101011100010" => rgb <= "000000";
					when "00100101011100011" => rgb <= "000000";
					when "00100101011100100" => rgb <= "000000";
					when "00100101011100101" => rgb <= "000000";
					when "00100101011100110" => rgb <= "000000";
					when "00100101011100111" => rgb <= "000000";
					when "00100101011101000" => rgb <= "000000";
					when "00100101011101001" => rgb <= "000000";
					when "00100101011101010" => rgb <= "000000";
					when "00100101011101011" => rgb <= "000000";
					when "00100101011101100" => rgb <= "000000";
					when "00100101011101101" => rgb <= "000000";
					when "00100101011101110" => rgb <= "000000";
					when "00100101011101111" => rgb <= "000000";
					when "00100101011110000" => rgb <= "000000";
					when "00100101011110001" => rgb <= "000000";
					when "00100101011110010" => rgb <= "000000";
					when "00100101011110011" => rgb <= "000000";
					when "00100101011110100" => rgb <= "000000";
					when "00100101011110101" => rgb <= "000000";
					when "00100101011110110" => rgb <= "000000";
					when "00100101011110111" => rgb <= "000000";
					when "00100101011111000" => rgb <= "000000";
					when "00100101011111001" => rgb <= "000000";
					when "00100101011111010" => rgb <= "000000";
					when "00100101011111011" => rgb <= "000000";
					when "00100101011111100" => rgb <= "000000";
					when "00100101011111101" => rgb <= "000000";
					when "00100101011111110" => rgb <= "000000";
					when "00100101011111111" => rgb <= "000000";
					when "00100101100000000" => rgb <= "000000";
					when "00100101100000001" => rgb <= "000000";
					when "00100101100000010" => rgb <= "000000";
					when "00100101100000011" => rgb <= "000000";
					when "00100101100000100" => rgb <= "000000";
					when "00100101100000101" => rgb <= "000000";
					when "00100101100000110" => rgb <= "000000";
					when "00100101100000111" => rgb <= "000000";
					when "00100101100001000" => rgb <= "000000";
					when "00100101100001001" => rgb <= "000000";
					when "00100101100001010" => rgb <= "000000";
					when "00100101100001011" => rgb <= "000000";
					when "00100101100001100" => rgb <= "000000";
					when "00100101100001101" => rgb <= "000000";
					when "00100101100001110" => rgb <= "000000";
					when "00100101100001111" => rgb <= "000000";
					when "00100101100010000" => rgb <= "000000";
					when "00100101100010001" => rgb <= "000000";
					when "00100101100010010" => rgb <= "000000";
					when "00100101100010011" => rgb <= "000000";
					when "00100101100010100" => rgb <= "000000";
					when "00100101100010101" => rgb <= "000000";
					when "00100101100010110" => rgb <= "000000";
					when "00100101100010111" => rgb <= "000000";
					when "00100101100011000" => rgb <= "000000";
					when "00100101100011001" => rgb <= "000000";
					when "00100101100011010" => rgb <= "000000";
					when "00100101100011011" => rgb <= "000000";
					when "00100101100011100" => rgb <= "000000";
					when "00100101100011101" => rgb <= "000000";
					when "00100101100011110" => rgb <= "000000";
					when "00100101100011111" => rgb <= "000000";
					when "00100101100100000" => rgb <= "000000";
					when "00100101100100001" => rgb <= "000000";
					when "00100101100100010" => rgb <= "000000";
					when "00100101100100011" => rgb <= "000000";
					when "00100101100100100" => rgb <= "000000";
					when "00100101100100101" => rgb <= "000000";
					when "00100101100100110" => rgb <= "000000";
					when "00100101100100111" => rgb <= "000000";
					when "00100101100101000" => rgb <= "000000";
					when "00100101100101001" => rgb <= "000000";
					when "00100101100101010" => rgb <= "000000";
					when "00100101100101011" => rgb <= "000000";
					when "00100101100101100" => rgb <= "000000";
					when "00100101100101101" => rgb <= "000000";
					when "00100101100101110" => rgb <= "000000";
					when "00100101100101111" => rgb <= "000000";
					when "00100101100110000" => rgb <= "000000";
					when "00100101100110001" => rgb <= "000000";
					when "00100101100110010" => rgb <= "000000";
					when "00100101100110011" => rgb <= "000000";
					when "00100101100110100" => rgb <= "000000";
					when "00100101100110101" => rgb <= "000000";
					when "00100101100110110" => rgb <= "000000";
					when "00100101100110111" => rgb <= "000000";
					when "00100101100111000" => rgb <= "000000";
					when "00100101100111001" => rgb <= "000000";
					when "00100101100111010" => rgb <= "000000";
					when "00100101100111011" => rgb <= "000000";
					when "00100101100111100" => rgb <= "000000";
					when "00100101100111101" => rgb <= "000000";
					when "00100101100111110" => rgb <= "000000";
					when "00100101100111111" => rgb <= "000000";
					when "00100110000000000" => rgb <= "000000";
					when "00100110000000001" => rgb <= "000000";
					when "00100110000000010" => rgb <= "000000";
					when "00100110000000011" => rgb <= "000000";
					when "00100110000000100" => rgb <= "000000";
					when "00100110000000101" => rgb <= "000000";
					when "00100110000000110" => rgb <= "000000";
					when "00100110000000111" => rgb <= "000000";
					when "00100110000001000" => rgb <= "000000";
					when "00100110000001001" => rgb <= "000000";
					when "00100110000001010" => rgb <= "000000";
					when "00100110000001011" => rgb <= "000000";
					when "00100110000001100" => rgb <= "000000";
					when "00100110000001101" => rgb <= "000000";
					when "00100110000001110" => rgb <= "000000";
					when "00100110000001111" => rgb <= "000000";
					when "00100110000010000" => rgb <= "000000";
					when "00100110000010001" => rgb <= "000000";
					when "00100110000010010" => rgb <= "000000";
					when "00100110000010011" => rgb <= "000000";
					when "00100110000010100" => rgb <= "000000";
					when "00100110000010101" => rgb <= "000000";
					when "00100110000010110" => rgb <= "000000";
					when "00100110000010111" => rgb <= "000000";
					when "00100110000011000" => rgb <= "000000";
					when "00100110000011001" => rgb <= "000000";
					when "00100110000011010" => rgb <= "000000";
					when "00100110000011011" => rgb <= "000000";
					when "00100110000011100" => rgb <= "000000";
					when "00100110000011101" => rgb <= "000000";
					when "00100110000011110" => rgb <= "000000";
					when "00100110000011111" => rgb <= "000000";
					when "00100110000100000" => rgb <= "000000";
					when "00100110000100001" => rgb <= "000000";
					when "00100110000100010" => rgb <= "000000";
					when "00100110000100011" => rgb <= "000000";
					when "00100110000100100" => rgb <= "000000";
					when "00100110000100101" => rgb <= "000000";
					when "00100110000100110" => rgb <= "000000";
					when "00100110000100111" => rgb <= "000000";
					when "00100110000101000" => rgb <= "000000";
					when "00100110000101001" => rgb <= "000000";
					when "00100110000101010" => rgb <= "000000";
					when "00100110000101011" => rgb <= "000000";
					when "00100110000101100" => rgb <= "000000";
					when "00100110000101101" => rgb <= "000000";
					when "00100110000101110" => rgb <= "000000";
					when "00100110000101111" => rgb <= "000000";
					when "00100110000110000" => rgb <= "000000";
					when "00100110000110001" => rgb <= "000000";
					when "00100110000110010" => rgb <= "000000";
					when "00100110000110011" => rgb <= "000000";
					when "00100110000110100" => rgb <= "000000";
					when "00100110000110101" => rgb <= "000000";
					when "00100110000110110" => rgb <= "000000";
					when "00100110000110111" => rgb <= "000000";
					when "00100110000111000" => rgb <= "000000";
					when "00100110000111001" => rgb <= "000000";
					when "00100110000111010" => rgb <= "000000";
					when "00100110000111011" => rgb <= "000000";
					when "00100110000111100" => rgb <= "000000";
					when "00100110000111101" => rgb <= "000000";
					when "00100110000111110" => rgb <= "000000";
					when "00100110000111111" => rgb <= "000000";
					when "00100110001000000" => rgb <= "000000";
					when "00100110001000001" => rgb <= "000000";
					when "00100110001000010" => rgb <= "000000";
					when "00100110001000011" => rgb <= "000000";
					when "00100110001000100" => rgb <= "000000";
					when "00100110001000101" => rgb <= "000000";
					when "00100110001000110" => rgb <= "000000";
					when "00100110001000111" => rgb <= "000000";
					when "00100110001001000" => rgb <= "000000";
					when "00100110001001001" => rgb <= "000000";
					when "00100110001001010" => rgb <= "000000";
					when "00100110001001011" => rgb <= "000000";
					when "00100110001001100" => rgb <= "000000";
					when "00100110001001101" => rgb <= "000000";
					when "00100110001001110" => rgb <= "000000";
					when "00100110001001111" => rgb <= "000000";
					when "00100110001010000" => rgb <= "000000";
					when "00100110001010001" => rgb <= "000000";
					when "00100110001010010" => rgb <= "000000";
					when "00100110001010011" => rgb <= "000000";
					when "00100110001010100" => rgb <= "000000";
					when "00100110001010101" => rgb <= "000000";
					when "00100110001010110" => rgb <= "000000";
					when "00100110001010111" => rgb <= "000000";
					when "00100110001011000" => rgb <= "000000";
					when "00100110001011001" => rgb <= "000000";
					when "00100110001011010" => rgb <= "000000";
					when "00100110001011011" => rgb <= "000000";
					when "00100110001011100" => rgb <= "000000";
					when "00100110001011101" => rgb <= "000000";
					when "00100110001011110" => rgb <= "000000";
					when "00100110001011111" => rgb <= "000000";
					when "00100110001100000" => rgb <= "000000";
					when "00100110001100001" => rgb <= "000000";
					when "00100110001100010" => rgb <= "000000";
					when "00100110001100011" => rgb <= "000000";
					when "00100110001100100" => rgb <= "000000";
					when "00100110001100101" => rgb <= "000000";
					when "00100110001100110" => rgb <= "000000";
					when "00100110001100111" => rgb <= "000000";
					when "00100110001101000" => rgb <= "000000";
					when "00100110001101001" => rgb <= "000000";
					when "00100110001101010" => rgb <= "000000";
					when "00100110001101011" => rgb <= "000000";
					when "00100110001101100" => rgb <= "000000";
					when "00100110001101101" => rgb <= "000000";
					when "00100110001101110" => rgb <= "000000";
					when "00100110001101111" => rgb <= "000000";
					when "00100110001110000" => rgb <= "000000";
					when "00100110001110001" => rgb <= "000000";
					when "00100110001110010" => rgb <= "000000";
					when "00100110001110011" => rgb <= "000000";
					when "00100110001110100" => rgb <= "000000";
					when "00100110001110101" => rgb <= "000000";
					when "00100110001110110" => rgb <= "000000";
					when "00100110001110111" => rgb <= "000000";
					when "00100110001111000" => rgb <= "000000";
					when "00100110001111001" => rgb <= "000000";
					when "00100110001111010" => rgb <= "000000";
					when "00100110001111011" => rgb <= "000000";
					when "00100110001111100" => rgb <= "000000";
					when "00100110001111101" => rgb <= "101000";
					when "00100110001111110" => rgb <= "101000";
					when "00100110001111111" => rgb <= "101000";
					when "00100110010000000" => rgb <= "101000";
					when "00100110010000001" => rgb <= "101000";
					when "00100110010000010" => rgb <= "101000";
					when "00100110010000011" => rgb <= "101000";
					when "00100110010000100" => rgb <= "101000";
					when "00100110010000101" => rgb <= "101000";
					when "00100110010000110" => rgb <= "101000";
					when "00100110010000111" => rgb <= "101000";
					when "00100110010001000" => rgb <= "101001";
					when "00100110010001001" => rgb <= "111001";
					when "00100110010001010" => rgb <= "101001";
					when "00100110010001011" => rgb <= "101001";
					when "00100110010001100" => rgb <= "111001";
					when "00100110010001101" => rgb <= "111001";
					when "00100110010001110" => rgb <= "111001";
					when "00100110010001111" => rgb <= "101001";
					when "00100110010010000" => rgb <= "111001";
					when "00100110010010001" => rgb <= "111001";
					when "00100110010010010" => rgb <= "111001";
					when "00100110010010011" => rgb <= "111001";
					when "00100110010010100" => rgb <= "111001";
					when "00100110010010101" => rgb <= "111001";
					when "00100110010010110" => rgb <= "101001";
					when "00100110010010111" => rgb <= "101001";
					when "00100110010011000" => rgb <= "111001";
					when "00100110010011001" => rgb <= "101001";
					when "00100110010011010" => rgb <= "101001";
					when "00100110010011011" => rgb <= "111001";
					when "00100110010011100" => rgb <= "111001";
					when "00100110010011101" => rgb <= "101001";
					when "00100110010011110" => rgb <= "111001";
					when "00100110010011111" => rgb <= "101000";
					when "00100110010100000" => rgb <= "101000";
					when "00100110010100001" => rgb <= "101000";
					when "00100110010100010" => rgb <= "101000";
					when "00100110010100011" => rgb <= "101000";
					when "00100110010100100" => rgb <= "101000";
					when "00100110010100101" => rgb <= "101000";
					when "00100110010100110" => rgb <= "101000";
					when "00100110010100111" => rgb <= "101000";
					when "00100110010101000" => rgb <= "101000";
					when "00100110010101001" => rgb <= "101000";
					when "00100110010101010" => rgb <= "101000";
					when "00100110010101011" => rgb <= "101000";
					when "00100110010101100" => rgb <= "101000";
					when "00100110010101101" => rgb <= "101000";
					when "00100110010101110" => rgb <= "101000";
					when "00100110010101111" => rgb <= "101000";
					when "00100110010110000" => rgb <= "101000";
					when "00100110010110001" => rgb <= "101000";
					when "00100110010110010" => rgb <= "101000";
					when "00100110010110011" => rgb <= "101000";
					when "00100110010110100" => rgb <= "101000";
					when "00100110010110101" => rgb <= "101000";
					when "00100110010110110" => rgb <= "101000";
					when "00100110010110111" => rgb <= "101000";
					when "00100110010111000" => rgb <= "101000";
					when "00100110010111001" => rgb <= "101000";
					when "00100110010111010" => rgb <= "101000";
					when "00100110010111011" => rgb <= "101000";
					when "00100110010111100" => rgb <= "101000";
					when "00100110010111101" => rgb <= "101000";
					when "00100110010111110" => rgb <= "101000";
					when "00100110010111111" => rgb <= "101000";
					when "00100110011000000" => rgb <= "100100";
					when "00100110011000001" => rgb <= "000000";
					when "00100110011000010" => rgb <= "000000";
					when "00100110011000011" => rgb <= "000000";
					when "00100110011000100" => rgb <= "000000";
					when "00100110011000101" => rgb <= "000000";
					when "00100110011000110" => rgb <= "000000";
					when "00100110011000111" => rgb <= "000000";
					when "00100110011001000" => rgb <= "000000";
					when "00100110011001001" => rgb <= "000000";
					when "00100110011001010" => rgb <= "000000";
					when "00100110011001011" => rgb <= "000000";
					when "00100110011001100" => rgb <= "000000";
					when "00100110011001101" => rgb <= "000000";
					when "00100110011001110" => rgb <= "000000";
					when "00100110011001111" => rgb <= "000000";
					when "00100110011010000" => rgb <= "000000";
					when "00100110011010001" => rgb <= "000000";
					when "00100110011010010" => rgb <= "000000";
					when "00100110011010011" => rgb <= "000000";
					when "00100110011010100" => rgb <= "000000";
					when "00100110011010101" => rgb <= "000000";
					when "00100110011010110" => rgb <= "000000";
					when "00100110011010111" => rgb <= "000000";
					when "00100110011011000" => rgb <= "000000";
					when "00100110011011001" => rgb <= "000000";
					when "00100110011011010" => rgb <= "000000";
					when "00100110011011011" => rgb <= "000000";
					when "00100110011011100" => rgb <= "000000";
					when "00100110011011101" => rgb <= "000000";
					when "00100110011011110" => rgb <= "000000";
					when "00100110011011111" => rgb <= "000000";
					when "00100110011100000" => rgb <= "000000";
					when "00100110011100001" => rgb <= "000000";
					when "00100110011100010" => rgb <= "000000";
					when "00100110011100011" => rgb <= "000000";
					when "00100110011100100" => rgb <= "000000";
					when "00100110011100101" => rgb <= "000000";
					when "00100110011100110" => rgb <= "000000";
					when "00100110011100111" => rgb <= "000000";
					when "00100110011101000" => rgb <= "000000";
					when "00100110011101001" => rgb <= "000000";
					when "00100110011101010" => rgb <= "000000";
					when "00100110011101011" => rgb <= "000000";
					when "00100110011101100" => rgb <= "000000";
					when "00100110011101101" => rgb <= "000000";
					when "00100110011101110" => rgb <= "000000";
					when "00100110011101111" => rgb <= "000000";
					when "00100110011110000" => rgb <= "000000";
					when "00100110011110001" => rgb <= "000000";
					when "00100110011110010" => rgb <= "000000";
					when "00100110011110011" => rgb <= "000000";
					when "00100110011110100" => rgb <= "000000";
					when "00100110011110101" => rgb <= "000000";
					when "00100110011110110" => rgb <= "000000";
					when "00100110011110111" => rgb <= "000000";
					when "00100110011111000" => rgb <= "000000";
					when "00100110011111001" => rgb <= "000000";
					when "00100110011111010" => rgb <= "000000";
					when "00100110011111011" => rgb <= "000000";
					when "00100110011111100" => rgb <= "000000";
					when "00100110011111101" => rgb <= "000000";
					when "00100110011111110" => rgb <= "000000";
					when "00100110011111111" => rgb <= "000000";
					when "00100110100000000" => rgb <= "000000";
					when "00100110100000001" => rgb <= "000000";
					when "00100110100000010" => rgb <= "000000";
					when "00100110100000011" => rgb <= "000000";
					when "00100110100000100" => rgb <= "000000";
					when "00100110100000101" => rgb <= "000000";
					when "00100110100000110" => rgb <= "000000";
					when "00100110100000111" => rgb <= "000000";
					when "00100110100001000" => rgb <= "000000";
					when "00100110100001001" => rgb <= "000000";
					when "00100110100001010" => rgb <= "000000";
					when "00100110100001011" => rgb <= "000000";
					when "00100110100001100" => rgb <= "000000";
					when "00100110100001101" => rgb <= "000000";
					when "00100110100001110" => rgb <= "000000";
					when "00100110100001111" => rgb <= "000000";
					when "00100110100010000" => rgb <= "000000";
					when "00100110100010001" => rgb <= "000000";
					when "00100110100010010" => rgb <= "000000";
					when "00100110100010011" => rgb <= "000000";
					when "00100110100010100" => rgb <= "000000";
					when "00100110100010101" => rgb <= "000000";
					when "00100110100010110" => rgb <= "000000";
					when "00100110100010111" => rgb <= "000000";
					when "00100110100011000" => rgb <= "000000";
					when "00100110100011001" => rgb <= "000000";
					when "00100110100011010" => rgb <= "000000";
					when "00100110100011011" => rgb <= "000000";
					when "00100110100011100" => rgb <= "000000";
					when "00100110100011101" => rgb <= "000000";
					when "00100110100011110" => rgb <= "000000";
					when "00100110100011111" => rgb <= "000000";
					when "00100110100100000" => rgb <= "000000";
					when "00100110100100001" => rgb <= "000000";
					when "00100110100100010" => rgb <= "000000";
					when "00100110100100011" => rgb <= "000000";
					when "00100110100100100" => rgb <= "000000";
					when "00100110100100101" => rgb <= "000000";
					when "00100110100100110" => rgb <= "000000";
					when "00100110100100111" => rgb <= "000000";
					when "00100110100101000" => rgb <= "000000";
					when "00100110100101001" => rgb <= "000000";
					when "00100110100101010" => rgb <= "000000";
					when "00100110100101011" => rgb <= "000000";
					when "00100110100101100" => rgb <= "000000";
					when "00100110100101101" => rgb <= "000000";
					when "00100110100101110" => rgb <= "000000";
					when "00100110100101111" => rgb <= "000000";
					when "00100110100110000" => rgb <= "000000";
					when "00100110100110001" => rgb <= "000000";
					when "00100110100110010" => rgb <= "000000";
					when "00100110100110011" => rgb <= "000000";
					when "00100110100110100" => rgb <= "000000";
					when "00100110100110101" => rgb <= "000000";
					when "00100110100110110" => rgb <= "000000";
					when "00100110100110111" => rgb <= "000000";
					when "00100110100111000" => rgb <= "000000";
					when "00100110100111001" => rgb <= "000000";
					when "00100110100111010" => rgb <= "000000";
					when "00100110100111011" => rgb <= "000000";
					when "00100110100111100" => rgb <= "000000";
					when "00100110100111101" => rgb <= "000000";
					when "00100110100111110" => rgb <= "000000";
					when "00100110100111111" => rgb <= "000000";
					when "00100111000000000" => rgb <= "000000";
					when "00100111000000001" => rgb <= "000000";
					when "00100111000000010" => rgb <= "000000";
					when "00100111000000011" => rgb <= "000000";
					when "00100111000000100" => rgb <= "000000";
					when "00100111000000101" => rgb <= "000000";
					when "00100111000000110" => rgb <= "000000";
					when "00100111000000111" => rgb <= "000000";
					when "00100111000001000" => rgb <= "000000";
					when "00100111000001001" => rgb <= "000000";
					when "00100111000001010" => rgb <= "000000";
					when "00100111000001011" => rgb <= "000000";
					when "00100111000001100" => rgb <= "000000";
					when "00100111000001101" => rgb <= "000000";
					when "00100111000001110" => rgb <= "000000";
					when "00100111000001111" => rgb <= "000000";
					when "00100111000010000" => rgb <= "000000";
					when "00100111000010001" => rgb <= "000000";
					when "00100111000010010" => rgb <= "000000";
					when "00100111000010011" => rgb <= "000000";
					when "00100111000010100" => rgb <= "000000";
					when "00100111000010101" => rgb <= "000000";
					when "00100111000010110" => rgb <= "000000";
					when "00100111000010111" => rgb <= "000000";
					when "00100111000011000" => rgb <= "000000";
					when "00100111000011001" => rgb <= "000000";
					when "00100111000011010" => rgb <= "000000";
					when "00100111000011011" => rgb <= "000000";
					when "00100111000011100" => rgb <= "000000";
					when "00100111000011101" => rgb <= "000000";
					when "00100111000011110" => rgb <= "000000";
					when "00100111000011111" => rgb <= "000000";
					when "00100111000100000" => rgb <= "000000";
					when "00100111000100001" => rgb <= "000000";
					when "00100111000100010" => rgb <= "000000";
					when "00100111000100011" => rgb <= "000000";
					when "00100111000100100" => rgb <= "000000";
					when "00100111000100101" => rgb <= "000000";
					when "00100111000100110" => rgb <= "000000";
					when "00100111000100111" => rgb <= "000000";
					when "00100111000101000" => rgb <= "000000";
					when "00100111000101001" => rgb <= "000000";
					when "00100111000101010" => rgb <= "000000";
					when "00100111000101011" => rgb <= "000000";
					when "00100111000101100" => rgb <= "000000";
					when "00100111000101101" => rgb <= "000000";
					when "00100111000101110" => rgb <= "000000";
					when "00100111000101111" => rgb <= "000000";
					when "00100111000110000" => rgb <= "000000";
					when "00100111000110001" => rgb <= "000000";
					when "00100111000110010" => rgb <= "000000";
					when "00100111000110011" => rgb <= "000000";
					when "00100111000110100" => rgb <= "000000";
					when "00100111000110101" => rgb <= "000000";
					when "00100111000110110" => rgb <= "000000";
					when "00100111000110111" => rgb <= "000000";
					when "00100111000111000" => rgb <= "000000";
					when "00100111000111001" => rgb <= "000000";
					when "00100111000111010" => rgb <= "000000";
					when "00100111000111011" => rgb <= "000000";
					when "00100111000111100" => rgb <= "000000";
					when "00100111000111101" => rgb <= "000000";
					when "00100111000111110" => rgb <= "000000";
					when "00100111000111111" => rgb <= "000000";
					when "00100111001000000" => rgb <= "000000";
					when "00100111001000001" => rgb <= "000000";
					when "00100111001000010" => rgb <= "000000";
					when "00100111001000011" => rgb <= "000000";
					when "00100111001000100" => rgb <= "000000";
					when "00100111001000101" => rgb <= "000000";
					when "00100111001000110" => rgb <= "000000";
					when "00100111001000111" => rgb <= "000000";
					when "00100111001001000" => rgb <= "000000";
					when "00100111001001001" => rgb <= "000000";
					when "00100111001001010" => rgb <= "000000";
					when "00100111001001011" => rgb <= "000000";
					when "00100111001001100" => rgb <= "000000";
					when "00100111001001101" => rgb <= "000000";
					when "00100111001001110" => rgb <= "000000";
					when "00100111001001111" => rgb <= "000000";
					when "00100111001010000" => rgb <= "000000";
					when "00100111001010001" => rgb <= "000000";
					when "00100111001010010" => rgb <= "000000";
					when "00100111001010011" => rgb <= "000000";
					when "00100111001010100" => rgb <= "000000";
					when "00100111001010101" => rgb <= "000000";
					when "00100111001010110" => rgb <= "000000";
					when "00100111001010111" => rgb <= "000000";
					when "00100111001011000" => rgb <= "000000";
					when "00100111001011001" => rgb <= "000000";
					when "00100111001011010" => rgb <= "000000";
					when "00100111001011011" => rgb <= "000000";
					when "00100111001011100" => rgb <= "000000";
					when "00100111001011101" => rgb <= "000000";
					when "00100111001011110" => rgb <= "000000";
					when "00100111001011111" => rgb <= "000000";
					when "00100111001100000" => rgb <= "000000";
					when "00100111001100001" => rgb <= "000000";
					when "00100111001100010" => rgb <= "000000";
					when "00100111001100011" => rgb <= "000000";
					when "00100111001100100" => rgb <= "000000";
					when "00100111001100101" => rgb <= "000000";
					when "00100111001100110" => rgb <= "000000";
					when "00100111001100111" => rgb <= "000000";
					when "00100111001101000" => rgb <= "000000";
					when "00100111001101001" => rgb <= "000000";
					when "00100111001101010" => rgb <= "000000";
					when "00100111001101011" => rgb <= "000000";
					when "00100111001101100" => rgb <= "000000";
					when "00100111001101101" => rgb <= "000000";
					when "00100111001101110" => rgb <= "000000";
					when "00100111001101111" => rgb <= "000000";
					when "00100111001110000" => rgb <= "000000";
					when "00100111001110001" => rgb <= "000000";
					when "00100111001110010" => rgb <= "000000";
					when "00100111001110011" => rgb <= "000000";
					when "00100111001110100" => rgb <= "000000";
					when "00100111001110101" => rgb <= "000000";
					when "00100111001110110" => rgb <= "000000";
					when "00100111001110111" => rgb <= "000000";
					when "00100111001111000" => rgb <= "000000";
					when "00100111001111001" => rgb <= "000000";
					when "00100111001111010" => rgb <= "000000";
					when "00100111001111011" => rgb <= "000000";
					when "00100111001111100" => rgb <= "010000";
					when "00100111001111101" => rgb <= "101000";
					when "00100111001111110" => rgb <= "101000";
					when "00100111001111111" => rgb <= "101000";
					when "00100111010000000" => rgb <= "101000";
					when "00100111010000001" => rgb <= "101000";
					when "00100111010000010" => rgb <= "101000";
					when "00100111010000011" => rgb <= "101000";
					when "00100111010000100" => rgb <= "101000";
					when "00100111010000101" => rgb <= "101000";
					when "00100111010000110" => rgb <= "101000";
					when "00100111010000111" => rgb <= "101000";
					when "00100111010001000" => rgb <= "101001";
					when "00100111010001001" => rgb <= "111001";
					when "00100111010001010" => rgb <= "101001";
					when "00100111010001011" => rgb <= "101001";
					when "00100111010001100" => rgb <= "111001";
					when "00100111010001101" => rgb <= "111001";
					when "00100111010001110" => rgb <= "111001";
					when "00100111010001111" => rgb <= "101001";
					when "00100111010010000" => rgb <= "111001";
					when "00100111010010001" => rgb <= "101001";
					when "00100111010010010" => rgb <= "101001";
					when "00100111010010011" => rgb <= "101001";
					when "00100111010010100" => rgb <= "101001";
					when "00100111010010101" => rgb <= "101001";
					when "00100111010010110" => rgb <= "101001";
					when "00100111010010111" => rgb <= "101001";
					when "00100111010011000" => rgb <= "101001";
					when "00100111010011001" => rgb <= "101001";
					when "00100111010011010" => rgb <= "101001";
					when "00100111010011011" => rgb <= "101001";
					when "00100111010011100" => rgb <= "101001";
					when "00100111010011101" => rgb <= "101001";
					when "00100111010011110" => rgb <= "101001";
					when "00100111010011111" => rgb <= "101000";
					when "00100111010100000" => rgb <= "101000";
					when "00100111010100001" => rgb <= "101000";
					when "00100111010100010" => rgb <= "101000";
					when "00100111010100011" => rgb <= "101000";
					when "00100111010100100" => rgb <= "101000";
					when "00100111010100101" => rgb <= "101000";
					when "00100111010100110" => rgb <= "101000";
					when "00100111010100111" => rgb <= "101000";
					when "00100111010101000" => rgb <= "101000";
					when "00100111010101001" => rgb <= "101000";
					when "00100111010101010" => rgb <= "101000";
					when "00100111010101011" => rgb <= "101000";
					when "00100111010101100" => rgb <= "101000";
					when "00100111010101101" => rgb <= "101000";
					when "00100111010101110" => rgb <= "101000";
					when "00100111010101111" => rgb <= "101000";
					when "00100111010110000" => rgb <= "101000";
					when "00100111010110001" => rgb <= "101000";
					when "00100111010110010" => rgb <= "101000";
					when "00100111010110011" => rgb <= "101000";
					when "00100111010110100" => rgb <= "101000";
					when "00100111010110101" => rgb <= "101000";
					when "00100111010110110" => rgb <= "101000";
					when "00100111010110111" => rgb <= "101000";
					when "00100111010111000" => rgb <= "101000";
					when "00100111010111001" => rgb <= "101000";
					when "00100111010111010" => rgb <= "101000";
					when "00100111010111011" => rgb <= "101000";
					when "00100111010111100" => rgb <= "101000";
					when "00100111010111101" => rgb <= "101000";
					when "00100111010111110" => rgb <= "101000";
					when "00100111010111111" => rgb <= "101000";
					when "00100111011000000" => rgb <= "101000";
					when "00100111011000001" => rgb <= "000000";
					when "00100111011000010" => rgb <= "000000";
					when "00100111011000011" => rgb <= "000000";
					when "00100111011000100" => rgb <= "000000";
					when "00100111011000101" => rgb <= "000000";
					when "00100111011000110" => rgb <= "000000";
					when "00100111011000111" => rgb <= "000000";
					when "00100111011001000" => rgb <= "000000";
					when "00100111011001001" => rgb <= "000000";
					when "00100111011001010" => rgb <= "000000";
					when "00100111011001011" => rgb <= "000000";
					when "00100111011001100" => rgb <= "000000";
					when "00100111011001101" => rgb <= "000000";
					when "00100111011001110" => rgb <= "000000";
					when "00100111011001111" => rgb <= "000000";
					when "00100111011010000" => rgb <= "000000";
					when "00100111011010001" => rgb <= "000000";
					when "00100111011010010" => rgb <= "000000";
					when "00100111011010011" => rgb <= "000000";
					when "00100111011010100" => rgb <= "000000";
					when "00100111011010101" => rgb <= "000000";
					when "00100111011010110" => rgb <= "000000";
					when "00100111011010111" => rgb <= "000000";
					when "00100111011011000" => rgb <= "000000";
					when "00100111011011001" => rgb <= "000000";
					when "00100111011011010" => rgb <= "000000";
					when "00100111011011011" => rgb <= "000000";
					when "00100111011011100" => rgb <= "000000";
					when "00100111011011101" => rgb <= "000000";
					when "00100111011011110" => rgb <= "000000";
					when "00100111011011111" => rgb <= "000000";
					when "00100111011100000" => rgb <= "000000";
					when "00100111011100001" => rgb <= "000000";
					when "00100111011100010" => rgb <= "000000";
					when "00100111011100011" => rgb <= "000000";
					when "00100111011100100" => rgb <= "000000";
					when "00100111011100101" => rgb <= "000000";
					when "00100111011100110" => rgb <= "000000";
					when "00100111011100111" => rgb <= "000000";
					when "00100111011101000" => rgb <= "000000";
					when "00100111011101001" => rgb <= "000000";
					when "00100111011101010" => rgb <= "000000";
					when "00100111011101011" => rgb <= "000000";
					when "00100111011101100" => rgb <= "000000";
					when "00100111011101101" => rgb <= "000000";
					when "00100111011101110" => rgb <= "000000";
					when "00100111011101111" => rgb <= "000000";
					when "00100111011110000" => rgb <= "000000";
					when "00100111011110001" => rgb <= "000000";
					when "00100111011110010" => rgb <= "000000";
					when "00100111011110011" => rgb <= "000000";
					when "00100111011110100" => rgb <= "000000";
					when "00100111011110101" => rgb <= "000000";
					when "00100111011110110" => rgb <= "000000";
					when "00100111011110111" => rgb <= "000000";
					when "00100111011111000" => rgb <= "000000";
					when "00100111011111001" => rgb <= "000000";
					when "00100111011111010" => rgb <= "000000";
					when "00100111011111011" => rgb <= "000000";
					when "00100111011111100" => rgb <= "000000";
					when "00100111011111101" => rgb <= "000000";
					when "00100111011111110" => rgb <= "000000";
					when "00100111011111111" => rgb <= "000000";
					when "00100111100000000" => rgb <= "000000";
					when "00100111100000001" => rgb <= "000000";
					when "00100111100000010" => rgb <= "000000";
					when "00100111100000011" => rgb <= "000000";
					when "00100111100000100" => rgb <= "000000";
					when "00100111100000101" => rgb <= "000000";
					when "00100111100000110" => rgb <= "000000";
					when "00100111100000111" => rgb <= "000000";
					when "00100111100001000" => rgb <= "000000";
					when "00100111100001001" => rgb <= "000000";
					when "00100111100001010" => rgb <= "000000";
					when "00100111100001011" => rgb <= "000000";
					when "00100111100001100" => rgb <= "000000";
					when "00100111100001101" => rgb <= "000000";
					when "00100111100001110" => rgb <= "000000";
					when "00100111100001111" => rgb <= "000000";
					when "00100111100010000" => rgb <= "000000";
					when "00100111100010001" => rgb <= "000000";
					when "00100111100010010" => rgb <= "000000";
					when "00100111100010011" => rgb <= "000000";
					when "00100111100010100" => rgb <= "000000";
					when "00100111100010101" => rgb <= "000000";
					when "00100111100010110" => rgb <= "000000";
					when "00100111100010111" => rgb <= "000000";
					when "00100111100011000" => rgb <= "000000";
					when "00100111100011001" => rgb <= "000000";
					when "00100111100011010" => rgb <= "000000";
					when "00100111100011011" => rgb <= "000000";
					when "00100111100011100" => rgb <= "000000";
					when "00100111100011101" => rgb <= "000000";
					when "00100111100011110" => rgb <= "000000";
					when "00100111100011111" => rgb <= "000000";
					when "00100111100100000" => rgb <= "000000";
					when "00100111100100001" => rgb <= "000000";
					when "00100111100100010" => rgb <= "000000";
					when "00100111100100011" => rgb <= "000000";
					when "00100111100100100" => rgb <= "000000";
					when "00100111100100101" => rgb <= "000000";
					when "00100111100100110" => rgb <= "000000";
					when "00100111100100111" => rgb <= "000000";
					when "00100111100101000" => rgb <= "000000";
					when "00100111100101001" => rgb <= "000000";
					when "00100111100101010" => rgb <= "000000";
					when "00100111100101011" => rgb <= "000000";
					when "00100111100101100" => rgb <= "000000";
					when "00100111100101101" => rgb <= "000000";
					when "00100111100101110" => rgb <= "000000";
					when "00100111100101111" => rgb <= "000000";
					when "00100111100110000" => rgb <= "000000";
					when "00100111100110001" => rgb <= "000000";
					when "00100111100110010" => rgb <= "000000";
					when "00100111100110011" => rgb <= "000000";
					when "00100111100110100" => rgb <= "000000";
					when "00100111100110101" => rgb <= "000000";
					when "00100111100110110" => rgb <= "000000";
					when "00100111100110111" => rgb <= "000000";
					when "00100111100111000" => rgb <= "000000";
					when "00100111100111001" => rgb <= "000000";
					when "00100111100111010" => rgb <= "000000";
					when "00100111100111011" => rgb <= "000000";
					when "00100111100111100" => rgb <= "000000";
					when "00100111100111101" => rgb <= "000000";
					when "00100111100111110" => rgb <= "000000";
					when "00100111100111111" => rgb <= "000000";
					when "00101000000000000" => rgb <= "000000";
					when "00101000000000001" => rgb <= "000000";
					when "00101000000000010" => rgb <= "000000";
					when "00101000000000011" => rgb <= "000000";
					when "00101000000000100" => rgb <= "000000";
					when "00101000000000101" => rgb <= "000000";
					when "00101000000000110" => rgb <= "000000";
					when "00101000000000111" => rgb <= "000000";
					when "00101000000001000" => rgb <= "000000";
					when "00101000000001001" => rgb <= "000000";
					when "00101000000001010" => rgb <= "000000";
					when "00101000000001011" => rgb <= "000000";
					when "00101000000001100" => rgb <= "000000";
					when "00101000000001101" => rgb <= "000000";
					when "00101000000001110" => rgb <= "000000";
					when "00101000000001111" => rgb <= "000000";
					when "00101000000010000" => rgb <= "000000";
					when "00101000000010001" => rgb <= "000000";
					when "00101000000010010" => rgb <= "000000";
					when "00101000000010011" => rgb <= "000000";
					when "00101000000010100" => rgb <= "000000";
					when "00101000000010101" => rgb <= "000000";
					when "00101000000010110" => rgb <= "000000";
					when "00101000000010111" => rgb <= "000000";
					when "00101000000011000" => rgb <= "000000";
					when "00101000000011001" => rgb <= "000000";
					when "00101000000011010" => rgb <= "000000";
					when "00101000000011011" => rgb <= "000000";
					when "00101000000011100" => rgb <= "000000";
					when "00101000000011101" => rgb <= "000000";
					when "00101000000011110" => rgb <= "000000";
					when "00101000000011111" => rgb <= "000000";
					when "00101000000100000" => rgb <= "000000";
					when "00101000000100001" => rgb <= "000000";
					when "00101000000100010" => rgb <= "000000";
					when "00101000000100011" => rgb <= "000000";
					when "00101000000100100" => rgb <= "000000";
					when "00101000000100101" => rgb <= "000000";
					when "00101000000100110" => rgb <= "000000";
					when "00101000000100111" => rgb <= "000000";
					when "00101000000101000" => rgb <= "000000";
					when "00101000000101001" => rgb <= "000000";
					when "00101000000101010" => rgb <= "000000";
					when "00101000000101011" => rgb <= "000000";
					when "00101000000101100" => rgb <= "000000";
					when "00101000000101101" => rgb <= "000000";
					when "00101000000101110" => rgb <= "000000";
					when "00101000000101111" => rgb <= "000000";
					when "00101000000110000" => rgb <= "000000";
					when "00101000000110001" => rgb <= "000000";
					when "00101000000110010" => rgb <= "000000";
					when "00101000000110011" => rgb <= "000000";
					when "00101000000110100" => rgb <= "000000";
					when "00101000000110101" => rgb <= "000000";
					when "00101000000110110" => rgb <= "000000";
					when "00101000000110111" => rgb <= "000000";
					when "00101000000111000" => rgb <= "000000";
					when "00101000000111001" => rgb <= "000000";
					when "00101000000111010" => rgb <= "000000";
					when "00101000000111011" => rgb <= "000000";
					when "00101000000111100" => rgb <= "000000";
					when "00101000000111101" => rgb <= "000000";
					when "00101000000111110" => rgb <= "000000";
					when "00101000000111111" => rgb <= "000000";
					when "00101000001000000" => rgb <= "000000";
					when "00101000001000001" => rgb <= "000000";
					when "00101000001000010" => rgb <= "000000";
					when "00101000001000011" => rgb <= "000000";
					when "00101000001000100" => rgb <= "000000";
					when "00101000001000101" => rgb <= "000000";
					when "00101000001000110" => rgb <= "000000";
					when "00101000001000111" => rgb <= "000000";
					when "00101000001001000" => rgb <= "000000";
					when "00101000001001001" => rgb <= "000000";
					when "00101000001001010" => rgb <= "000000";
					when "00101000001001011" => rgb <= "000000";
					when "00101000001001100" => rgb <= "000000";
					when "00101000001001101" => rgb <= "000000";
					when "00101000001001110" => rgb <= "000000";
					when "00101000001001111" => rgb <= "000000";
					when "00101000001010000" => rgb <= "000000";
					when "00101000001010001" => rgb <= "000000";
					when "00101000001010010" => rgb <= "000000";
					when "00101000001010011" => rgb <= "000000";
					when "00101000001010100" => rgb <= "000000";
					when "00101000001010101" => rgb <= "000000";
					when "00101000001010110" => rgb <= "000000";
					when "00101000001010111" => rgb <= "000000";
					when "00101000001011000" => rgb <= "000000";
					when "00101000001011001" => rgb <= "000000";
					when "00101000001011010" => rgb <= "000000";
					when "00101000001011011" => rgb <= "000000";
					when "00101000001011100" => rgb <= "000000";
					when "00101000001011101" => rgb <= "000000";
					when "00101000001011110" => rgb <= "000000";
					when "00101000001011111" => rgb <= "000000";
					when "00101000001100000" => rgb <= "000000";
					when "00101000001100001" => rgb <= "000000";
					when "00101000001100010" => rgb <= "000000";
					when "00101000001100011" => rgb <= "000000";
					when "00101000001100100" => rgb <= "000000";
					when "00101000001100101" => rgb <= "000000";
					when "00101000001100110" => rgb <= "010100";
					when "00101000001100111" => rgb <= "111000";
					when "00101000001101000" => rgb <= "101000";
					when "00101000001101001" => rgb <= "101000";
					when "00101000001101010" => rgb <= "101000";
					when "00101000001101011" => rgb <= "101000";
					when "00101000001101100" => rgb <= "101000";
					when "00101000001101101" => rgb <= "101000";
					when "00101000001101110" => rgb <= "101000";
					when "00101000001101111" => rgb <= "101000";
					when "00101000001110000" => rgb <= "101000";
					when "00101000001110001" => rgb <= "101000";
					when "00101000001110010" => rgb <= "101000";
					when "00101000001110011" => rgb <= "101000";
					when "00101000001110100" => rgb <= "101000";
					when "00101000001110101" => rgb <= "101000";
					when "00101000001110110" => rgb <= "101000";
					when "00101000001110111" => rgb <= "101000";
					when "00101000001111000" => rgb <= "101000";
					when "00101000001111001" => rgb <= "101000";
					when "00101000001111010" => rgb <= "101000";
					when "00101000001111011" => rgb <= "101000";
					when "00101000001111100" => rgb <= "101000";
					when "00101000001111101" => rgb <= "101000";
					when "00101000001111110" => rgb <= "101000";
					when "00101000001111111" => rgb <= "101000";
					when "00101000010000000" => rgb <= "101000";
					when "00101000010000001" => rgb <= "101000";
					when "00101000010000010" => rgb <= "101000";
					when "00101000010000011" => rgb <= "101000";
					when "00101000010000100" => rgb <= "101000";
					when "00101000010000101" => rgb <= "101000";
					when "00101000010000110" => rgb <= "101000";
					when "00101000010000111" => rgb <= "101000";
					when "00101000010001000" => rgb <= "101001";
					when "00101000010001001" => rgb <= "111001";
					when "00101000010001010" => rgb <= "101001";
					when "00101000010001011" => rgb <= "101001";
					when "00101000010001100" => rgb <= "111001";
					when "00101000010001101" => rgb <= "111001";
					when "00101000010001110" => rgb <= "111001";
					when "00101000010001111" => rgb <= "101001";
					when "00101000010010000" => rgb <= "101001";
					when "00101000010010001" => rgb <= "101001";
					when "00101000010010010" => rgb <= "111001";
					when "00101000010010011" => rgb <= "101001";
					when "00101000010010100" => rgb <= "101000";
					when "00101000010010101" => rgb <= "101000";
					when "00101000010010110" => rgb <= "101000";
					when "00101000010010111" => rgb <= "101000";
					when "00101000010011000" => rgb <= "101000";
					when "00101000010011001" => rgb <= "101000";
					when "00101000010011010" => rgb <= "101000";
					when "00101000010011011" => rgb <= "101000";
					when "00101000010011100" => rgb <= "101000";
					when "00101000010011101" => rgb <= "101000";
					when "00101000010011110" => rgb <= "101000";
					when "00101000010011111" => rgb <= "101000";
					when "00101000010100000" => rgb <= "101000";
					when "00101000010100001" => rgb <= "101000";
					when "00101000010100010" => rgb <= "101000";
					when "00101000010100011" => rgb <= "101000";
					when "00101000010100100" => rgb <= "101000";
					when "00101000010100101" => rgb <= "101000";
					when "00101000010100110" => rgb <= "101000";
					when "00101000010100111" => rgb <= "101000";
					when "00101000010101000" => rgb <= "101000";
					when "00101000010101001" => rgb <= "101000";
					when "00101000010101010" => rgb <= "101000";
					when "00101000010101011" => rgb <= "101000";
					when "00101000010101100" => rgb <= "101000";
					when "00101000010101101" => rgb <= "101000";
					when "00101000010101110" => rgb <= "101000";
					when "00101000010101111" => rgb <= "101000";
					when "00101000010110000" => rgb <= "101000";
					when "00101000010110001" => rgb <= "101000";
					when "00101000010110010" => rgb <= "101000";
					when "00101000010110011" => rgb <= "101000";
					when "00101000010110100" => rgb <= "101000";
					when "00101000010110101" => rgb <= "101000";
					when "00101000010110110" => rgb <= "101000";
					when "00101000010110111" => rgb <= "101000";
					when "00101000010111000" => rgb <= "101000";
					when "00101000010111001" => rgb <= "101000";
					when "00101000010111010" => rgb <= "101000";
					when "00101000010111011" => rgb <= "101000";
					when "00101000010111100" => rgb <= "101000";
					when "00101000010111101" => rgb <= "101000";
					when "00101000010111110" => rgb <= "101000";
					when "00101000010111111" => rgb <= "101000";
					when "00101000011000000" => rgb <= "101000";
					when "00101000011000001" => rgb <= "101000";
					when "00101000011000010" => rgb <= "101000";
					when "00101000011000011" => rgb <= "101000";
					when "00101000011000100" => rgb <= "101000";
					when "00101000011000101" => rgb <= "101000";
					when "00101000011000110" => rgb <= "101000";
					when "00101000011000111" => rgb <= "101000";
					when "00101000011001000" => rgb <= "101000";
					when "00101000011001001" => rgb <= "101000";
					when "00101000011001010" => rgb <= "101000";
					when "00101000011001011" => rgb <= "101000";
					when "00101000011001100" => rgb <= "101000";
					when "00101000011001101" => rgb <= "101000";
					when "00101000011001110" => rgb <= "101000";
					when "00101000011001111" => rgb <= "101000";
					when "00101000011010000" => rgb <= "101000";
					when "00101000011010001" => rgb <= "101000";
					when "00101000011010010" => rgb <= "101000";
					when "00101000011010011" => rgb <= "101000";
					when "00101000011010100" => rgb <= "101000";
					when "00101000011010101" => rgb <= "101000";
					when "00101000011010110" => rgb <= "101000";
					when "00101000011010111" => rgb <= "010100";
					when "00101000011011000" => rgb <= "000000";
					when "00101000011011001" => rgb <= "000000";
					when "00101000011011010" => rgb <= "000000";
					when "00101000011011011" => rgb <= "000000";
					when "00101000011011100" => rgb <= "000000";
					when "00101000011011101" => rgb <= "000000";
					when "00101000011011110" => rgb <= "000000";
					when "00101000011011111" => rgb <= "000000";
					when "00101000011100000" => rgb <= "000000";
					when "00101000011100001" => rgb <= "000000";
					when "00101000011100010" => rgb <= "000000";
					when "00101000011100011" => rgb <= "000000";
					when "00101000011100100" => rgb <= "000000";
					when "00101000011100101" => rgb <= "000000";
					when "00101000011100110" => rgb <= "000000";
					when "00101000011100111" => rgb <= "000000";
					when "00101000011101000" => rgb <= "000000";
					when "00101000011101001" => rgb <= "000000";
					when "00101000011101010" => rgb <= "000000";
					when "00101000011101011" => rgb <= "000000";
					when "00101000011101100" => rgb <= "000000";
					when "00101000011101101" => rgb <= "000000";
					when "00101000011101110" => rgb <= "000000";
					when "00101000011101111" => rgb <= "000000";
					when "00101000011110000" => rgb <= "000000";
					when "00101000011110001" => rgb <= "000000";
					when "00101000011110010" => rgb <= "000000";
					when "00101000011110011" => rgb <= "000000";
					when "00101000011110100" => rgb <= "000000";
					when "00101000011110101" => rgb <= "000000";
					when "00101000011110110" => rgb <= "000000";
					when "00101000011110111" => rgb <= "000000";
					when "00101000011111000" => rgb <= "000000";
					when "00101000011111001" => rgb <= "000000";
					when "00101000011111010" => rgb <= "000000";
					when "00101000011111011" => rgb <= "000000";
					when "00101000011111100" => rgb <= "000000";
					when "00101000011111101" => rgb <= "000000";
					when "00101000011111110" => rgb <= "000000";
					when "00101000011111111" => rgb <= "000000";
					when "00101000100000000" => rgb <= "000000";
					when "00101000100000001" => rgb <= "000000";
					when "00101000100000010" => rgb <= "000000";
					when "00101000100000011" => rgb <= "000000";
					when "00101000100000100" => rgb <= "000000";
					when "00101000100000101" => rgb <= "000000";
					when "00101000100000110" => rgb <= "000000";
					when "00101000100000111" => rgb <= "000000";
					when "00101000100001000" => rgb <= "000000";
					when "00101000100001001" => rgb <= "000000";
					when "00101000100001010" => rgb <= "000000";
					when "00101000100001011" => rgb <= "000000";
					when "00101000100001100" => rgb <= "000000";
					when "00101000100001101" => rgb <= "000000";
					when "00101000100001110" => rgb <= "000000";
					when "00101000100001111" => rgb <= "000000";
					when "00101000100010000" => rgb <= "000000";
					when "00101000100010001" => rgb <= "000000";
					when "00101000100010010" => rgb <= "000000";
					when "00101000100010011" => rgb <= "000000";
					when "00101000100010100" => rgb <= "000000";
					when "00101000100010101" => rgb <= "000000";
					when "00101000100010110" => rgb <= "000000";
					when "00101000100010111" => rgb <= "000000";
					when "00101000100011000" => rgb <= "000000";
					when "00101000100011001" => rgb <= "000000";
					when "00101000100011010" => rgb <= "000000";
					when "00101000100011011" => rgb <= "000000";
					when "00101000100011100" => rgb <= "000000";
					when "00101000100011101" => rgb <= "000000";
					when "00101000100011110" => rgb <= "000000";
					when "00101000100011111" => rgb <= "000000";
					when "00101000100100000" => rgb <= "000000";
					when "00101000100100001" => rgb <= "000000";
					when "00101000100100010" => rgb <= "000000";
					when "00101000100100011" => rgb <= "000000";
					when "00101000100100100" => rgb <= "000000";
					when "00101000100100101" => rgb <= "000000";
					when "00101000100100110" => rgb <= "000000";
					when "00101000100100111" => rgb <= "000000";
					when "00101000100101000" => rgb <= "000000";
					when "00101000100101001" => rgb <= "000000";
					when "00101000100101010" => rgb <= "000000";
					when "00101000100101011" => rgb <= "000000";
					when "00101000100101100" => rgb <= "000000";
					when "00101000100101101" => rgb <= "000000";
					when "00101000100101110" => rgb <= "000000";
					when "00101000100101111" => rgb <= "000000";
					when "00101000100110000" => rgb <= "000000";
					when "00101000100110001" => rgb <= "000000";
					when "00101000100110010" => rgb <= "000000";
					when "00101000100110011" => rgb <= "000000";
					when "00101000100110100" => rgb <= "000000";
					when "00101000100110101" => rgb <= "000000";
					when "00101000100110110" => rgb <= "000000";
					when "00101000100110111" => rgb <= "000000";
					when "00101000100111000" => rgb <= "000000";
					when "00101000100111001" => rgb <= "000000";
					when "00101000100111010" => rgb <= "000000";
					when "00101000100111011" => rgb <= "000000";
					when "00101000100111100" => rgb <= "000000";
					when "00101000100111101" => rgb <= "000000";
					when "00101000100111110" => rgb <= "000000";
					when "00101000100111111" => rgb <= "000000";
					when "00101001000000000" => rgb <= "000000";
					when "00101001000000001" => rgb <= "000000";
					when "00101001000000010" => rgb <= "000000";
					when "00101001000000011" => rgb <= "000000";
					when "00101001000000100" => rgb <= "000000";
					when "00101001000000101" => rgb <= "000000";
					when "00101001000000110" => rgb <= "000000";
					when "00101001000000111" => rgb <= "000000";
					when "00101001000001000" => rgb <= "000000";
					when "00101001000001001" => rgb <= "000000";
					when "00101001000001010" => rgb <= "000000";
					when "00101001000001011" => rgb <= "000000";
					when "00101001000001100" => rgb <= "000000";
					when "00101001000001101" => rgb <= "000000";
					when "00101001000001110" => rgb <= "000000";
					when "00101001000001111" => rgb <= "000000";
					when "00101001000010000" => rgb <= "000000";
					when "00101001000010001" => rgb <= "000000";
					when "00101001000010010" => rgb <= "000000";
					when "00101001000010011" => rgb <= "000000";
					when "00101001000010100" => rgb <= "000000";
					when "00101001000010101" => rgb <= "000000";
					when "00101001000010110" => rgb <= "000000";
					when "00101001000010111" => rgb <= "000000";
					when "00101001000011000" => rgb <= "000000";
					when "00101001000011001" => rgb <= "000000";
					when "00101001000011010" => rgb <= "000000";
					when "00101001000011011" => rgb <= "000000";
					when "00101001000011100" => rgb <= "000000";
					when "00101001000011101" => rgb <= "000000";
					when "00101001000011110" => rgb <= "000000";
					when "00101001000011111" => rgb <= "000000";
					when "00101001000100000" => rgb <= "000000";
					when "00101001000100001" => rgb <= "000000";
					when "00101001000100010" => rgb <= "000000";
					when "00101001000100011" => rgb <= "000000";
					when "00101001000100100" => rgb <= "000000";
					when "00101001000100101" => rgb <= "000000";
					when "00101001000100110" => rgb <= "000000";
					when "00101001000100111" => rgb <= "000000";
					when "00101001000101000" => rgb <= "000000";
					when "00101001000101001" => rgb <= "000000";
					when "00101001000101010" => rgb <= "000000";
					when "00101001000101011" => rgb <= "000000";
					when "00101001000101100" => rgb <= "000000";
					when "00101001000101101" => rgb <= "000000";
					when "00101001000101110" => rgb <= "000000";
					when "00101001000101111" => rgb <= "000000";
					when "00101001000110000" => rgb <= "000000";
					when "00101001000110001" => rgb <= "000000";
					when "00101001000110010" => rgb <= "000000";
					when "00101001000110011" => rgb <= "000000";
					when "00101001000110100" => rgb <= "000000";
					when "00101001000110101" => rgb <= "000000";
					when "00101001000110110" => rgb <= "000000";
					when "00101001000110111" => rgb <= "000000";
					when "00101001000111000" => rgb <= "000000";
					when "00101001000111001" => rgb <= "000000";
					when "00101001000111010" => rgb <= "000000";
					when "00101001000111011" => rgb <= "000000";
					when "00101001000111100" => rgb <= "000000";
					when "00101001000111101" => rgb <= "000000";
					when "00101001000111110" => rgb <= "000000";
					when "00101001000111111" => rgb <= "000000";
					when "00101001001000000" => rgb <= "000000";
					when "00101001001000001" => rgb <= "000000";
					when "00101001001000010" => rgb <= "000000";
					when "00101001001000011" => rgb <= "000000";
					when "00101001001000100" => rgb <= "000000";
					when "00101001001000101" => rgb <= "000000";
					when "00101001001000110" => rgb <= "000000";
					when "00101001001000111" => rgb <= "000000";
					when "00101001001001000" => rgb <= "000000";
					when "00101001001001001" => rgb <= "000000";
					when "00101001001001010" => rgb <= "000000";
					when "00101001001001011" => rgb <= "000000";
					when "00101001001001100" => rgb <= "000000";
					when "00101001001001101" => rgb <= "000000";
					when "00101001001001110" => rgb <= "000000";
					when "00101001001001111" => rgb <= "000000";
					when "00101001001010000" => rgb <= "000000";
					when "00101001001010001" => rgb <= "000000";
					when "00101001001010010" => rgb <= "000000";
					when "00101001001010011" => rgb <= "000000";
					when "00101001001010100" => rgb <= "000000";
					when "00101001001010101" => rgb <= "000000";
					when "00101001001010110" => rgb <= "000000";
					when "00101001001010111" => rgb <= "000000";
					when "00101001001011000" => rgb <= "000000";
					when "00101001001011001" => rgb <= "000000";
					when "00101001001011010" => rgb <= "000000";
					when "00101001001011011" => rgb <= "000000";
					when "00101001001011100" => rgb <= "000000";
					when "00101001001011101" => rgb <= "000000";
					when "00101001001011110" => rgb <= "000000";
					when "00101001001011111" => rgb <= "000000";
					when "00101001001100000" => rgb <= "000000";
					when "00101001001100001" => rgb <= "000000";
					when "00101001001100010" => rgb <= "000000";
					when "00101001001100011" => rgb <= "000000";
					when "00101001001100100" => rgb <= "000000";
					when "00101001001100101" => rgb <= "000000";
					when "00101001001100110" => rgb <= "010100";
					when "00101001001100111" => rgb <= "111000";
					when "00101001001101000" => rgb <= "101000";
					when "00101001001101001" => rgb <= "101000";
					when "00101001001101010" => rgb <= "101000";
					when "00101001001101011" => rgb <= "101000";
					when "00101001001101100" => rgb <= "101000";
					when "00101001001101101" => rgb <= "101000";
					when "00101001001101110" => rgb <= "101000";
					when "00101001001101111" => rgb <= "101000";
					when "00101001001110000" => rgb <= "101000";
					when "00101001001110001" => rgb <= "101000";
					when "00101001001110010" => rgb <= "101000";
					when "00101001001110011" => rgb <= "101000";
					when "00101001001110100" => rgb <= "101000";
					when "00101001001110101" => rgb <= "101000";
					when "00101001001110110" => rgb <= "101000";
					when "00101001001110111" => rgb <= "101000";
					when "00101001001111000" => rgb <= "101000";
					when "00101001001111001" => rgb <= "101000";
					when "00101001001111010" => rgb <= "101000";
					when "00101001001111011" => rgb <= "101000";
					when "00101001001111100" => rgb <= "101000";
					when "00101001001111101" => rgb <= "101000";
					when "00101001001111110" => rgb <= "101000";
					when "00101001001111111" => rgb <= "101000";
					when "00101001010000000" => rgb <= "101000";
					when "00101001010000001" => rgb <= "101000";
					when "00101001010000010" => rgb <= "101000";
					when "00101001010000011" => rgb <= "101000";
					when "00101001010000100" => rgb <= "101000";
					when "00101001010000101" => rgb <= "101000";
					when "00101001010000110" => rgb <= "101000";
					when "00101001010000111" => rgb <= "101000";
					when "00101001010001000" => rgb <= "101001";
					when "00101001010001001" => rgb <= "111001";
					when "00101001010001010" => rgb <= "101001";
					when "00101001010001011" => rgb <= "101001";
					when "00101001010001100" => rgb <= "111001";
					when "00101001010001101" => rgb <= "111001";
					when "00101001010001110" => rgb <= "111001";
					when "00101001010001111" => rgb <= "101001";
					when "00101001010010000" => rgb <= "111001";
					when "00101001010010001" => rgb <= "101001";
					when "00101001010010010" => rgb <= "111001";
					when "00101001010010011" => rgb <= "101001";
					when "00101001010010100" => rgb <= "101000";
					when "00101001010010101" => rgb <= "101000";
					when "00101001010010110" => rgb <= "101000";
					when "00101001010010111" => rgb <= "101000";
					when "00101001010011000" => rgb <= "101000";
					when "00101001010011001" => rgb <= "101000";
					when "00101001010011010" => rgb <= "101000";
					when "00101001010011011" => rgb <= "101000";
					when "00101001010011100" => rgb <= "101000";
					when "00101001010011101" => rgb <= "101000";
					when "00101001010011110" => rgb <= "101000";
					when "00101001010011111" => rgb <= "101000";
					when "00101001010100000" => rgb <= "101000";
					when "00101001010100001" => rgb <= "101000";
					when "00101001010100010" => rgb <= "101000";
					when "00101001010100011" => rgb <= "101000";
					when "00101001010100100" => rgb <= "101000";
					when "00101001010100101" => rgb <= "101000";
					when "00101001010100110" => rgb <= "101000";
					when "00101001010100111" => rgb <= "101000";
					when "00101001010101000" => rgb <= "101000";
					when "00101001010101001" => rgb <= "101000";
					when "00101001010101010" => rgb <= "101000";
					when "00101001010101011" => rgb <= "101000";
					when "00101001010101100" => rgb <= "101000";
					when "00101001010101101" => rgb <= "101000";
					when "00101001010101110" => rgb <= "101000";
					when "00101001010101111" => rgb <= "101000";
					when "00101001010110000" => rgb <= "101000";
					when "00101001010110001" => rgb <= "101000";
					when "00101001010110010" => rgb <= "101000";
					when "00101001010110011" => rgb <= "101000";
					when "00101001010110100" => rgb <= "101000";
					when "00101001010110101" => rgb <= "101000";
					when "00101001010110110" => rgb <= "101000";
					when "00101001010110111" => rgb <= "101000";
					when "00101001010111000" => rgb <= "101000";
					when "00101001010111001" => rgb <= "101000";
					when "00101001010111010" => rgb <= "101000";
					when "00101001010111011" => rgb <= "101000";
					when "00101001010111100" => rgb <= "101000";
					when "00101001010111101" => rgb <= "101000";
					when "00101001010111110" => rgb <= "101000";
					when "00101001010111111" => rgb <= "101000";
					when "00101001011000000" => rgb <= "101000";
					when "00101001011000001" => rgb <= "101000";
					when "00101001011000010" => rgb <= "101000";
					when "00101001011000011" => rgb <= "101000";
					when "00101001011000100" => rgb <= "101000";
					when "00101001011000101" => rgb <= "101000";
					when "00101001011000110" => rgb <= "101000";
					when "00101001011000111" => rgb <= "101000";
					when "00101001011001000" => rgb <= "101000";
					when "00101001011001001" => rgb <= "101000";
					when "00101001011001010" => rgb <= "101000";
					when "00101001011001011" => rgb <= "101000";
					when "00101001011001100" => rgb <= "101000";
					when "00101001011001101" => rgb <= "101000";
					when "00101001011001110" => rgb <= "101000";
					when "00101001011001111" => rgb <= "101000";
					when "00101001011010000" => rgb <= "101000";
					when "00101001011010001" => rgb <= "101000";
					when "00101001011010010" => rgb <= "101000";
					when "00101001011010011" => rgb <= "101000";
					when "00101001011010100" => rgb <= "101000";
					when "00101001011010101" => rgb <= "101000";
					when "00101001011010110" => rgb <= "101000";
					when "00101001011010111" => rgb <= "010100";
					when "00101001011011000" => rgb <= "000000";
					when "00101001011011001" => rgb <= "000000";
					when "00101001011011010" => rgb <= "000000";
					when "00101001011011011" => rgb <= "000000";
					when "00101001011011100" => rgb <= "000000";
					when "00101001011011101" => rgb <= "000000";
					when "00101001011011110" => rgb <= "000000";
					when "00101001011011111" => rgb <= "000000";
					when "00101001011100000" => rgb <= "000000";
					when "00101001011100001" => rgb <= "000000";
					when "00101001011100010" => rgb <= "000000";
					when "00101001011100011" => rgb <= "000000";
					when "00101001011100100" => rgb <= "000000";
					when "00101001011100101" => rgb <= "000000";
					when "00101001011100110" => rgb <= "000000";
					when "00101001011100111" => rgb <= "000000";
					when "00101001011101000" => rgb <= "000000";
					when "00101001011101001" => rgb <= "000000";
					when "00101001011101010" => rgb <= "000000";
					when "00101001011101011" => rgb <= "000000";
					when "00101001011101100" => rgb <= "000000";
					when "00101001011101101" => rgb <= "000000";
					when "00101001011101110" => rgb <= "000000";
					when "00101001011101111" => rgb <= "000000";
					when "00101001011110000" => rgb <= "000000";
					when "00101001011110001" => rgb <= "000000";
					when "00101001011110010" => rgb <= "000000";
					when "00101001011110011" => rgb <= "000000";
					when "00101001011110100" => rgb <= "000000";
					when "00101001011110101" => rgb <= "000000";
					when "00101001011110110" => rgb <= "000000";
					when "00101001011110111" => rgb <= "000000";
					when "00101001011111000" => rgb <= "000000";
					when "00101001011111001" => rgb <= "000000";
					when "00101001011111010" => rgb <= "000000";
					when "00101001011111011" => rgb <= "000000";
					when "00101001011111100" => rgb <= "000000";
					when "00101001011111101" => rgb <= "000000";
					when "00101001011111110" => rgb <= "000000";
					when "00101001011111111" => rgb <= "000000";
					when "00101001100000000" => rgb <= "000000";
					when "00101001100000001" => rgb <= "000000";
					when "00101001100000010" => rgb <= "000000";
					when "00101001100000011" => rgb <= "000000";
					when "00101001100000100" => rgb <= "000000";
					when "00101001100000101" => rgb <= "000000";
					when "00101001100000110" => rgb <= "000000";
					when "00101001100000111" => rgb <= "000000";
					when "00101001100001000" => rgb <= "000000";
					when "00101001100001001" => rgb <= "000000";
					when "00101001100001010" => rgb <= "000000";
					when "00101001100001011" => rgb <= "000000";
					when "00101001100001100" => rgb <= "000000";
					when "00101001100001101" => rgb <= "000000";
					when "00101001100001110" => rgb <= "000000";
					when "00101001100001111" => rgb <= "000000";
					when "00101001100010000" => rgb <= "000000";
					when "00101001100010001" => rgb <= "000000";
					when "00101001100010010" => rgb <= "000000";
					when "00101001100010011" => rgb <= "000000";
					when "00101001100010100" => rgb <= "000000";
					when "00101001100010101" => rgb <= "000000";
					when "00101001100010110" => rgb <= "000000";
					when "00101001100010111" => rgb <= "000000";
					when "00101001100011000" => rgb <= "000000";
					when "00101001100011001" => rgb <= "000000";
					when "00101001100011010" => rgb <= "000000";
					when "00101001100011011" => rgb <= "000000";
					when "00101001100011100" => rgb <= "000000";
					when "00101001100011101" => rgb <= "000000";
					when "00101001100011110" => rgb <= "000000";
					when "00101001100011111" => rgb <= "000000";
					when "00101001100100000" => rgb <= "000000";
					when "00101001100100001" => rgb <= "000000";
					when "00101001100100010" => rgb <= "000000";
					when "00101001100100011" => rgb <= "000000";
					when "00101001100100100" => rgb <= "000000";
					when "00101001100100101" => rgb <= "000000";
					when "00101001100100110" => rgb <= "000000";
					when "00101001100100111" => rgb <= "000000";
					when "00101001100101000" => rgb <= "000000";
					when "00101001100101001" => rgb <= "000000";
					when "00101001100101010" => rgb <= "000000";
					when "00101001100101011" => rgb <= "000000";
					when "00101001100101100" => rgb <= "000000";
					when "00101001100101101" => rgb <= "000000";
					when "00101001100101110" => rgb <= "000000";
					when "00101001100101111" => rgb <= "000000";
					when "00101001100110000" => rgb <= "000000";
					when "00101001100110001" => rgb <= "000000";
					when "00101001100110010" => rgb <= "000000";
					when "00101001100110011" => rgb <= "000000";
					when "00101001100110100" => rgb <= "000000";
					when "00101001100110101" => rgb <= "000000";
					when "00101001100110110" => rgb <= "000000";
					when "00101001100110111" => rgb <= "000000";
					when "00101001100111000" => rgb <= "000000";
					when "00101001100111001" => rgb <= "000000";
					when "00101001100111010" => rgb <= "000000";
					when "00101001100111011" => rgb <= "000000";
					when "00101001100111100" => rgb <= "000000";
					when "00101001100111101" => rgb <= "000000";
					when "00101001100111110" => rgb <= "000000";
					when "00101001100111111" => rgb <= "000000";
					when "00101010000000000" => rgb <= "000000";
					when "00101010000000001" => rgb <= "000000";
					when "00101010000000010" => rgb <= "000000";
					when "00101010000000011" => rgb <= "000000";
					when "00101010000000100" => rgb <= "000000";
					when "00101010000000101" => rgb <= "000000";
					when "00101010000000110" => rgb <= "000000";
					when "00101010000000111" => rgb <= "000000";
					when "00101010000001000" => rgb <= "000000";
					when "00101010000001001" => rgb <= "000000";
					when "00101010000001010" => rgb <= "000000";
					when "00101010000001011" => rgb <= "000000";
					when "00101010000001100" => rgb <= "000000";
					when "00101010000001101" => rgb <= "000000";
					when "00101010000001110" => rgb <= "000000";
					when "00101010000001111" => rgb <= "000000";
					when "00101010000010000" => rgb <= "000000";
					when "00101010000010001" => rgb <= "000000";
					when "00101010000010010" => rgb <= "000000";
					when "00101010000010011" => rgb <= "000000";
					when "00101010000010100" => rgb <= "000000";
					when "00101010000010101" => rgb <= "000000";
					when "00101010000010110" => rgb <= "000000";
					when "00101010000010111" => rgb <= "000000";
					when "00101010000011000" => rgb <= "000000";
					when "00101010000011001" => rgb <= "000000";
					when "00101010000011010" => rgb <= "000000";
					when "00101010000011011" => rgb <= "000000";
					when "00101010000011100" => rgb <= "000000";
					when "00101010000011101" => rgb <= "000000";
					when "00101010000011110" => rgb <= "000000";
					when "00101010000011111" => rgb <= "000000";
					when "00101010000100000" => rgb <= "000000";
					when "00101010000100001" => rgb <= "000000";
					when "00101010000100010" => rgb <= "000000";
					when "00101010000100011" => rgb <= "000000";
					when "00101010000100100" => rgb <= "000000";
					when "00101010000100101" => rgb <= "000000";
					when "00101010000100110" => rgb <= "000000";
					when "00101010000100111" => rgb <= "000000";
					when "00101010000101000" => rgb <= "000000";
					when "00101010000101001" => rgb <= "000000";
					when "00101010000101010" => rgb <= "000000";
					when "00101010000101011" => rgb <= "000000";
					when "00101010000101100" => rgb <= "000000";
					when "00101010000101101" => rgb <= "000000";
					when "00101010000101110" => rgb <= "000000";
					when "00101010000101111" => rgb <= "000000";
					when "00101010000110000" => rgb <= "000000";
					when "00101010000110001" => rgb <= "000000";
					when "00101010000110010" => rgb <= "000000";
					when "00101010000110011" => rgb <= "000000";
					when "00101010000110100" => rgb <= "000000";
					when "00101010000110101" => rgb <= "000000";
					when "00101010000110110" => rgb <= "000000";
					when "00101010000110111" => rgb <= "000000";
					when "00101010000111000" => rgb <= "000000";
					when "00101010000111001" => rgb <= "000000";
					when "00101010000111010" => rgb <= "000000";
					when "00101010000111011" => rgb <= "000000";
					when "00101010000111100" => rgb <= "000000";
					when "00101010000111101" => rgb <= "000000";
					when "00101010000111110" => rgb <= "000000";
					when "00101010000111111" => rgb <= "000000";
					when "00101010001000000" => rgb <= "000000";
					when "00101010001000001" => rgb <= "000000";
					when "00101010001000010" => rgb <= "000000";
					when "00101010001000011" => rgb <= "000000";
					when "00101010001000100" => rgb <= "000000";
					when "00101010001000101" => rgb <= "000000";
					when "00101010001000110" => rgb <= "000000";
					when "00101010001000111" => rgb <= "000000";
					when "00101010001001000" => rgb <= "000000";
					when "00101010001001001" => rgb <= "000000";
					when "00101010001001010" => rgb <= "000000";
					when "00101010001001011" => rgb <= "000000";
					when "00101010001001100" => rgb <= "000000";
					when "00101010001001101" => rgb <= "000000";
					when "00101010001001110" => rgb <= "000000";
					when "00101010001001111" => rgb <= "000000";
					when "00101010001010000" => rgb <= "000000";
					when "00101010001010001" => rgb <= "000000";
					when "00101010001010010" => rgb <= "000000";
					when "00101010001010011" => rgb <= "000000";
					when "00101010001010100" => rgb <= "000000";
					when "00101010001010101" => rgb <= "000000";
					when "00101010001010110" => rgb <= "000000";
					when "00101010001010111" => rgb <= "000000";
					when "00101010001011000" => rgb <= "000000";
					when "00101010001011001" => rgb <= "000000";
					when "00101010001011010" => rgb <= "000000";
					when "00101010001011011" => rgb <= "000000";
					when "00101010001011100" => rgb <= "000000";
					when "00101010001011101" => rgb <= "000000";
					when "00101010001011110" => rgb <= "000000";
					when "00101010001011111" => rgb <= "000000";
					when "00101010001100000" => rgb <= "000000";
					when "00101010001100001" => rgb <= "000000";
					when "00101010001100010" => rgb <= "000000";
					when "00101010001100011" => rgb <= "000000";
					when "00101010001100100" => rgb <= "000000";
					when "00101010001100101" => rgb <= "000000";
					when "00101010001100110" => rgb <= "010100";
					when "00101010001100111" => rgb <= "111000";
					when "00101010001101000" => rgb <= "101000";
					when "00101010001101001" => rgb <= "101000";
					when "00101010001101010" => rgb <= "101000";
					when "00101010001101011" => rgb <= "101000";
					when "00101010001101100" => rgb <= "101000";
					when "00101010001101101" => rgb <= "101000";
					when "00101010001101110" => rgb <= "101000";
					when "00101010001101111" => rgb <= "101000";
					when "00101010001110000" => rgb <= "101000";
					when "00101010001110001" => rgb <= "101000";
					when "00101010001110010" => rgb <= "101000";
					when "00101010001110011" => rgb <= "101000";
					when "00101010001110100" => rgb <= "101000";
					when "00101010001110101" => rgb <= "101000";
					when "00101010001110110" => rgb <= "101000";
					when "00101010001110111" => rgb <= "101000";
					when "00101010001111000" => rgb <= "101000";
					when "00101010001111001" => rgb <= "101000";
					when "00101010001111010" => rgb <= "101000";
					when "00101010001111011" => rgb <= "101000";
					when "00101010001111100" => rgb <= "101000";
					when "00101010001111101" => rgb <= "101000";
					when "00101010001111110" => rgb <= "101000";
					when "00101010001111111" => rgb <= "101000";
					when "00101010010000000" => rgb <= "101000";
					when "00101010010000001" => rgb <= "101000";
					when "00101010010000010" => rgb <= "101000";
					when "00101010010000011" => rgb <= "101000";
					when "00101010010000100" => rgb <= "101000";
					when "00101010010000101" => rgb <= "101000";
					when "00101010010000110" => rgb <= "101000";
					when "00101010010000111" => rgb <= "101000";
					when "00101010010001000" => rgb <= "101001";
					when "00101010010001001" => rgb <= "111001";
					when "00101010010001010" => rgb <= "101001";
					when "00101010010001011" => rgb <= "101001";
					when "00101010010001100" => rgb <= "111001";
					when "00101010010001101" => rgb <= "111001";
					when "00101010010001110" => rgb <= "111001";
					when "00101010010001111" => rgb <= "101001";
					when "00101010010010000" => rgb <= "111001";
					when "00101010010010001" => rgb <= "101001";
					when "00101010010010010" => rgb <= "111001";
					when "00101010010010011" => rgb <= "101001";
					when "00101010010010100" => rgb <= "101000";
					when "00101010010010101" => rgb <= "101000";
					when "00101010010010110" => rgb <= "101000";
					when "00101010010010111" => rgb <= "101000";
					when "00101010010011000" => rgb <= "101000";
					when "00101010010011001" => rgb <= "101000";
					when "00101010010011010" => rgb <= "101000";
					when "00101010010011011" => rgb <= "101000";
					when "00101010010011100" => rgb <= "101000";
					when "00101010010011101" => rgb <= "101000";
					when "00101010010011110" => rgb <= "101000";
					when "00101010010011111" => rgb <= "101000";
					when "00101010010100000" => rgb <= "101000";
					when "00101010010100001" => rgb <= "101000";
					when "00101010010100010" => rgb <= "101000";
					when "00101010010100011" => rgb <= "101000";
					when "00101010010100100" => rgb <= "101000";
					when "00101010010100101" => rgb <= "101000";
					when "00101010010100110" => rgb <= "101000";
					when "00101010010100111" => rgb <= "101000";
					when "00101010010101000" => rgb <= "101000";
					when "00101010010101001" => rgb <= "101000";
					when "00101010010101010" => rgb <= "101000";
					when "00101010010101011" => rgb <= "101000";
					when "00101010010101100" => rgb <= "101000";
					when "00101010010101101" => rgb <= "101000";
					when "00101010010101110" => rgb <= "101000";
					when "00101010010101111" => rgb <= "101000";
					when "00101010010110000" => rgb <= "101000";
					when "00101010010110001" => rgb <= "101000";
					when "00101010010110010" => rgb <= "101000";
					when "00101010010110011" => rgb <= "101000";
					when "00101010010110100" => rgb <= "101000";
					when "00101010010110101" => rgb <= "101000";
					when "00101010010110110" => rgb <= "101000";
					when "00101010010110111" => rgb <= "101000";
					when "00101010010111000" => rgb <= "101000";
					when "00101010010111001" => rgb <= "101000";
					when "00101010010111010" => rgb <= "101000";
					when "00101010010111011" => rgb <= "101000";
					when "00101010010111100" => rgb <= "101000";
					when "00101010010111101" => rgb <= "101000";
					when "00101010010111110" => rgb <= "101000";
					when "00101010010111111" => rgb <= "101000";
					when "00101010011000000" => rgb <= "101000";
					when "00101010011000001" => rgb <= "101000";
					when "00101010011000010" => rgb <= "101000";
					when "00101010011000011" => rgb <= "101000";
					when "00101010011000100" => rgb <= "101000";
					when "00101010011000101" => rgb <= "101000";
					when "00101010011000110" => rgb <= "101000";
					when "00101010011000111" => rgb <= "101000";
					when "00101010011001000" => rgb <= "101000";
					when "00101010011001001" => rgb <= "101000";
					when "00101010011001010" => rgb <= "101000";
					when "00101010011001011" => rgb <= "101000";
					when "00101010011001100" => rgb <= "101000";
					when "00101010011001101" => rgb <= "101000";
					when "00101010011001110" => rgb <= "101000";
					when "00101010011001111" => rgb <= "101000";
					when "00101010011010000" => rgb <= "101000";
					when "00101010011010001" => rgb <= "101000";
					when "00101010011010010" => rgb <= "101000";
					when "00101010011010011" => rgb <= "101000";
					when "00101010011010100" => rgb <= "101000";
					when "00101010011010101" => rgb <= "101000";
					when "00101010011010110" => rgb <= "101000";
					when "00101010011010111" => rgb <= "010100";
					when "00101010011011000" => rgb <= "000000";
					when "00101010011011001" => rgb <= "000000";
					when "00101010011011010" => rgb <= "000000";
					when "00101010011011011" => rgb <= "000000";
					when "00101010011011100" => rgb <= "000000";
					when "00101010011011101" => rgb <= "000000";
					when "00101010011011110" => rgb <= "000000";
					when "00101010011011111" => rgb <= "000000";
					when "00101010011100000" => rgb <= "000000";
					when "00101010011100001" => rgb <= "000000";
					when "00101010011100010" => rgb <= "000000";
					when "00101010011100011" => rgb <= "000000";
					when "00101010011100100" => rgb <= "000000";
					when "00101010011100101" => rgb <= "000000";
					when "00101010011100110" => rgb <= "000000";
					when "00101010011100111" => rgb <= "000000";
					when "00101010011101000" => rgb <= "000000";
					when "00101010011101001" => rgb <= "000000";
					when "00101010011101010" => rgb <= "000000";
					when "00101010011101011" => rgb <= "000000";
					when "00101010011101100" => rgb <= "000000";
					when "00101010011101101" => rgb <= "000000";
					when "00101010011101110" => rgb <= "000000";
					when "00101010011101111" => rgb <= "000000";
					when "00101010011110000" => rgb <= "000000";
					when "00101010011110001" => rgb <= "000000";
					when "00101010011110010" => rgb <= "000000";
					when "00101010011110011" => rgb <= "000000";
					when "00101010011110100" => rgb <= "000000";
					when "00101010011110101" => rgb <= "000000";
					when "00101010011110110" => rgb <= "000000";
					when "00101010011110111" => rgb <= "000000";
					when "00101010011111000" => rgb <= "000000";
					when "00101010011111001" => rgb <= "000000";
					when "00101010011111010" => rgb <= "000000";
					when "00101010011111011" => rgb <= "000000";
					when "00101010011111100" => rgb <= "000000";
					when "00101010011111101" => rgb <= "000000";
					when "00101010011111110" => rgb <= "000000";
					when "00101010011111111" => rgb <= "000000";
					when "00101010100000000" => rgb <= "000000";
					when "00101010100000001" => rgb <= "000000";
					when "00101010100000010" => rgb <= "000000";
					when "00101010100000011" => rgb <= "000000";
					when "00101010100000100" => rgb <= "000000";
					when "00101010100000101" => rgb <= "000000";
					when "00101010100000110" => rgb <= "000000";
					when "00101010100000111" => rgb <= "000000";
					when "00101010100001000" => rgb <= "000000";
					when "00101010100001001" => rgb <= "000000";
					when "00101010100001010" => rgb <= "000000";
					when "00101010100001011" => rgb <= "000000";
					when "00101010100001100" => rgb <= "000000";
					when "00101010100001101" => rgb <= "000000";
					when "00101010100001110" => rgb <= "000000";
					when "00101010100001111" => rgb <= "000000";
					when "00101010100010000" => rgb <= "000000";
					when "00101010100010001" => rgb <= "000000";
					when "00101010100010010" => rgb <= "000000";
					when "00101010100010011" => rgb <= "000000";
					when "00101010100010100" => rgb <= "000000";
					when "00101010100010101" => rgb <= "000000";
					when "00101010100010110" => rgb <= "000000";
					when "00101010100010111" => rgb <= "000000";
					when "00101010100011000" => rgb <= "000000";
					when "00101010100011001" => rgb <= "000000";
					when "00101010100011010" => rgb <= "000000";
					when "00101010100011011" => rgb <= "000000";
					when "00101010100011100" => rgb <= "000000";
					when "00101010100011101" => rgb <= "000000";
					when "00101010100011110" => rgb <= "000000";
					when "00101010100011111" => rgb <= "000000";
					when "00101010100100000" => rgb <= "000000";
					when "00101010100100001" => rgb <= "000000";
					when "00101010100100010" => rgb <= "000000";
					when "00101010100100011" => rgb <= "000000";
					when "00101010100100100" => rgb <= "000000";
					when "00101010100100101" => rgb <= "000000";
					when "00101010100100110" => rgb <= "000000";
					when "00101010100100111" => rgb <= "000000";
					when "00101010100101000" => rgb <= "000000";
					when "00101010100101001" => rgb <= "000000";
					when "00101010100101010" => rgb <= "000000";
					when "00101010100101011" => rgb <= "000000";
					when "00101010100101100" => rgb <= "000000";
					when "00101010100101101" => rgb <= "000000";
					when "00101010100101110" => rgb <= "000000";
					when "00101010100101111" => rgb <= "000000";
					when "00101010100110000" => rgb <= "000000";
					when "00101010100110001" => rgb <= "000000";
					when "00101010100110010" => rgb <= "000000";
					when "00101010100110011" => rgb <= "000000";
					when "00101010100110100" => rgb <= "000000";
					when "00101010100110101" => rgb <= "000000";
					when "00101010100110110" => rgb <= "000000";
					when "00101010100110111" => rgb <= "000000";
					when "00101010100111000" => rgb <= "000000";
					when "00101010100111001" => rgb <= "000000";
					when "00101010100111010" => rgb <= "000000";
					when "00101010100111011" => rgb <= "000000";
					when "00101010100111100" => rgb <= "000000";
					when "00101010100111101" => rgb <= "000000";
					when "00101010100111110" => rgb <= "000000";
					when "00101010100111111" => rgb <= "000000";
					when "00101011000000000" => rgb <= "000000";
					when "00101011000000001" => rgb <= "000000";
					when "00101011000000010" => rgb <= "000000";
					when "00101011000000011" => rgb <= "000000";
					when "00101011000000100" => rgb <= "000000";
					when "00101011000000101" => rgb <= "000000";
					when "00101011000000110" => rgb <= "000000";
					when "00101011000000111" => rgb <= "000000";
					when "00101011000001000" => rgb <= "000000";
					when "00101011000001001" => rgb <= "000000";
					when "00101011000001010" => rgb <= "000000";
					when "00101011000001011" => rgb <= "000000";
					when "00101011000001100" => rgb <= "000000";
					when "00101011000001101" => rgb <= "000000";
					when "00101011000001110" => rgb <= "000000";
					when "00101011000001111" => rgb <= "000000";
					when "00101011000010000" => rgb <= "000000";
					when "00101011000010001" => rgb <= "000000";
					when "00101011000010010" => rgb <= "000000";
					when "00101011000010011" => rgb <= "000000";
					when "00101011000010100" => rgb <= "000000";
					when "00101011000010101" => rgb <= "000000";
					when "00101011000010110" => rgb <= "000000";
					when "00101011000010111" => rgb <= "000000";
					when "00101011000011000" => rgb <= "000000";
					when "00101011000011001" => rgb <= "000000";
					when "00101011000011010" => rgb <= "000000";
					when "00101011000011011" => rgb <= "000000";
					when "00101011000011100" => rgb <= "000000";
					when "00101011000011101" => rgb <= "000000";
					when "00101011000011110" => rgb <= "000000";
					when "00101011000011111" => rgb <= "000000";
					when "00101011000100000" => rgb <= "000000";
					when "00101011000100001" => rgb <= "000000";
					when "00101011000100010" => rgb <= "000000";
					when "00101011000100011" => rgb <= "000000";
					when "00101011000100100" => rgb <= "000000";
					when "00101011000100101" => rgb <= "000000";
					when "00101011000100110" => rgb <= "000000";
					when "00101011000100111" => rgb <= "000000";
					when "00101011000101000" => rgb <= "000000";
					when "00101011000101001" => rgb <= "000000";
					when "00101011000101010" => rgb <= "000000";
					when "00101011000101011" => rgb <= "000000";
					when "00101011000101100" => rgb <= "000000";
					when "00101011000101101" => rgb <= "000000";
					when "00101011000101110" => rgb <= "000000";
					when "00101011000101111" => rgb <= "000000";
					when "00101011000110000" => rgb <= "000000";
					when "00101011000110001" => rgb <= "000000";
					when "00101011000110010" => rgb <= "000000";
					when "00101011000110011" => rgb <= "000000";
					when "00101011000110100" => rgb <= "000000";
					when "00101011000110101" => rgb <= "000000";
					when "00101011000110110" => rgb <= "000000";
					when "00101011000110111" => rgb <= "000000";
					when "00101011000111000" => rgb <= "000000";
					when "00101011000111001" => rgb <= "000000";
					when "00101011000111010" => rgb <= "000000";
					when "00101011000111011" => rgb <= "000000";
					when "00101011000111100" => rgb <= "000000";
					when "00101011000111101" => rgb <= "000000";
					when "00101011000111110" => rgb <= "000000";
					when "00101011000111111" => rgb <= "000000";
					when "00101011001000000" => rgb <= "000000";
					when "00101011001000001" => rgb <= "000000";
					when "00101011001000010" => rgb <= "000000";
					when "00101011001000011" => rgb <= "000000";
					when "00101011001000100" => rgb <= "000000";
					when "00101011001000101" => rgb <= "000000";
					when "00101011001000110" => rgb <= "000000";
					when "00101011001000111" => rgb <= "000000";
					when "00101011001001000" => rgb <= "000000";
					when "00101011001001001" => rgb <= "000000";
					when "00101011001001010" => rgb <= "000000";
					when "00101011001001011" => rgb <= "000000";
					when "00101011001001100" => rgb <= "000000";
					when "00101011001001101" => rgb <= "000000";
					when "00101011001001110" => rgb <= "000000";
					when "00101011001001111" => rgb <= "000000";
					when "00101011001010000" => rgb <= "000000";
					when "00101011001010001" => rgb <= "000000";
					when "00101011001010010" => rgb <= "000000";
					when "00101011001010011" => rgb <= "000000";
					when "00101011001010100" => rgb <= "000000";
					when "00101011001010101" => rgb <= "000000";
					when "00101011001010110" => rgb <= "000000";
					when "00101011001010111" => rgb <= "000000";
					when "00101011001011000" => rgb <= "000000";
					when "00101011001011001" => rgb <= "000000";
					when "00101011001011010" => rgb <= "000000";
					when "00101011001011011" => rgb <= "000000";
					when "00101011001011100" => rgb <= "000000";
					when "00101011001011101" => rgb <= "000000";
					when "00101011001011110" => rgb <= "000000";
					when "00101011001011111" => rgb <= "000000";
					when "00101011001100000" => rgb <= "000000";
					when "00101011001100001" => rgb <= "000000";
					when "00101011001100010" => rgb <= "000000";
					when "00101011001100011" => rgb <= "000000";
					when "00101011001100100" => rgb <= "000000";
					when "00101011001100101" => rgb <= "000000";
					when "00101011001100110" => rgb <= "010100";
					when "00101011001100111" => rgb <= "111000";
					when "00101011001101000" => rgb <= "101000";
					when "00101011001101001" => rgb <= "101000";
					when "00101011001101010" => rgb <= "101000";
					when "00101011001101011" => rgb <= "101000";
					when "00101011001101100" => rgb <= "101000";
					when "00101011001101101" => rgb <= "101000";
					when "00101011001101110" => rgb <= "101000";
					when "00101011001101111" => rgb <= "101000";
					when "00101011001110000" => rgb <= "101000";
					when "00101011001110001" => rgb <= "101000";
					when "00101011001110010" => rgb <= "101000";
					when "00101011001110011" => rgb <= "101000";
					when "00101011001110100" => rgb <= "101000";
					when "00101011001110101" => rgb <= "101000";
					when "00101011001110110" => rgb <= "101000";
					when "00101011001110111" => rgb <= "101000";
					when "00101011001111000" => rgb <= "101000";
					when "00101011001111001" => rgb <= "101000";
					when "00101011001111010" => rgb <= "101000";
					when "00101011001111011" => rgb <= "101000";
					when "00101011001111100" => rgb <= "101000";
					when "00101011001111101" => rgb <= "101000";
					when "00101011001111110" => rgb <= "101000";
					when "00101011001111111" => rgb <= "101000";
					when "00101011010000000" => rgb <= "101000";
					when "00101011010000001" => rgb <= "101000";
					when "00101011010000010" => rgb <= "101000";
					when "00101011010000011" => rgb <= "101000";
					when "00101011010000100" => rgb <= "101000";
					when "00101011010000101" => rgb <= "101000";
					when "00101011010000110" => rgb <= "101000";
					when "00101011010000111" => rgb <= "101000";
					when "00101011010001000" => rgb <= "101001";
					when "00101011010001001" => rgb <= "111001";
					when "00101011010001010" => rgb <= "101001";
					when "00101011010001011" => rgb <= "101001";
					when "00101011010001100" => rgb <= "111001";
					when "00101011010001101" => rgb <= "111001";
					when "00101011010001110" => rgb <= "111001";
					when "00101011010001111" => rgb <= "101001";
					when "00101011010010000" => rgb <= "111001";
					when "00101011010010001" => rgb <= "101001";
					when "00101011010010010" => rgb <= "111001";
					when "00101011010010011" => rgb <= "101001";
					when "00101011010010100" => rgb <= "101000";
					when "00101011010010101" => rgb <= "101000";
					when "00101011010010110" => rgb <= "101000";
					when "00101011010010111" => rgb <= "101000";
					when "00101011010011000" => rgb <= "101000";
					when "00101011010011001" => rgb <= "101000";
					when "00101011010011010" => rgb <= "101000";
					when "00101011010011011" => rgb <= "101000";
					when "00101011010011100" => rgb <= "101000";
					when "00101011010011101" => rgb <= "101000";
					when "00101011010011110" => rgb <= "101000";
					when "00101011010011111" => rgb <= "101000";
					when "00101011010100000" => rgb <= "101000";
					when "00101011010100001" => rgb <= "101000";
					when "00101011010100010" => rgb <= "101000";
					when "00101011010100011" => rgb <= "101000";
					when "00101011010100100" => rgb <= "101000";
					when "00101011010100101" => rgb <= "101000";
					when "00101011010100110" => rgb <= "101000";
					when "00101011010100111" => rgb <= "101000";
					when "00101011010101000" => rgb <= "101000";
					when "00101011010101001" => rgb <= "101000";
					when "00101011010101010" => rgb <= "101000";
					when "00101011010101011" => rgb <= "101000";
					when "00101011010101100" => rgb <= "101000";
					when "00101011010101101" => rgb <= "101000";
					when "00101011010101110" => rgb <= "101000";
					when "00101011010101111" => rgb <= "101000";
					when "00101011010110000" => rgb <= "101000";
					when "00101011010110001" => rgb <= "101000";
					when "00101011010110010" => rgb <= "101000";
					when "00101011010110011" => rgb <= "101000";
					when "00101011010110100" => rgb <= "101000";
					when "00101011010110101" => rgb <= "101000";
					when "00101011010110110" => rgb <= "101000";
					when "00101011010110111" => rgb <= "101000";
					when "00101011010111000" => rgb <= "101000";
					when "00101011010111001" => rgb <= "101000";
					when "00101011010111010" => rgb <= "101000";
					when "00101011010111011" => rgb <= "101000";
					when "00101011010111100" => rgb <= "101000";
					when "00101011010111101" => rgb <= "101000";
					when "00101011010111110" => rgb <= "101000";
					when "00101011010111111" => rgb <= "101000";
					when "00101011011000000" => rgb <= "101000";
					when "00101011011000001" => rgb <= "101000";
					when "00101011011000010" => rgb <= "101000";
					when "00101011011000011" => rgb <= "101000";
					when "00101011011000100" => rgb <= "101000";
					when "00101011011000101" => rgb <= "101000";
					when "00101011011000110" => rgb <= "101000";
					when "00101011011000111" => rgb <= "101000";
					when "00101011011001000" => rgb <= "101000";
					when "00101011011001001" => rgb <= "101000";
					when "00101011011001010" => rgb <= "101000";
					when "00101011011001011" => rgb <= "101000";
					when "00101011011001100" => rgb <= "101000";
					when "00101011011001101" => rgb <= "101000";
					when "00101011011001110" => rgb <= "101000";
					when "00101011011001111" => rgb <= "101000";
					when "00101011011010000" => rgb <= "101000";
					when "00101011011010001" => rgb <= "101000";
					when "00101011011010010" => rgb <= "101000";
					when "00101011011010011" => rgb <= "101000";
					when "00101011011010100" => rgb <= "101000";
					when "00101011011010101" => rgb <= "101000";
					when "00101011011010110" => rgb <= "101000";
					when "00101011011010111" => rgb <= "010100";
					when "00101011011011000" => rgb <= "000000";
					when "00101011011011001" => rgb <= "000000";
					when "00101011011011010" => rgb <= "000000";
					when "00101011011011011" => rgb <= "000000";
					when "00101011011011100" => rgb <= "000000";
					when "00101011011011101" => rgb <= "000000";
					when "00101011011011110" => rgb <= "000000";
					when "00101011011011111" => rgb <= "000000";
					when "00101011011100000" => rgb <= "000000";
					when "00101011011100001" => rgb <= "000000";
					when "00101011011100010" => rgb <= "000000";
					when "00101011011100011" => rgb <= "000000";
					when "00101011011100100" => rgb <= "000000";
					when "00101011011100101" => rgb <= "000000";
					when "00101011011100110" => rgb <= "000000";
					when "00101011011100111" => rgb <= "000000";
					when "00101011011101000" => rgb <= "000000";
					when "00101011011101001" => rgb <= "000000";
					when "00101011011101010" => rgb <= "000000";
					when "00101011011101011" => rgb <= "000000";
					when "00101011011101100" => rgb <= "000000";
					when "00101011011101101" => rgb <= "000000";
					when "00101011011101110" => rgb <= "000000";
					when "00101011011101111" => rgb <= "000000";
					when "00101011011110000" => rgb <= "000000";
					when "00101011011110001" => rgb <= "000000";
					when "00101011011110010" => rgb <= "000000";
					when "00101011011110011" => rgb <= "000000";
					when "00101011011110100" => rgb <= "000000";
					when "00101011011110101" => rgb <= "000000";
					when "00101011011110110" => rgb <= "000000";
					when "00101011011110111" => rgb <= "000000";
					when "00101011011111000" => rgb <= "000000";
					when "00101011011111001" => rgb <= "000000";
					when "00101011011111010" => rgb <= "000000";
					when "00101011011111011" => rgb <= "000000";
					when "00101011011111100" => rgb <= "000000";
					when "00101011011111101" => rgb <= "000000";
					when "00101011011111110" => rgb <= "000000";
					when "00101011011111111" => rgb <= "000000";
					when "00101011100000000" => rgb <= "000000";
					when "00101011100000001" => rgb <= "000000";
					when "00101011100000010" => rgb <= "000000";
					when "00101011100000011" => rgb <= "000000";
					when "00101011100000100" => rgb <= "000000";
					when "00101011100000101" => rgb <= "000000";
					when "00101011100000110" => rgb <= "000000";
					when "00101011100000111" => rgb <= "000000";
					when "00101011100001000" => rgb <= "000000";
					when "00101011100001001" => rgb <= "000000";
					when "00101011100001010" => rgb <= "000000";
					when "00101011100001011" => rgb <= "000000";
					when "00101011100001100" => rgb <= "000000";
					when "00101011100001101" => rgb <= "000000";
					when "00101011100001110" => rgb <= "000000";
					when "00101011100001111" => rgb <= "000000";
					when "00101011100010000" => rgb <= "000000";
					when "00101011100010001" => rgb <= "000000";
					when "00101011100010010" => rgb <= "000000";
					when "00101011100010011" => rgb <= "000000";
					when "00101011100010100" => rgb <= "000000";
					when "00101011100010101" => rgb <= "000000";
					when "00101011100010110" => rgb <= "000000";
					when "00101011100010111" => rgb <= "000000";
					when "00101011100011000" => rgb <= "000000";
					when "00101011100011001" => rgb <= "000000";
					when "00101011100011010" => rgb <= "000000";
					when "00101011100011011" => rgb <= "000000";
					when "00101011100011100" => rgb <= "000000";
					when "00101011100011101" => rgb <= "000000";
					when "00101011100011110" => rgb <= "000000";
					when "00101011100011111" => rgb <= "000000";
					when "00101011100100000" => rgb <= "000000";
					when "00101011100100001" => rgb <= "000000";
					when "00101011100100010" => rgb <= "000000";
					when "00101011100100011" => rgb <= "000000";
					when "00101011100100100" => rgb <= "000000";
					when "00101011100100101" => rgb <= "000000";
					when "00101011100100110" => rgb <= "000000";
					when "00101011100100111" => rgb <= "000000";
					when "00101011100101000" => rgb <= "000000";
					when "00101011100101001" => rgb <= "000000";
					when "00101011100101010" => rgb <= "000000";
					when "00101011100101011" => rgb <= "000000";
					when "00101011100101100" => rgb <= "000000";
					when "00101011100101101" => rgb <= "000000";
					when "00101011100101110" => rgb <= "000000";
					when "00101011100101111" => rgb <= "000000";
					when "00101011100110000" => rgb <= "000000";
					when "00101011100110001" => rgb <= "000000";
					when "00101011100110010" => rgb <= "000000";
					when "00101011100110011" => rgb <= "000000";
					when "00101011100110100" => rgb <= "000000";
					when "00101011100110101" => rgb <= "000000";
					when "00101011100110110" => rgb <= "000000";
					when "00101011100110111" => rgb <= "000000";
					when "00101011100111000" => rgb <= "000000";
					when "00101011100111001" => rgb <= "000000";
					when "00101011100111010" => rgb <= "000000";
					when "00101011100111011" => rgb <= "000000";
					when "00101011100111100" => rgb <= "000000";
					when "00101011100111101" => rgb <= "000000";
					when "00101011100111110" => rgb <= "000000";
					when "00101011100111111" => rgb <= "000000";
					when "00101100000000000" => rgb <= "000000";
					when "00101100000000001" => rgb <= "000000";
					when "00101100000000010" => rgb <= "000000";
					when "00101100000000011" => rgb <= "000000";
					when "00101100000000100" => rgb <= "000000";
					when "00101100000000101" => rgb <= "000000";
					when "00101100000000110" => rgb <= "000000";
					when "00101100000000111" => rgb <= "000000";
					when "00101100000001000" => rgb <= "000000";
					when "00101100000001001" => rgb <= "000000";
					when "00101100000001010" => rgb <= "000000";
					when "00101100000001011" => rgb <= "000000";
					when "00101100000001100" => rgb <= "000000";
					when "00101100000001101" => rgb <= "000000";
					when "00101100000001110" => rgb <= "000000";
					when "00101100000001111" => rgb <= "000000";
					when "00101100000010000" => rgb <= "000000";
					when "00101100000010001" => rgb <= "000000";
					when "00101100000010010" => rgb <= "000000";
					when "00101100000010011" => rgb <= "000000";
					when "00101100000010100" => rgb <= "000000";
					when "00101100000010101" => rgb <= "000000";
					when "00101100000010110" => rgb <= "000000";
					when "00101100000010111" => rgb <= "000000";
					when "00101100000011000" => rgb <= "000000";
					when "00101100000011001" => rgb <= "000000";
					when "00101100000011010" => rgb <= "000000";
					when "00101100000011011" => rgb <= "000000";
					when "00101100000011100" => rgb <= "000000";
					when "00101100000011101" => rgb <= "000000";
					when "00101100000011110" => rgb <= "000000";
					when "00101100000011111" => rgb <= "000000";
					when "00101100000100000" => rgb <= "000000";
					when "00101100000100001" => rgb <= "000000";
					when "00101100000100010" => rgb <= "000000";
					when "00101100000100011" => rgb <= "000000";
					when "00101100000100100" => rgb <= "000000";
					when "00101100000100101" => rgb <= "000000";
					when "00101100000100110" => rgb <= "000000";
					when "00101100000100111" => rgb <= "000000";
					when "00101100000101000" => rgb <= "000000";
					when "00101100000101001" => rgb <= "000000";
					when "00101100000101010" => rgb <= "000000";
					when "00101100000101011" => rgb <= "000000";
					when "00101100000101100" => rgb <= "000000";
					when "00101100000101101" => rgb <= "000000";
					when "00101100000101110" => rgb <= "000000";
					when "00101100000101111" => rgb <= "000000";
					when "00101100000110000" => rgb <= "000000";
					when "00101100000110001" => rgb <= "000000";
					when "00101100000110010" => rgb <= "000000";
					when "00101100000110011" => rgb <= "000000";
					when "00101100000110100" => rgb <= "000000";
					when "00101100000110101" => rgb <= "000000";
					when "00101100000110110" => rgb <= "000000";
					when "00101100000110111" => rgb <= "000000";
					when "00101100000111000" => rgb <= "000000";
					when "00101100000111001" => rgb <= "000000";
					when "00101100000111010" => rgb <= "000000";
					when "00101100000111011" => rgb <= "000000";
					when "00101100000111100" => rgb <= "000000";
					when "00101100000111101" => rgb <= "000000";
					when "00101100000111110" => rgb <= "000000";
					when "00101100000111111" => rgb <= "000000";
					when "00101100001000000" => rgb <= "000000";
					when "00101100001000001" => rgb <= "000000";
					when "00101100001000010" => rgb <= "000000";
					when "00101100001000011" => rgb <= "000000";
					when "00101100001000100" => rgb <= "000000";
					when "00101100001000101" => rgb <= "000000";
					when "00101100001000110" => rgb <= "000000";
					when "00101100001000111" => rgb <= "000000";
					when "00101100001001000" => rgb <= "000000";
					when "00101100001001001" => rgb <= "000000";
					when "00101100001001010" => rgb <= "000000";
					when "00101100001001011" => rgb <= "000000";
					when "00101100001001100" => rgb <= "000000";
					when "00101100001001101" => rgb <= "000000";
					when "00101100001001110" => rgb <= "000000";
					when "00101100001001111" => rgb <= "000000";
					when "00101100001010000" => rgb <= "000000";
					when "00101100001010001" => rgb <= "000000";
					when "00101100001010010" => rgb <= "000000";
					when "00101100001010011" => rgb <= "000000";
					when "00101100001010100" => rgb <= "000000";
					when "00101100001010101" => rgb <= "000000";
					when "00101100001010110" => rgb <= "000000";
					when "00101100001010111" => rgb <= "000000";
					when "00101100001011000" => rgb <= "000000";
					when "00101100001011001" => rgb <= "000000";
					when "00101100001011010" => rgb <= "000000";
					when "00101100001011011" => rgb <= "000000";
					when "00101100001011100" => rgb <= "000000";
					when "00101100001011101" => rgb <= "000000";
					when "00101100001011110" => rgb <= "000000";
					when "00101100001011111" => rgb <= "000000";
					when "00101100001100000" => rgb <= "000000";
					when "00101100001100001" => rgb <= "000000";
					when "00101100001100010" => rgb <= "000000";
					when "00101100001100011" => rgb <= "000000";
					when "00101100001100100" => rgb <= "000000";
					when "00101100001100101" => rgb <= "000000";
					when "00101100001100110" => rgb <= "010100";
					when "00101100001100111" => rgb <= "111000";
					when "00101100001101000" => rgb <= "101000";
					when "00101100001101001" => rgb <= "101000";
					when "00101100001101010" => rgb <= "101000";
					when "00101100001101011" => rgb <= "101000";
					when "00101100001101100" => rgb <= "101000";
					when "00101100001101101" => rgb <= "101000";
					when "00101100001101110" => rgb <= "101000";
					when "00101100001101111" => rgb <= "101000";
					when "00101100001110000" => rgb <= "101000";
					when "00101100001110001" => rgb <= "101000";
					when "00101100001110010" => rgb <= "101000";
					when "00101100001110011" => rgb <= "101000";
					when "00101100001110100" => rgb <= "101000";
					when "00101100001110101" => rgb <= "101000";
					when "00101100001110110" => rgb <= "101000";
					when "00101100001110111" => rgb <= "101000";
					when "00101100001111000" => rgb <= "101000";
					when "00101100001111001" => rgb <= "101000";
					when "00101100001111010" => rgb <= "101000";
					when "00101100001111011" => rgb <= "101000";
					when "00101100001111100" => rgb <= "101000";
					when "00101100001111101" => rgb <= "101000";
					when "00101100001111110" => rgb <= "101000";
					when "00101100001111111" => rgb <= "101000";
					when "00101100010000000" => rgb <= "101000";
					when "00101100010000001" => rgb <= "101000";
					when "00101100010000010" => rgb <= "101000";
					when "00101100010000011" => rgb <= "101000";
					when "00101100010000100" => rgb <= "101000";
					when "00101100010000101" => rgb <= "101000";
					when "00101100010000110" => rgb <= "101000";
					when "00101100010000111" => rgb <= "101000";
					when "00101100010001000" => rgb <= "101001";
					when "00101100010001001" => rgb <= "111001";
					when "00101100010001010" => rgb <= "101001";
					when "00101100010001011" => rgb <= "101001";
					when "00101100010001100" => rgb <= "111001";
					when "00101100010001101" => rgb <= "111001";
					when "00101100010001110" => rgb <= "111001";
					when "00101100010001111" => rgb <= "101001";
					when "00101100010010000" => rgb <= "111001";
					when "00101100010010001" => rgb <= "101001";
					when "00101100010010010" => rgb <= "111001";
					when "00101100010010011" => rgb <= "101001";
					when "00101100010010100" => rgb <= "101000";
					when "00101100010010101" => rgb <= "101000";
					when "00101100010010110" => rgb <= "101000";
					when "00101100010010111" => rgb <= "101000";
					when "00101100010011000" => rgb <= "101000";
					when "00101100010011001" => rgb <= "101000";
					when "00101100010011010" => rgb <= "101000";
					when "00101100010011011" => rgb <= "101000";
					when "00101100010011100" => rgb <= "101000";
					when "00101100010011101" => rgb <= "101000";
					when "00101100010011110" => rgb <= "101000";
					when "00101100010011111" => rgb <= "101000";
					when "00101100010100000" => rgb <= "101000";
					when "00101100010100001" => rgb <= "101000";
					when "00101100010100010" => rgb <= "101000";
					when "00101100010100011" => rgb <= "101000";
					when "00101100010100100" => rgb <= "101000";
					when "00101100010100101" => rgb <= "101000";
					when "00101100010100110" => rgb <= "101000";
					when "00101100010100111" => rgb <= "101000";
					when "00101100010101000" => rgb <= "101000";
					when "00101100010101001" => rgb <= "101000";
					when "00101100010101010" => rgb <= "101000";
					when "00101100010101011" => rgb <= "101000";
					when "00101100010101100" => rgb <= "101000";
					when "00101100010101101" => rgb <= "101000";
					when "00101100010101110" => rgb <= "101000";
					when "00101100010101111" => rgb <= "101000";
					when "00101100010110000" => rgb <= "101000";
					when "00101100010110001" => rgb <= "101000";
					when "00101100010110010" => rgb <= "101000";
					when "00101100010110011" => rgb <= "101000";
					when "00101100010110100" => rgb <= "101000";
					when "00101100010110101" => rgb <= "101000";
					when "00101100010110110" => rgb <= "101000";
					when "00101100010110111" => rgb <= "101000";
					when "00101100010111000" => rgb <= "101000";
					when "00101100010111001" => rgb <= "101000";
					when "00101100010111010" => rgb <= "101000";
					when "00101100010111011" => rgb <= "101000";
					when "00101100010111100" => rgb <= "101000";
					when "00101100010111101" => rgb <= "101000";
					when "00101100010111110" => rgb <= "101000";
					when "00101100010111111" => rgb <= "101000";
					when "00101100011000000" => rgb <= "101000";
					when "00101100011000001" => rgb <= "101000";
					when "00101100011000010" => rgb <= "101000";
					when "00101100011000011" => rgb <= "101000";
					when "00101100011000100" => rgb <= "101000";
					when "00101100011000101" => rgb <= "101000";
					when "00101100011000110" => rgb <= "101000";
					when "00101100011000111" => rgb <= "101000";
					when "00101100011001000" => rgb <= "101000";
					when "00101100011001001" => rgb <= "101000";
					when "00101100011001010" => rgb <= "101000";
					when "00101100011001011" => rgb <= "101000";
					when "00101100011001100" => rgb <= "101000";
					when "00101100011001101" => rgb <= "101000";
					when "00101100011001110" => rgb <= "101000";
					when "00101100011001111" => rgb <= "101000";
					when "00101100011010000" => rgb <= "101000";
					when "00101100011010001" => rgb <= "101000";
					when "00101100011010010" => rgb <= "101000";
					when "00101100011010011" => rgb <= "101000";
					when "00101100011010100" => rgb <= "101000";
					when "00101100011010101" => rgb <= "101000";
					when "00101100011010110" => rgb <= "101000";
					when "00101100011010111" => rgb <= "010100";
					when "00101100011011000" => rgb <= "000000";
					when "00101100011011001" => rgb <= "000000";
					when "00101100011011010" => rgb <= "000000";
					when "00101100011011011" => rgb <= "000000";
					when "00101100011011100" => rgb <= "000000";
					when "00101100011011101" => rgb <= "000000";
					when "00101100011011110" => rgb <= "000000";
					when "00101100011011111" => rgb <= "000000";
					when "00101100011100000" => rgb <= "000000";
					when "00101100011100001" => rgb <= "000000";
					when "00101100011100010" => rgb <= "000000";
					when "00101100011100011" => rgb <= "000000";
					when "00101100011100100" => rgb <= "000000";
					when "00101100011100101" => rgb <= "000000";
					when "00101100011100110" => rgb <= "000000";
					when "00101100011100111" => rgb <= "000000";
					when "00101100011101000" => rgb <= "000000";
					when "00101100011101001" => rgb <= "000000";
					when "00101100011101010" => rgb <= "000000";
					when "00101100011101011" => rgb <= "000000";
					when "00101100011101100" => rgb <= "000000";
					when "00101100011101101" => rgb <= "000000";
					when "00101100011101110" => rgb <= "000000";
					when "00101100011101111" => rgb <= "000000";
					when "00101100011110000" => rgb <= "000000";
					when "00101100011110001" => rgb <= "000000";
					when "00101100011110010" => rgb <= "000000";
					when "00101100011110011" => rgb <= "000000";
					when "00101100011110100" => rgb <= "000000";
					when "00101100011110101" => rgb <= "000000";
					when "00101100011110110" => rgb <= "000000";
					when "00101100011110111" => rgb <= "000000";
					when "00101100011111000" => rgb <= "000000";
					when "00101100011111001" => rgb <= "000000";
					when "00101100011111010" => rgb <= "000000";
					when "00101100011111011" => rgb <= "000000";
					when "00101100011111100" => rgb <= "000000";
					when "00101100011111101" => rgb <= "000000";
					when "00101100011111110" => rgb <= "000000";
					when "00101100011111111" => rgb <= "000000";
					when "00101100100000000" => rgb <= "000000";
					when "00101100100000001" => rgb <= "000000";
					when "00101100100000010" => rgb <= "000000";
					when "00101100100000011" => rgb <= "000000";
					when "00101100100000100" => rgb <= "000000";
					when "00101100100000101" => rgb <= "000000";
					when "00101100100000110" => rgb <= "000000";
					when "00101100100000111" => rgb <= "000000";
					when "00101100100001000" => rgb <= "000000";
					when "00101100100001001" => rgb <= "000000";
					when "00101100100001010" => rgb <= "000000";
					when "00101100100001011" => rgb <= "000000";
					when "00101100100001100" => rgb <= "000000";
					when "00101100100001101" => rgb <= "000000";
					when "00101100100001110" => rgb <= "000000";
					when "00101100100001111" => rgb <= "000000";
					when "00101100100010000" => rgb <= "000000";
					when "00101100100010001" => rgb <= "000000";
					when "00101100100010010" => rgb <= "000000";
					when "00101100100010011" => rgb <= "000000";
					when "00101100100010100" => rgb <= "000000";
					when "00101100100010101" => rgb <= "000000";
					when "00101100100010110" => rgb <= "000000";
					when "00101100100010111" => rgb <= "000000";
					when "00101100100011000" => rgb <= "000000";
					when "00101100100011001" => rgb <= "000000";
					when "00101100100011010" => rgb <= "000000";
					when "00101100100011011" => rgb <= "000000";
					when "00101100100011100" => rgb <= "000000";
					when "00101100100011101" => rgb <= "000000";
					when "00101100100011110" => rgb <= "000000";
					when "00101100100011111" => rgb <= "000000";
					when "00101100100100000" => rgb <= "000000";
					when "00101100100100001" => rgb <= "000000";
					when "00101100100100010" => rgb <= "000000";
					when "00101100100100011" => rgb <= "000000";
					when "00101100100100100" => rgb <= "000000";
					when "00101100100100101" => rgb <= "000000";
					when "00101100100100110" => rgb <= "000000";
					when "00101100100100111" => rgb <= "000000";
					when "00101100100101000" => rgb <= "000000";
					when "00101100100101001" => rgb <= "000000";
					when "00101100100101010" => rgb <= "000000";
					when "00101100100101011" => rgb <= "000000";
					when "00101100100101100" => rgb <= "000000";
					when "00101100100101101" => rgb <= "000000";
					when "00101100100101110" => rgb <= "000000";
					when "00101100100101111" => rgb <= "000000";
					when "00101100100110000" => rgb <= "000000";
					when "00101100100110001" => rgb <= "000000";
					when "00101100100110010" => rgb <= "000000";
					when "00101100100110011" => rgb <= "000000";
					when "00101100100110100" => rgb <= "000000";
					when "00101100100110101" => rgb <= "000000";
					when "00101100100110110" => rgb <= "000000";
					when "00101100100110111" => rgb <= "000000";
					when "00101100100111000" => rgb <= "000000";
					when "00101100100111001" => rgb <= "000000";
					when "00101100100111010" => rgb <= "000000";
					when "00101100100111011" => rgb <= "000000";
					when "00101100100111100" => rgb <= "000000";
					when "00101100100111101" => rgb <= "000000";
					when "00101100100111110" => rgb <= "000000";
					when "00101100100111111" => rgb <= "000000";
					when "00101101000000000" => rgb <= "000000";
					when "00101101000000001" => rgb <= "000000";
					when "00101101000000010" => rgb <= "000000";
					when "00101101000000011" => rgb <= "000000";
					when "00101101000000100" => rgb <= "000000";
					when "00101101000000101" => rgb <= "000000";
					when "00101101000000110" => rgb <= "000000";
					when "00101101000000111" => rgb <= "000000";
					when "00101101000001000" => rgb <= "000000";
					when "00101101000001001" => rgb <= "000000";
					when "00101101000001010" => rgb <= "000000";
					when "00101101000001011" => rgb <= "000000";
					when "00101101000001100" => rgb <= "000000";
					when "00101101000001101" => rgb <= "000000";
					when "00101101000001110" => rgb <= "000000";
					when "00101101000001111" => rgb <= "000000";
					when "00101101000010000" => rgb <= "000000";
					when "00101101000010001" => rgb <= "000000";
					when "00101101000010010" => rgb <= "000000";
					when "00101101000010011" => rgb <= "000000";
					when "00101101000010100" => rgb <= "000000";
					when "00101101000010101" => rgb <= "000000";
					when "00101101000010110" => rgb <= "000000";
					when "00101101000010111" => rgb <= "000000";
					when "00101101000011000" => rgb <= "000000";
					when "00101101000011001" => rgb <= "000000";
					when "00101101000011010" => rgb <= "000000";
					when "00101101000011011" => rgb <= "000000";
					when "00101101000011100" => rgb <= "000000";
					when "00101101000011101" => rgb <= "000000";
					when "00101101000011110" => rgb <= "000000";
					when "00101101000011111" => rgb <= "000000";
					when "00101101000100000" => rgb <= "000000";
					when "00101101000100001" => rgb <= "000000";
					when "00101101000100010" => rgb <= "000000";
					when "00101101000100011" => rgb <= "000000";
					when "00101101000100100" => rgb <= "000000";
					when "00101101000100101" => rgb <= "000000";
					when "00101101000100110" => rgb <= "000000";
					when "00101101000100111" => rgb <= "000000";
					when "00101101000101000" => rgb <= "000000";
					when "00101101000101001" => rgb <= "000000";
					when "00101101000101010" => rgb <= "000000";
					when "00101101000101011" => rgb <= "000000";
					when "00101101000101100" => rgb <= "000000";
					when "00101101000101101" => rgb <= "000000";
					when "00101101000101110" => rgb <= "000000";
					when "00101101000101111" => rgb <= "000000";
					when "00101101000110000" => rgb <= "000000";
					when "00101101000110001" => rgb <= "000000";
					when "00101101000110010" => rgb <= "000000";
					when "00101101000110011" => rgb <= "000000";
					when "00101101000110100" => rgb <= "000000";
					when "00101101000110101" => rgb <= "000000";
					when "00101101000110110" => rgb <= "000000";
					when "00101101000110111" => rgb <= "000000";
					when "00101101000111000" => rgb <= "000000";
					when "00101101000111001" => rgb <= "000000";
					when "00101101000111010" => rgb <= "000000";
					when "00101101000111011" => rgb <= "000000";
					when "00101101000111100" => rgb <= "000000";
					when "00101101000111101" => rgb <= "000000";
					when "00101101000111110" => rgb <= "000000";
					when "00101101000111111" => rgb <= "000000";
					when "00101101001000000" => rgb <= "000000";
					when "00101101001000001" => rgb <= "000000";
					when "00101101001000010" => rgb <= "000000";
					when "00101101001000011" => rgb <= "000000";
					when "00101101001000100" => rgb <= "000000";
					when "00101101001000101" => rgb <= "000000";
					when "00101101001000110" => rgb <= "000000";
					when "00101101001000111" => rgb <= "000000";
					when "00101101001001000" => rgb <= "000000";
					when "00101101001001001" => rgb <= "000000";
					when "00101101001001010" => rgb <= "000000";
					when "00101101001001011" => rgb <= "000000";
					when "00101101001001100" => rgb <= "000000";
					when "00101101001001101" => rgb <= "000000";
					when "00101101001001110" => rgb <= "000000";
					when "00101101001001111" => rgb <= "000000";
					when "00101101001010000" => rgb <= "000000";
					when "00101101001010001" => rgb <= "000000";
					when "00101101001010010" => rgb <= "000000";
					when "00101101001010011" => rgb <= "000000";
					when "00101101001010100" => rgb <= "000000";
					when "00101101001010101" => rgb <= "000000";
					when "00101101001010110" => rgb <= "000000";
					when "00101101001010111" => rgb <= "000000";
					when "00101101001011000" => rgb <= "000000";
					when "00101101001011001" => rgb <= "000000";
					when "00101101001011010" => rgb <= "000000";
					when "00101101001011011" => rgb <= "000000";
					when "00101101001011100" => rgb <= "000000";
					when "00101101001011101" => rgb <= "000000";
					when "00101101001011110" => rgb <= "000000";
					when "00101101001011111" => rgb <= "000000";
					when "00101101001100000" => rgb <= "000000";
					when "00101101001100001" => rgb <= "000000";
					when "00101101001100010" => rgb <= "000000";
					when "00101101001100011" => rgb <= "000000";
					when "00101101001100100" => rgb <= "000000";
					when "00101101001100101" => rgb <= "000000";
					when "00101101001100110" => rgb <= "010100";
					when "00101101001100111" => rgb <= "111000";
					when "00101101001101000" => rgb <= "101000";
					when "00101101001101001" => rgb <= "101000";
					when "00101101001101010" => rgb <= "101000";
					when "00101101001101011" => rgb <= "101000";
					when "00101101001101100" => rgb <= "101000";
					when "00101101001101101" => rgb <= "101000";
					when "00101101001101110" => rgb <= "101000";
					when "00101101001101111" => rgb <= "101000";
					when "00101101001110000" => rgb <= "101000";
					when "00101101001110001" => rgb <= "101000";
					when "00101101001110010" => rgb <= "101000";
					when "00101101001110011" => rgb <= "101000";
					when "00101101001110100" => rgb <= "101000";
					when "00101101001110101" => rgb <= "101000";
					when "00101101001110110" => rgb <= "101000";
					when "00101101001110111" => rgb <= "101000";
					when "00101101001111000" => rgb <= "101000";
					when "00101101001111001" => rgb <= "101000";
					when "00101101001111010" => rgb <= "101000";
					when "00101101001111011" => rgb <= "101000";
					when "00101101001111100" => rgb <= "101000";
					when "00101101001111101" => rgb <= "101000";
					when "00101101001111110" => rgb <= "101000";
					when "00101101001111111" => rgb <= "101000";
					when "00101101010000000" => rgb <= "101000";
					when "00101101010000001" => rgb <= "101000";
					when "00101101010000010" => rgb <= "101000";
					when "00101101010000011" => rgb <= "101000";
					when "00101101010000100" => rgb <= "101000";
					when "00101101010000101" => rgb <= "101000";
					when "00101101010000110" => rgb <= "101000";
					when "00101101010000111" => rgb <= "101000";
					when "00101101010001000" => rgb <= "101001";
					when "00101101010001001" => rgb <= "111001";
					when "00101101010001010" => rgb <= "101001";
					when "00101101010001011" => rgb <= "101001";
					when "00101101010001100" => rgb <= "111001";
					when "00101101010001101" => rgb <= "111001";
					when "00101101010001110" => rgb <= "111001";
					when "00101101010001111" => rgb <= "101001";
					when "00101101010010000" => rgb <= "111001";
					when "00101101010010001" => rgb <= "101001";
					when "00101101010010010" => rgb <= "111001";
					when "00101101010010011" => rgb <= "101001";
					when "00101101010010100" => rgb <= "101000";
					when "00101101010010101" => rgb <= "101000";
					when "00101101010010110" => rgb <= "101000";
					when "00101101010010111" => rgb <= "101000";
					when "00101101010011000" => rgb <= "101000";
					when "00101101010011001" => rgb <= "101000";
					when "00101101010011010" => rgb <= "101000";
					when "00101101010011011" => rgb <= "101000";
					when "00101101010011100" => rgb <= "101000";
					when "00101101010011101" => rgb <= "101000";
					when "00101101010011110" => rgb <= "101000";
					when "00101101010011111" => rgb <= "101000";
					when "00101101010100000" => rgb <= "101000";
					when "00101101010100001" => rgb <= "101000";
					when "00101101010100010" => rgb <= "101000";
					when "00101101010100011" => rgb <= "101000";
					when "00101101010100100" => rgb <= "101000";
					when "00101101010100101" => rgb <= "101000";
					when "00101101010100110" => rgb <= "101000";
					when "00101101010100111" => rgb <= "101000";
					when "00101101010101000" => rgb <= "101000";
					when "00101101010101001" => rgb <= "101000";
					when "00101101010101010" => rgb <= "101000";
					when "00101101010101011" => rgb <= "101000";
					when "00101101010101100" => rgb <= "101000";
					when "00101101010101101" => rgb <= "101000";
					when "00101101010101110" => rgb <= "101000";
					when "00101101010101111" => rgb <= "101000";
					when "00101101010110000" => rgb <= "101000";
					when "00101101010110001" => rgb <= "101000";
					when "00101101010110010" => rgb <= "101000";
					when "00101101010110011" => rgb <= "101000";
					when "00101101010110100" => rgb <= "101000";
					when "00101101010110101" => rgb <= "101000";
					when "00101101010110110" => rgb <= "101000";
					when "00101101010110111" => rgb <= "101000";
					when "00101101010111000" => rgb <= "101000";
					when "00101101010111001" => rgb <= "101000";
					when "00101101010111010" => rgb <= "101000";
					when "00101101010111011" => rgb <= "101000";
					when "00101101010111100" => rgb <= "101000";
					when "00101101010111101" => rgb <= "101000";
					when "00101101010111110" => rgb <= "101000";
					when "00101101010111111" => rgb <= "101000";
					when "00101101011000000" => rgb <= "101000";
					when "00101101011000001" => rgb <= "101000";
					when "00101101011000010" => rgb <= "101000";
					when "00101101011000011" => rgb <= "101000";
					when "00101101011000100" => rgb <= "101000";
					when "00101101011000101" => rgb <= "101000";
					when "00101101011000110" => rgb <= "101000";
					when "00101101011000111" => rgb <= "101000";
					when "00101101011001000" => rgb <= "101000";
					when "00101101011001001" => rgb <= "101000";
					when "00101101011001010" => rgb <= "101000";
					when "00101101011001011" => rgb <= "101000";
					when "00101101011001100" => rgb <= "101000";
					when "00101101011001101" => rgb <= "101000";
					when "00101101011001110" => rgb <= "101000";
					when "00101101011001111" => rgb <= "101000";
					when "00101101011010000" => rgb <= "101000";
					when "00101101011010001" => rgb <= "101000";
					when "00101101011010010" => rgb <= "101000";
					when "00101101011010011" => rgb <= "101000";
					when "00101101011010100" => rgb <= "101000";
					when "00101101011010101" => rgb <= "101000";
					when "00101101011010110" => rgb <= "101000";
					when "00101101011010111" => rgb <= "010100";
					when "00101101011011000" => rgb <= "000000";
					when "00101101011011001" => rgb <= "000000";
					when "00101101011011010" => rgb <= "000000";
					when "00101101011011011" => rgb <= "000000";
					when "00101101011011100" => rgb <= "000000";
					when "00101101011011101" => rgb <= "000000";
					when "00101101011011110" => rgb <= "000000";
					when "00101101011011111" => rgb <= "000000";
					when "00101101011100000" => rgb <= "000000";
					when "00101101011100001" => rgb <= "000000";
					when "00101101011100010" => rgb <= "000000";
					when "00101101011100011" => rgb <= "000000";
					when "00101101011100100" => rgb <= "000000";
					when "00101101011100101" => rgb <= "000000";
					when "00101101011100110" => rgb <= "000000";
					when "00101101011100111" => rgb <= "000000";
					when "00101101011101000" => rgb <= "000000";
					when "00101101011101001" => rgb <= "000000";
					when "00101101011101010" => rgb <= "000000";
					when "00101101011101011" => rgb <= "000000";
					when "00101101011101100" => rgb <= "000000";
					when "00101101011101101" => rgb <= "000000";
					when "00101101011101110" => rgb <= "000000";
					when "00101101011101111" => rgb <= "000000";
					when "00101101011110000" => rgb <= "000000";
					when "00101101011110001" => rgb <= "000000";
					when "00101101011110010" => rgb <= "000000";
					when "00101101011110011" => rgb <= "000000";
					when "00101101011110100" => rgb <= "000000";
					when "00101101011110101" => rgb <= "000000";
					when "00101101011110110" => rgb <= "000000";
					when "00101101011110111" => rgb <= "000000";
					when "00101101011111000" => rgb <= "000000";
					when "00101101011111001" => rgb <= "000000";
					when "00101101011111010" => rgb <= "000000";
					when "00101101011111011" => rgb <= "000000";
					when "00101101011111100" => rgb <= "000000";
					when "00101101011111101" => rgb <= "000000";
					when "00101101011111110" => rgb <= "000000";
					when "00101101011111111" => rgb <= "000000";
					when "00101101100000000" => rgb <= "000000";
					when "00101101100000001" => rgb <= "000000";
					when "00101101100000010" => rgb <= "000000";
					when "00101101100000011" => rgb <= "000000";
					when "00101101100000100" => rgb <= "000000";
					when "00101101100000101" => rgb <= "000000";
					when "00101101100000110" => rgb <= "000000";
					when "00101101100000111" => rgb <= "000000";
					when "00101101100001000" => rgb <= "000000";
					when "00101101100001001" => rgb <= "000000";
					when "00101101100001010" => rgb <= "000000";
					when "00101101100001011" => rgb <= "000000";
					when "00101101100001100" => rgb <= "000000";
					when "00101101100001101" => rgb <= "000000";
					when "00101101100001110" => rgb <= "000000";
					when "00101101100001111" => rgb <= "000000";
					when "00101101100010000" => rgb <= "000000";
					when "00101101100010001" => rgb <= "000000";
					when "00101101100010010" => rgb <= "000000";
					when "00101101100010011" => rgb <= "000000";
					when "00101101100010100" => rgb <= "000000";
					when "00101101100010101" => rgb <= "000000";
					when "00101101100010110" => rgb <= "000000";
					when "00101101100010111" => rgb <= "000000";
					when "00101101100011000" => rgb <= "000000";
					when "00101101100011001" => rgb <= "000000";
					when "00101101100011010" => rgb <= "000000";
					when "00101101100011011" => rgb <= "000000";
					when "00101101100011100" => rgb <= "000000";
					when "00101101100011101" => rgb <= "000000";
					when "00101101100011110" => rgb <= "000000";
					when "00101101100011111" => rgb <= "000000";
					when "00101101100100000" => rgb <= "000000";
					when "00101101100100001" => rgb <= "000000";
					when "00101101100100010" => rgb <= "000000";
					when "00101101100100011" => rgb <= "000000";
					when "00101101100100100" => rgb <= "000000";
					when "00101101100100101" => rgb <= "000000";
					when "00101101100100110" => rgb <= "000000";
					when "00101101100100111" => rgb <= "000000";
					when "00101101100101000" => rgb <= "000000";
					when "00101101100101001" => rgb <= "000000";
					when "00101101100101010" => rgb <= "000000";
					when "00101101100101011" => rgb <= "000000";
					when "00101101100101100" => rgb <= "000000";
					when "00101101100101101" => rgb <= "000000";
					when "00101101100101110" => rgb <= "000000";
					when "00101101100101111" => rgb <= "000000";
					when "00101101100110000" => rgb <= "000000";
					when "00101101100110001" => rgb <= "000000";
					when "00101101100110010" => rgb <= "000000";
					when "00101101100110011" => rgb <= "000000";
					when "00101101100110100" => rgb <= "000000";
					when "00101101100110101" => rgb <= "000000";
					when "00101101100110110" => rgb <= "000000";
					when "00101101100110111" => rgb <= "000000";
					when "00101101100111000" => rgb <= "000000";
					when "00101101100111001" => rgb <= "000000";
					when "00101101100111010" => rgb <= "000000";
					when "00101101100111011" => rgb <= "000000";
					when "00101101100111100" => rgb <= "000000";
					when "00101101100111101" => rgb <= "000000";
					when "00101101100111110" => rgb <= "000000";
					when "00101101100111111" => rgb <= "000000";
					when "00101110000000000" => rgb <= "000000";
					when "00101110000000001" => rgb <= "000000";
					when "00101110000000010" => rgb <= "000000";
					when "00101110000000011" => rgb <= "000000";
					when "00101110000000100" => rgb <= "000000";
					when "00101110000000101" => rgb <= "000000";
					when "00101110000000110" => rgb <= "000000";
					when "00101110000000111" => rgb <= "000000";
					when "00101110000001000" => rgb <= "000000";
					when "00101110000001001" => rgb <= "000000";
					when "00101110000001010" => rgb <= "000000";
					when "00101110000001011" => rgb <= "000000";
					when "00101110000001100" => rgb <= "000000";
					when "00101110000001101" => rgb <= "000000";
					when "00101110000001110" => rgb <= "000000";
					when "00101110000001111" => rgb <= "000000";
					when "00101110000010000" => rgb <= "000000";
					when "00101110000010001" => rgb <= "000000";
					when "00101110000010010" => rgb <= "000000";
					when "00101110000010011" => rgb <= "000000";
					when "00101110000010100" => rgb <= "000000";
					when "00101110000010101" => rgb <= "000000";
					when "00101110000010110" => rgb <= "000000";
					when "00101110000010111" => rgb <= "000000";
					when "00101110000011000" => rgb <= "000000";
					when "00101110000011001" => rgb <= "000000";
					when "00101110000011010" => rgb <= "000000";
					when "00101110000011011" => rgb <= "000000";
					when "00101110000011100" => rgb <= "000000";
					when "00101110000011101" => rgb <= "000000";
					when "00101110000011110" => rgb <= "000000";
					when "00101110000011111" => rgb <= "000000";
					when "00101110000100000" => rgb <= "000000";
					when "00101110000100001" => rgb <= "000000";
					when "00101110000100010" => rgb <= "000000";
					when "00101110000100011" => rgb <= "000000";
					when "00101110000100100" => rgb <= "000000";
					when "00101110000100101" => rgb <= "000000";
					when "00101110000100110" => rgb <= "000000";
					when "00101110000100111" => rgb <= "000000";
					when "00101110000101000" => rgb <= "000000";
					when "00101110000101001" => rgb <= "000000";
					when "00101110000101010" => rgb <= "000000";
					when "00101110000101011" => rgb <= "000000";
					when "00101110000101100" => rgb <= "000000";
					when "00101110000101101" => rgb <= "000000";
					when "00101110000101110" => rgb <= "000000";
					when "00101110000101111" => rgb <= "000000";
					when "00101110000110000" => rgb <= "000000";
					when "00101110000110001" => rgb <= "000000";
					when "00101110000110010" => rgb <= "000000";
					when "00101110000110011" => rgb <= "000000";
					when "00101110000110100" => rgb <= "000000";
					when "00101110000110101" => rgb <= "000000";
					when "00101110000110110" => rgb <= "000000";
					when "00101110000110111" => rgb <= "000000";
					when "00101110000111000" => rgb <= "000000";
					when "00101110000111001" => rgb <= "000000";
					when "00101110000111010" => rgb <= "000000";
					when "00101110000111011" => rgb <= "000000";
					when "00101110000111100" => rgb <= "000000";
					when "00101110000111101" => rgb <= "000000";
					when "00101110000111110" => rgb <= "000000";
					when "00101110000111111" => rgb <= "000000";
					when "00101110001000000" => rgb <= "000000";
					when "00101110001000001" => rgb <= "000000";
					when "00101110001000010" => rgb <= "000000";
					when "00101110001000011" => rgb <= "000000";
					when "00101110001000100" => rgb <= "000000";
					when "00101110001000101" => rgb <= "000000";
					when "00101110001000110" => rgb <= "000000";
					when "00101110001000111" => rgb <= "000000";
					when "00101110001001000" => rgb <= "000000";
					when "00101110001001001" => rgb <= "000000";
					when "00101110001001010" => rgb <= "000000";
					when "00101110001001011" => rgb <= "000000";
					when "00101110001001100" => rgb <= "000000";
					when "00101110001001101" => rgb <= "000000";
					when "00101110001001110" => rgb <= "000000";
					when "00101110001001111" => rgb <= "000000";
					when "00101110001010000" => rgb <= "000000";
					when "00101110001010001" => rgb <= "000000";
					when "00101110001010010" => rgb <= "000000";
					when "00101110001010011" => rgb <= "000000";
					when "00101110001010100" => rgb <= "000000";
					when "00101110001010101" => rgb <= "000000";
					when "00101110001010110" => rgb <= "000000";
					when "00101110001010111" => rgb <= "000000";
					when "00101110001011000" => rgb <= "000000";
					when "00101110001011001" => rgb <= "000000";
					when "00101110001011010" => rgb <= "000000";
					when "00101110001011011" => rgb <= "000000";
					when "00101110001011100" => rgb <= "000000";
					when "00101110001011101" => rgb <= "000000";
					when "00101110001011110" => rgb <= "000000";
					when "00101110001011111" => rgb <= "000000";
					when "00101110001100000" => rgb <= "000000";
					when "00101110001100001" => rgb <= "000000";
					when "00101110001100010" => rgb <= "000000";
					when "00101110001100011" => rgb <= "000000";
					when "00101110001100100" => rgb <= "000000";
					when "00101110001100101" => rgb <= "000000";
					when "00101110001100110" => rgb <= "010100";
					when "00101110001100111" => rgb <= "111000";
					when "00101110001101000" => rgb <= "101000";
					when "00101110001101001" => rgb <= "101000";
					when "00101110001101010" => rgb <= "101000";
					when "00101110001101011" => rgb <= "101000";
					when "00101110001101100" => rgb <= "101000";
					when "00101110001101101" => rgb <= "101000";
					when "00101110001101110" => rgb <= "101000";
					when "00101110001101111" => rgb <= "101000";
					when "00101110001110000" => rgb <= "101000";
					when "00101110001110001" => rgb <= "101000";
					when "00101110001110010" => rgb <= "101000";
					when "00101110001110011" => rgb <= "101000";
					when "00101110001110100" => rgb <= "101000";
					when "00101110001110101" => rgb <= "101000";
					when "00101110001110110" => rgb <= "101000";
					when "00101110001110111" => rgb <= "101000";
					when "00101110001111000" => rgb <= "101000";
					when "00101110001111001" => rgb <= "101000";
					when "00101110001111010" => rgb <= "101000";
					when "00101110001111011" => rgb <= "101000";
					when "00101110001111100" => rgb <= "101000";
					when "00101110001111101" => rgb <= "101000";
					when "00101110001111110" => rgb <= "101000";
					when "00101110001111111" => rgb <= "101000";
					when "00101110010000000" => rgb <= "101000";
					when "00101110010000001" => rgb <= "101000";
					when "00101110010000010" => rgb <= "101000";
					when "00101110010000011" => rgb <= "101000";
					when "00101110010000100" => rgb <= "101000";
					when "00101110010000101" => rgb <= "101000";
					when "00101110010000110" => rgb <= "101000";
					when "00101110010000111" => rgb <= "101000";
					when "00101110010001000" => rgb <= "101001";
					when "00101110010001001" => rgb <= "111001";
					when "00101110010001010" => rgb <= "101001";
					when "00101110010001011" => rgb <= "101001";
					when "00101110010001100" => rgb <= "111001";
					when "00101110010001101" => rgb <= "111001";
					when "00101110010001110" => rgb <= "111001";
					when "00101110010001111" => rgb <= "101001";
					when "00101110010010000" => rgb <= "111001";
					when "00101110010010001" => rgb <= "101001";
					when "00101110010010010" => rgb <= "111001";
					when "00101110010010011" => rgb <= "101001";
					when "00101110010010100" => rgb <= "101000";
					when "00101110010010101" => rgb <= "101000";
					when "00101110010010110" => rgb <= "101000";
					when "00101110010010111" => rgb <= "101000";
					when "00101110010011000" => rgb <= "101000";
					when "00101110010011001" => rgb <= "101000";
					when "00101110010011010" => rgb <= "101000";
					when "00101110010011011" => rgb <= "101000";
					when "00101110010011100" => rgb <= "101000";
					when "00101110010011101" => rgb <= "101000";
					when "00101110010011110" => rgb <= "101000";
					when "00101110010011111" => rgb <= "101000";
					when "00101110010100000" => rgb <= "101000";
					when "00101110010100001" => rgb <= "101000";
					when "00101110010100010" => rgb <= "101000";
					when "00101110010100011" => rgb <= "101000";
					when "00101110010100100" => rgb <= "101000";
					when "00101110010100101" => rgb <= "101000";
					when "00101110010100110" => rgb <= "101000";
					when "00101110010100111" => rgb <= "101000";
					when "00101110010101000" => rgb <= "101000";
					when "00101110010101001" => rgb <= "101000";
					when "00101110010101010" => rgb <= "101000";
					when "00101110010101011" => rgb <= "101000";
					when "00101110010101100" => rgb <= "101000";
					when "00101110010101101" => rgb <= "101000";
					when "00101110010101110" => rgb <= "101000";
					when "00101110010101111" => rgb <= "101000";
					when "00101110010110000" => rgb <= "101000";
					when "00101110010110001" => rgb <= "101000";
					when "00101110010110010" => rgb <= "101000";
					when "00101110010110011" => rgb <= "101000";
					when "00101110010110100" => rgb <= "101000";
					when "00101110010110101" => rgb <= "101000";
					when "00101110010110110" => rgb <= "101000";
					when "00101110010110111" => rgb <= "101000";
					when "00101110010111000" => rgb <= "101000";
					when "00101110010111001" => rgb <= "101000";
					when "00101110010111010" => rgb <= "101000";
					when "00101110010111011" => rgb <= "101000";
					when "00101110010111100" => rgb <= "101000";
					when "00101110010111101" => rgb <= "101000";
					when "00101110010111110" => rgb <= "101000";
					when "00101110010111111" => rgb <= "101000";
					when "00101110011000000" => rgb <= "101000";
					when "00101110011000001" => rgb <= "101000";
					when "00101110011000010" => rgb <= "101000";
					when "00101110011000011" => rgb <= "101000";
					when "00101110011000100" => rgb <= "101000";
					when "00101110011000101" => rgb <= "101000";
					when "00101110011000110" => rgb <= "101000";
					when "00101110011000111" => rgb <= "101000";
					when "00101110011001000" => rgb <= "101000";
					when "00101110011001001" => rgb <= "101000";
					when "00101110011001010" => rgb <= "101000";
					when "00101110011001011" => rgb <= "101000";
					when "00101110011001100" => rgb <= "101000";
					when "00101110011001101" => rgb <= "101000";
					when "00101110011001110" => rgb <= "101000";
					when "00101110011001111" => rgb <= "101000";
					when "00101110011010000" => rgb <= "101000";
					when "00101110011010001" => rgb <= "101000";
					when "00101110011010010" => rgb <= "101000";
					when "00101110011010011" => rgb <= "101000";
					when "00101110011010100" => rgb <= "101000";
					when "00101110011010101" => rgb <= "101000";
					when "00101110011010110" => rgb <= "101000";
					when "00101110011010111" => rgb <= "010100";
					when "00101110011011000" => rgb <= "000000";
					when "00101110011011001" => rgb <= "000000";
					when "00101110011011010" => rgb <= "000000";
					when "00101110011011011" => rgb <= "000000";
					when "00101110011011100" => rgb <= "000000";
					when "00101110011011101" => rgb <= "000000";
					when "00101110011011110" => rgb <= "000000";
					when "00101110011011111" => rgb <= "000000";
					when "00101110011100000" => rgb <= "000000";
					when "00101110011100001" => rgb <= "000000";
					when "00101110011100010" => rgb <= "000000";
					when "00101110011100011" => rgb <= "000000";
					when "00101110011100100" => rgb <= "000000";
					when "00101110011100101" => rgb <= "000000";
					when "00101110011100110" => rgb <= "000000";
					when "00101110011100111" => rgb <= "000000";
					when "00101110011101000" => rgb <= "000000";
					when "00101110011101001" => rgb <= "000000";
					when "00101110011101010" => rgb <= "000000";
					when "00101110011101011" => rgb <= "000000";
					when "00101110011101100" => rgb <= "000000";
					when "00101110011101101" => rgb <= "000000";
					when "00101110011101110" => rgb <= "000000";
					when "00101110011101111" => rgb <= "000000";
					when "00101110011110000" => rgb <= "000000";
					when "00101110011110001" => rgb <= "000000";
					when "00101110011110010" => rgb <= "000000";
					when "00101110011110011" => rgb <= "000000";
					when "00101110011110100" => rgb <= "000000";
					when "00101110011110101" => rgb <= "000000";
					when "00101110011110110" => rgb <= "000000";
					when "00101110011110111" => rgb <= "000000";
					when "00101110011111000" => rgb <= "000000";
					when "00101110011111001" => rgb <= "000000";
					when "00101110011111010" => rgb <= "000000";
					when "00101110011111011" => rgb <= "000000";
					when "00101110011111100" => rgb <= "000000";
					when "00101110011111101" => rgb <= "000000";
					when "00101110011111110" => rgb <= "000000";
					when "00101110011111111" => rgb <= "000000";
					when "00101110100000000" => rgb <= "000000";
					when "00101110100000001" => rgb <= "000000";
					when "00101110100000010" => rgb <= "000000";
					when "00101110100000011" => rgb <= "000000";
					when "00101110100000100" => rgb <= "000000";
					when "00101110100000101" => rgb <= "000000";
					when "00101110100000110" => rgb <= "000000";
					when "00101110100000111" => rgb <= "000000";
					when "00101110100001000" => rgb <= "000000";
					when "00101110100001001" => rgb <= "000000";
					when "00101110100001010" => rgb <= "000000";
					when "00101110100001011" => rgb <= "000000";
					when "00101110100001100" => rgb <= "000000";
					when "00101110100001101" => rgb <= "000000";
					when "00101110100001110" => rgb <= "000000";
					when "00101110100001111" => rgb <= "000000";
					when "00101110100010000" => rgb <= "000000";
					when "00101110100010001" => rgb <= "000000";
					when "00101110100010010" => rgb <= "000000";
					when "00101110100010011" => rgb <= "000000";
					when "00101110100010100" => rgb <= "000000";
					when "00101110100010101" => rgb <= "000000";
					when "00101110100010110" => rgb <= "000000";
					when "00101110100010111" => rgb <= "000000";
					when "00101110100011000" => rgb <= "000000";
					when "00101110100011001" => rgb <= "000000";
					when "00101110100011010" => rgb <= "000000";
					when "00101110100011011" => rgb <= "000000";
					when "00101110100011100" => rgb <= "000000";
					when "00101110100011101" => rgb <= "000000";
					when "00101110100011110" => rgb <= "000000";
					when "00101110100011111" => rgb <= "000000";
					when "00101110100100000" => rgb <= "000000";
					when "00101110100100001" => rgb <= "000000";
					when "00101110100100010" => rgb <= "000000";
					when "00101110100100011" => rgb <= "000000";
					when "00101110100100100" => rgb <= "000000";
					when "00101110100100101" => rgb <= "000000";
					when "00101110100100110" => rgb <= "000000";
					when "00101110100100111" => rgb <= "000000";
					when "00101110100101000" => rgb <= "000000";
					when "00101110100101001" => rgb <= "000000";
					when "00101110100101010" => rgb <= "000000";
					when "00101110100101011" => rgb <= "000000";
					when "00101110100101100" => rgb <= "000000";
					when "00101110100101101" => rgb <= "000000";
					when "00101110100101110" => rgb <= "000000";
					when "00101110100101111" => rgb <= "000000";
					when "00101110100110000" => rgb <= "000000";
					when "00101110100110001" => rgb <= "000000";
					when "00101110100110010" => rgb <= "000000";
					when "00101110100110011" => rgb <= "000000";
					when "00101110100110100" => rgb <= "000000";
					when "00101110100110101" => rgb <= "000000";
					when "00101110100110110" => rgb <= "000000";
					when "00101110100110111" => rgb <= "000000";
					when "00101110100111000" => rgb <= "000000";
					when "00101110100111001" => rgb <= "000000";
					when "00101110100111010" => rgb <= "000000";
					when "00101110100111011" => rgb <= "000000";
					when "00101110100111100" => rgb <= "000000";
					when "00101110100111101" => rgb <= "000000";
					when "00101110100111110" => rgb <= "000000";
					when "00101110100111111" => rgb <= "000000";
					when "00101111000000000" => rgb <= "000000";
					when "00101111000000001" => rgb <= "000000";
					when "00101111000000010" => rgb <= "000000";
					when "00101111000000011" => rgb <= "000000";
					when "00101111000000100" => rgb <= "000000";
					when "00101111000000101" => rgb <= "000000";
					when "00101111000000110" => rgb <= "000000";
					when "00101111000000111" => rgb <= "000000";
					when "00101111000001000" => rgb <= "000000";
					when "00101111000001001" => rgb <= "000000";
					when "00101111000001010" => rgb <= "000000";
					when "00101111000001011" => rgb <= "000000";
					when "00101111000001100" => rgb <= "000000";
					when "00101111000001101" => rgb <= "000000";
					when "00101111000001110" => rgb <= "000000";
					when "00101111000001111" => rgb <= "000000";
					when "00101111000010000" => rgb <= "000000";
					when "00101111000010001" => rgb <= "000000";
					when "00101111000010010" => rgb <= "000000";
					when "00101111000010011" => rgb <= "000000";
					when "00101111000010100" => rgb <= "000000";
					when "00101111000010101" => rgb <= "000000";
					when "00101111000010110" => rgb <= "000000";
					when "00101111000010111" => rgb <= "000000";
					when "00101111000011000" => rgb <= "000000";
					when "00101111000011001" => rgb <= "000000";
					when "00101111000011010" => rgb <= "000000";
					when "00101111000011011" => rgb <= "000000";
					when "00101111000011100" => rgb <= "000000";
					when "00101111000011101" => rgb <= "000000";
					when "00101111000011110" => rgb <= "000000";
					when "00101111000011111" => rgb <= "000000";
					when "00101111000100000" => rgb <= "000000";
					when "00101111000100001" => rgb <= "000000";
					when "00101111000100010" => rgb <= "000000";
					when "00101111000100011" => rgb <= "000000";
					when "00101111000100100" => rgb <= "000000";
					when "00101111000100101" => rgb <= "000000";
					when "00101111000100110" => rgb <= "000000";
					when "00101111000100111" => rgb <= "000000";
					when "00101111000101000" => rgb <= "000000";
					when "00101111000101001" => rgb <= "000000";
					when "00101111000101010" => rgb <= "000000";
					when "00101111000101011" => rgb <= "000000";
					when "00101111000101100" => rgb <= "000000";
					when "00101111000101101" => rgb <= "000000";
					when "00101111000101110" => rgb <= "000000";
					when "00101111000101111" => rgb <= "000000";
					when "00101111000110000" => rgb <= "000000";
					when "00101111000110001" => rgb <= "000000";
					when "00101111000110010" => rgb <= "000000";
					when "00101111000110011" => rgb <= "000000";
					when "00101111000110100" => rgb <= "000000";
					when "00101111000110101" => rgb <= "000000";
					when "00101111000110110" => rgb <= "000000";
					when "00101111000110111" => rgb <= "000000";
					when "00101111000111000" => rgb <= "000000";
					when "00101111000111001" => rgb <= "000000";
					when "00101111000111010" => rgb <= "000000";
					when "00101111000111011" => rgb <= "000000";
					when "00101111000111100" => rgb <= "000000";
					when "00101111000111101" => rgb <= "000000";
					when "00101111000111110" => rgb <= "000000";
					when "00101111000111111" => rgb <= "000000";
					when "00101111001000000" => rgb <= "000000";
					when "00101111001000001" => rgb <= "000000";
					when "00101111001000010" => rgb <= "000000";
					when "00101111001000011" => rgb <= "000000";
					when "00101111001000100" => rgb <= "000000";
					when "00101111001000101" => rgb <= "000000";
					when "00101111001000110" => rgb <= "000000";
					when "00101111001000111" => rgb <= "000000";
					when "00101111001001000" => rgb <= "000000";
					when "00101111001001001" => rgb <= "000000";
					when "00101111001001010" => rgb <= "000000";
					when "00101111001001011" => rgb <= "000000";
					when "00101111001001100" => rgb <= "000000";
					when "00101111001001101" => rgb <= "000000";
					when "00101111001001110" => rgb <= "000000";
					when "00101111001001111" => rgb <= "000000";
					when "00101111001010000" => rgb <= "000000";
					when "00101111001010001" => rgb <= "000000";
					when "00101111001010010" => rgb <= "000000";
					when "00101111001010011" => rgb <= "000000";
					when "00101111001010100" => rgb <= "000000";
					when "00101111001010101" => rgb <= "000000";
					when "00101111001010110" => rgb <= "000000";
					when "00101111001010111" => rgb <= "000000";
					when "00101111001011000" => rgb <= "000000";
					when "00101111001011001" => rgb <= "000000";
					when "00101111001011010" => rgb <= "000000";
					when "00101111001011011" => rgb <= "000000";
					when "00101111001011100" => rgb <= "000000";
					when "00101111001011101" => rgb <= "000000";
					when "00101111001011110" => rgb <= "000000";
					when "00101111001011111" => rgb <= "000000";
					when "00101111001100000" => rgb <= "000000";
					when "00101111001100001" => rgb <= "000000";
					when "00101111001100010" => rgb <= "000000";
					when "00101111001100011" => rgb <= "000000";
					when "00101111001100100" => rgb <= "000000";
					when "00101111001100101" => rgb <= "000000";
					when "00101111001100110" => rgb <= "010100";
					when "00101111001100111" => rgb <= "111000";
					when "00101111001101000" => rgb <= "101000";
					when "00101111001101001" => rgb <= "101000";
					when "00101111001101010" => rgb <= "101000";
					when "00101111001101011" => rgb <= "101000";
					when "00101111001101100" => rgb <= "101000";
					when "00101111001101101" => rgb <= "101000";
					when "00101111001101110" => rgb <= "101000";
					when "00101111001101111" => rgb <= "101000";
					when "00101111001110000" => rgb <= "101000";
					when "00101111001110001" => rgb <= "101000";
					when "00101111001110010" => rgb <= "101000";
					when "00101111001110011" => rgb <= "101000";
					when "00101111001110100" => rgb <= "101000";
					when "00101111001110101" => rgb <= "101000";
					when "00101111001110110" => rgb <= "101000";
					when "00101111001110111" => rgb <= "101000";
					when "00101111001111000" => rgb <= "101000";
					when "00101111001111001" => rgb <= "101000";
					when "00101111001111010" => rgb <= "101000";
					when "00101111001111011" => rgb <= "101000";
					when "00101111001111100" => rgb <= "101000";
					when "00101111001111101" => rgb <= "101000";
					when "00101111001111110" => rgb <= "101000";
					when "00101111001111111" => rgb <= "101000";
					when "00101111010000000" => rgb <= "101000";
					when "00101111010000001" => rgb <= "101000";
					when "00101111010000010" => rgb <= "101000";
					when "00101111010000011" => rgb <= "101000";
					when "00101111010000100" => rgb <= "101000";
					when "00101111010000101" => rgb <= "101000";
					when "00101111010000110" => rgb <= "101000";
					when "00101111010000111" => rgb <= "101000";
					when "00101111010001000" => rgb <= "101001";
					when "00101111010001001" => rgb <= "111001";
					when "00101111010001010" => rgb <= "101001";
					when "00101111010001011" => rgb <= "101001";
					when "00101111010001100" => rgb <= "111001";
					when "00101111010001101" => rgb <= "111001";
					when "00101111010001110" => rgb <= "111001";
					when "00101111010001111" => rgb <= "101001";
					when "00101111010010000" => rgb <= "111001";
					when "00101111010010001" => rgb <= "101001";
					when "00101111010010010" => rgb <= "111001";
					when "00101111010010011" => rgb <= "101001";
					when "00101111010010100" => rgb <= "101000";
					when "00101111010010101" => rgb <= "101000";
					when "00101111010010110" => rgb <= "101000";
					when "00101111010010111" => rgb <= "101000";
					when "00101111010011000" => rgb <= "101000";
					when "00101111010011001" => rgb <= "101000";
					when "00101111010011010" => rgb <= "101000";
					when "00101111010011011" => rgb <= "101000";
					when "00101111010011100" => rgb <= "101000";
					when "00101111010011101" => rgb <= "101000";
					when "00101111010011110" => rgb <= "101000";
					when "00101111010011111" => rgb <= "101000";
					when "00101111010100000" => rgb <= "101000";
					when "00101111010100001" => rgb <= "101000";
					when "00101111010100010" => rgb <= "101000";
					when "00101111010100011" => rgb <= "101000";
					when "00101111010100100" => rgb <= "101000";
					when "00101111010100101" => rgb <= "101000";
					when "00101111010100110" => rgb <= "101000";
					when "00101111010100111" => rgb <= "101000";
					when "00101111010101000" => rgb <= "101000";
					when "00101111010101001" => rgb <= "101000";
					when "00101111010101010" => rgb <= "101000";
					when "00101111010101011" => rgb <= "101000";
					when "00101111010101100" => rgb <= "101000";
					when "00101111010101101" => rgb <= "101000";
					when "00101111010101110" => rgb <= "101000";
					when "00101111010101111" => rgb <= "101000";
					when "00101111010110000" => rgb <= "101000";
					when "00101111010110001" => rgb <= "101000";
					when "00101111010110010" => rgb <= "101000";
					when "00101111010110011" => rgb <= "101000";
					when "00101111010110100" => rgb <= "101000";
					when "00101111010110101" => rgb <= "101000";
					when "00101111010110110" => rgb <= "101000";
					when "00101111010110111" => rgb <= "101000";
					when "00101111010111000" => rgb <= "101000";
					when "00101111010111001" => rgb <= "101000";
					when "00101111010111010" => rgb <= "101000";
					when "00101111010111011" => rgb <= "101000";
					when "00101111010111100" => rgb <= "101000";
					when "00101111010111101" => rgb <= "101000";
					when "00101111010111110" => rgb <= "101000";
					when "00101111010111111" => rgb <= "101000";
					when "00101111011000000" => rgb <= "101000";
					when "00101111011000001" => rgb <= "101000";
					when "00101111011000010" => rgb <= "101000";
					when "00101111011000011" => rgb <= "101000";
					when "00101111011000100" => rgb <= "101000";
					when "00101111011000101" => rgb <= "101000";
					when "00101111011000110" => rgb <= "101000";
					when "00101111011000111" => rgb <= "101000";
					when "00101111011001000" => rgb <= "101000";
					when "00101111011001001" => rgb <= "101000";
					when "00101111011001010" => rgb <= "101000";
					when "00101111011001011" => rgb <= "101000";
					when "00101111011001100" => rgb <= "101000";
					when "00101111011001101" => rgb <= "101000";
					when "00101111011001110" => rgb <= "101000";
					when "00101111011001111" => rgb <= "101000";
					when "00101111011010000" => rgb <= "101000";
					when "00101111011010001" => rgb <= "101000";
					when "00101111011010010" => rgb <= "101000";
					when "00101111011010011" => rgb <= "101000";
					when "00101111011010100" => rgb <= "101000";
					when "00101111011010101" => rgb <= "101000";
					when "00101111011010110" => rgb <= "101000";
					when "00101111011010111" => rgb <= "010100";
					when "00101111011011000" => rgb <= "000000";
					when "00101111011011001" => rgb <= "000000";
					when "00101111011011010" => rgb <= "000000";
					when "00101111011011011" => rgb <= "000000";
					when "00101111011011100" => rgb <= "000000";
					when "00101111011011101" => rgb <= "000000";
					when "00101111011011110" => rgb <= "000000";
					when "00101111011011111" => rgb <= "000000";
					when "00101111011100000" => rgb <= "000000";
					when "00101111011100001" => rgb <= "000000";
					when "00101111011100010" => rgb <= "000000";
					when "00101111011100011" => rgb <= "000000";
					when "00101111011100100" => rgb <= "000000";
					when "00101111011100101" => rgb <= "000000";
					when "00101111011100110" => rgb <= "000000";
					when "00101111011100111" => rgb <= "000000";
					when "00101111011101000" => rgb <= "000000";
					when "00101111011101001" => rgb <= "000000";
					when "00101111011101010" => rgb <= "000000";
					when "00101111011101011" => rgb <= "000000";
					when "00101111011101100" => rgb <= "000000";
					when "00101111011101101" => rgb <= "000000";
					when "00101111011101110" => rgb <= "000000";
					when "00101111011101111" => rgb <= "000000";
					when "00101111011110000" => rgb <= "000000";
					when "00101111011110001" => rgb <= "000000";
					when "00101111011110010" => rgb <= "000000";
					when "00101111011110011" => rgb <= "000000";
					when "00101111011110100" => rgb <= "000000";
					when "00101111011110101" => rgb <= "000000";
					when "00101111011110110" => rgb <= "000000";
					when "00101111011110111" => rgb <= "000000";
					when "00101111011111000" => rgb <= "000000";
					when "00101111011111001" => rgb <= "000000";
					when "00101111011111010" => rgb <= "000000";
					when "00101111011111011" => rgb <= "000000";
					when "00101111011111100" => rgb <= "000000";
					when "00101111011111101" => rgb <= "000000";
					when "00101111011111110" => rgb <= "000000";
					when "00101111011111111" => rgb <= "000000";
					when "00101111100000000" => rgb <= "000000";
					when "00101111100000001" => rgb <= "000000";
					when "00101111100000010" => rgb <= "000000";
					when "00101111100000011" => rgb <= "000000";
					when "00101111100000100" => rgb <= "000000";
					when "00101111100000101" => rgb <= "000000";
					when "00101111100000110" => rgb <= "000000";
					when "00101111100000111" => rgb <= "000000";
					when "00101111100001000" => rgb <= "000000";
					when "00101111100001001" => rgb <= "000000";
					when "00101111100001010" => rgb <= "000000";
					when "00101111100001011" => rgb <= "000000";
					when "00101111100001100" => rgb <= "000000";
					when "00101111100001101" => rgb <= "000000";
					when "00101111100001110" => rgb <= "000000";
					when "00101111100001111" => rgb <= "000000";
					when "00101111100010000" => rgb <= "000000";
					when "00101111100010001" => rgb <= "000000";
					when "00101111100010010" => rgb <= "000000";
					when "00101111100010011" => rgb <= "000000";
					when "00101111100010100" => rgb <= "000000";
					when "00101111100010101" => rgb <= "000000";
					when "00101111100010110" => rgb <= "000000";
					when "00101111100010111" => rgb <= "000000";
					when "00101111100011000" => rgb <= "000000";
					when "00101111100011001" => rgb <= "000000";
					when "00101111100011010" => rgb <= "000000";
					when "00101111100011011" => rgb <= "000000";
					when "00101111100011100" => rgb <= "000000";
					when "00101111100011101" => rgb <= "000000";
					when "00101111100011110" => rgb <= "000000";
					when "00101111100011111" => rgb <= "000000";
					when "00101111100100000" => rgb <= "000000";
					when "00101111100100001" => rgb <= "000000";
					when "00101111100100010" => rgb <= "000000";
					when "00101111100100011" => rgb <= "000000";
					when "00101111100100100" => rgb <= "000000";
					when "00101111100100101" => rgb <= "000000";
					when "00101111100100110" => rgb <= "000000";
					when "00101111100100111" => rgb <= "000000";
					when "00101111100101000" => rgb <= "000000";
					when "00101111100101001" => rgb <= "000000";
					when "00101111100101010" => rgb <= "000000";
					when "00101111100101011" => rgb <= "000000";
					when "00101111100101100" => rgb <= "000000";
					when "00101111100101101" => rgb <= "000000";
					when "00101111100101110" => rgb <= "000000";
					when "00101111100101111" => rgb <= "000000";
					when "00101111100110000" => rgb <= "000000";
					when "00101111100110001" => rgb <= "000000";
					when "00101111100110010" => rgb <= "000000";
					when "00101111100110011" => rgb <= "000000";
					when "00101111100110100" => rgb <= "000000";
					when "00101111100110101" => rgb <= "000000";
					when "00101111100110110" => rgb <= "000000";
					when "00101111100110111" => rgb <= "000000";
					when "00101111100111000" => rgb <= "000000";
					when "00101111100111001" => rgb <= "000000";
					when "00101111100111010" => rgb <= "000000";
					when "00101111100111011" => rgb <= "000000";
					when "00101111100111100" => rgb <= "000000";
					when "00101111100111101" => rgb <= "000000";
					when "00101111100111110" => rgb <= "000000";
					when "00101111100111111" => rgb <= "000000";
					when "00110000000000000" => rgb <= "000000";
					when "00110000000000001" => rgb <= "000000";
					when "00110000000000010" => rgb <= "000000";
					when "00110000000000011" => rgb <= "000000";
					when "00110000000000100" => rgb <= "000000";
					when "00110000000000101" => rgb <= "000000";
					when "00110000000000110" => rgb <= "000000";
					when "00110000000000111" => rgb <= "000000";
					when "00110000000001000" => rgb <= "000000";
					when "00110000000001001" => rgb <= "000000";
					when "00110000000001010" => rgb <= "000000";
					when "00110000000001011" => rgb <= "000000";
					when "00110000000001100" => rgb <= "000000";
					when "00110000000001101" => rgb <= "000000";
					when "00110000000001110" => rgb <= "000000";
					when "00110000000001111" => rgb <= "000000";
					when "00110000000010000" => rgb <= "000000";
					when "00110000000010001" => rgb <= "000000";
					when "00110000000010010" => rgb <= "000000";
					when "00110000000010011" => rgb <= "000000";
					when "00110000000010100" => rgb <= "000000";
					when "00110000000010101" => rgb <= "000000";
					when "00110000000010110" => rgb <= "000000";
					when "00110000000010111" => rgb <= "000000";
					when "00110000000011000" => rgb <= "000000";
					when "00110000000011001" => rgb <= "000000";
					when "00110000000011010" => rgb <= "000000";
					when "00110000000011011" => rgb <= "000000";
					when "00110000000011100" => rgb <= "000000";
					when "00110000000011101" => rgb <= "000000";
					when "00110000000011110" => rgb <= "000000";
					when "00110000000011111" => rgb <= "000000";
					when "00110000000100000" => rgb <= "000000";
					when "00110000000100001" => rgb <= "000000";
					when "00110000000100010" => rgb <= "000000";
					when "00110000000100011" => rgb <= "000000";
					when "00110000000100100" => rgb <= "000000";
					when "00110000000100101" => rgb <= "000000";
					when "00110000000100110" => rgb <= "000000";
					when "00110000000100111" => rgb <= "000000";
					when "00110000000101000" => rgb <= "000000";
					when "00110000000101001" => rgb <= "000000";
					when "00110000000101010" => rgb <= "000000";
					when "00110000000101011" => rgb <= "000000";
					when "00110000000101100" => rgb <= "000000";
					when "00110000000101101" => rgb <= "000000";
					when "00110000000101110" => rgb <= "000000";
					when "00110000000101111" => rgb <= "000000";
					when "00110000000110000" => rgb <= "000000";
					when "00110000000110001" => rgb <= "000000";
					when "00110000000110010" => rgb <= "000000";
					when "00110000000110011" => rgb <= "000000";
					when "00110000000110100" => rgb <= "000000";
					when "00110000000110101" => rgb <= "000000";
					when "00110000000110110" => rgb <= "000000";
					when "00110000000110111" => rgb <= "000000";
					when "00110000000111000" => rgb <= "000000";
					when "00110000000111001" => rgb <= "000000";
					when "00110000000111010" => rgb <= "000000";
					when "00110000000111011" => rgb <= "000000";
					when "00110000000111100" => rgb <= "000000";
					when "00110000000111101" => rgb <= "000000";
					when "00110000000111110" => rgb <= "000000";
					when "00110000000111111" => rgb <= "000000";
					when "00110000001000000" => rgb <= "000000";
					when "00110000001000001" => rgb <= "000000";
					when "00110000001000010" => rgb <= "000000";
					when "00110000001000011" => rgb <= "000000";
					when "00110000001000100" => rgb <= "000000";
					when "00110000001000101" => rgb <= "000000";
					when "00110000001000110" => rgb <= "000000";
					when "00110000001000111" => rgb <= "000000";
					when "00110000001001000" => rgb <= "000000";
					when "00110000001001001" => rgb <= "000000";
					when "00110000001001010" => rgb <= "000000";
					when "00110000001001011" => rgb <= "000000";
					when "00110000001001100" => rgb <= "000000";
					when "00110000001001101" => rgb <= "000000";
					when "00110000001001110" => rgb <= "000000";
					when "00110000001001111" => rgb <= "000000";
					when "00110000001010000" => rgb <= "000000";
					when "00110000001010001" => rgb <= "000000";
					when "00110000001010010" => rgb <= "000000";
					when "00110000001010011" => rgb <= "000000";
					when "00110000001010100" => rgb <= "000000";
					when "00110000001010101" => rgb <= "000000";
					when "00110000001010110" => rgb <= "000000";
					when "00110000001010111" => rgb <= "000000";
					when "00110000001011000" => rgb <= "000000";
					when "00110000001011001" => rgb <= "000000";
					when "00110000001011010" => rgb <= "000000";
					when "00110000001011011" => rgb <= "000000";
					when "00110000001011100" => rgb <= "000000";
					when "00110000001011101" => rgb <= "000000";
					when "00110000001011110" => rgb <= "000000";
					when "00110000001011111" => rgb <= "000000";
					when "00110000001100000" => rgb <= "000000";
					when "00110000001100001" => rgb <= "000000";
					when "00110000001100010" => rgb <= "000000";
					when "00110000001100011" => rgb <= "000000";
					when "00110000001100100" => rgb <= "000000";
					when "00110000001100101" => rgb <= "000000";
					when "00110000001100110" => rgb <= "010100";
					when "00110000001100111" => rgb <= "111000";
					when "00110000001101000" => rgb <= "101000";
					when "00110000001101001" => rgb <= "101000";
					when "00110000001101010" => rgb <= "101000";
					when "00110000001101011" => rgb <= "101000";
					when "00110000001101100" => rgb <= "101000";
					when "00110000001101101" => rgb <= "101000";
					when "00110000001101110" => rgb <= "101000";
					when "00110000001101111" => rgb <= "101000";
					when "00110000001110000" => rgb <= "101000";
					when "00110000001110001" => rgb <= "101000";
					when "00110000001110010" => rgb <= "101000";
					when "00110000001110011" => rgb <= "101000";
					when "00110000001110100" => rgb <= "101000";
					when "00110000001110101" => rgb <= "101000";
					when "00110000001110110" => rgb <= "101000";
					when "00110000001110111" => rgb <= "101000";
					when "00110000001111000" => rgb <= "101000";
					when "00110000001111001" => rgb <= "101000";
					when "00110000001111010" => rgb <= "101000";
					when "00110000001111011" => rgb <= "101000";
					when "00110000001111100" => rgb <= "101000";
					when "00110000001111101" => rgb <= "111001";
					when "00110000001111110" => rgb <= "101000";
					when "00110000001111111" => rgb <= "101000";
					when "00110000010000000" => rgb <= "101000";
					when "00110000010000001" => rgb <= "101000";
					when "00110000010000010" => rgb <= "101000";
					when "00110000010000011" => rgb <= "101000";
					when "00110000010000100" => rgb <= "101000";
					when "00110000010000101" => rgb <= "101000";
					when "00110000010000110" => rgb <= "101000";
					when "00110000010000111" => rgb <= "101000";
					when "00110000010001000" => rgb <= "101001";
					when "00110000010001001" => rgb <= "111001";
					when "00110000010001010" => rgb <= "111001";
					when "00110000010001011" => rgb <= "111001";
					when "00110000010001100" => rgb <= "111001";
					when "00110000010001101" => rgb <= "111001";
					when "00110000010001110" => rgb <= "111001";
					when "00110000010001111" => rgb <= "111001";
					when "00110000010010000" => rgb <= "101001";
					when "00110000010010001" => rgb <= "101001";
					when "00110000010010010" => rgb <= "101001";
					when "00110000010010011" => rgb <= "101001";
					when "00110000010010100" => rgb <= "101000";
					when "00110000010010101" => rgb <= "101000";
					when "00110000010010110" => rgb <= "101000";
					when "00110000010010111" => rgb <= "101000";
					when "00110000010011000" => rgb <= "101000";
					when "00110000010011001" => rgb <= "101000";
					when "00110000010011010" => rgb <= "101000";
					when "00110000010011011" => rgb <= "101000";
					when "00110000010011100" => rgb <= "101000";
					when "00110000010011101" => rgb <= "101000";
					when "00110000010011110" => rgb <= "101000";
					when "00110000010011111" => rgb <= "101000";
					when "00110000010100000" => rgb <= "101000";
					when "00110000010100001" => rgb <= "101000";
					when "00110000010100010" => rgb <= "101000";
					when "00110000010100011" => rgb <= "101000";
					when "00110000010100100" => rgb <= "101000";
					when "00110000010100101" => rgb <= "101000";
					when "00110000010100110" => rgb <= "101000";
					when "00110000010100111" => rgb <= "101000";
					when "00110000010101000" => rgb <= "101000";
					when "00110000010101001" => rgb <= "101000";
					when "00110000010101010" => rgb <= "101000";
					when "00110000010101011" => rgb <= "101000";
					when "00110000010101100" => rgb <= "101000";
					when "00110000010101101" => rgb <= "101000";
					when "00110000010101110" => rgb <= "101000";
					when "00110000010101111" => rgb <= "101000";
					when "00110000010110000" => rgb <= "101000";
					when "00110000010110001" => rgb <= "101000";
					when "00110000010110010" => rgb <= "101000";
					when "00110000010110011" => rgb <= "101000";
					when "00110000010110100" => rgb <= "101000";
					when "00110000010110101" => rgb <= "101000";
					when "00110000010110110" => rgb <= "101000";
					when "00110000010110111" => rgb <= "101000";
					when "00110000010111000" => rgb <= "101000";
					when "00110000010111001" => rgb <= "101000";
					when "00110000010111010" => rgb <= "101000";
					when "00110000010111011" => rgb <= "101000";
					when "00110000010111100" => rgb <= "101000";
					when "00110000010111101" => rgb <= "101000";
					when "00110000010111110" => rgb <= "101000";
					when "00110000010111111" => rgb <= "101000";
					when "00110000011000000" => rgb <= "101000";
					when "00110000011000001" => rgb <= "101000";
					when "00110000011000010" => rgb <= "101000";
					when "00110000011000011" => rgb <= "101000";
					when "00110000011000100" => rgb <= "101000";
					when "00110000011000101" => rgb <= "101000";
					when "00110000011000110" => rgb <= "111000";
					when "00110000011000111" => rgb <= "101000";
					when "00110000011001000" => rgb <= "101000";
					when "00110000011001001" => rgb <= "101000";
					when "00110000011001010" => rgb <= "101000";
					when "00110000011001011" => rgb <= "101000";
					when "00110000011001100" => rgb <= "101000";
					when "00110000011001101" => rgb <= "101000";
					when "00110000011001110" => rgb <= "101000";
					when "00110000011001111" => rgb <= "101000";
					when "00110000011010000" => rgb <= "101000";
					when "00110000011010001" => rgb <= "101000";
					when "00110000011010010" => rgb <= "101000";
					when "00110000011010011" => rgb <= "101000";
					when "00110000011010100" => rgb <= "101000";
					when "00110000011010101" => rgb <= "101000";
					when "00110000011010110" => rgb <= "101000";
					when "00110000011010111" => rgb <= "010100";
					when "00110000011011000" => rgb <= "000000";
					when "00110000011011001" => rgb <= "000000";
					when "00110000011011010" => rgb <= "000000";
					when "00110000011011011" => rgb <= "000000";
					when "00110000011011100" => rgb <= "000000";
					when "00110000011011101" => rgb <= "000000";
					when "00110000011011110" => rgb <= "000000";
					when "00110000011011111" => rgb <= "000000";
					when "00110000011100000" => rgb <= "000000";
					when "00110000011100001" => rgb <= "000000";
					when "00110000011100010" => rgb <= "000000";
					when "00110000011100011" => rgb <= "000000";
					when "00110000011100100" => rgb <= "000000";
					when "00110000011100101" => rgb <= "000000";
					when "00110000011100110" => rgb <= "000000";
					when "00110000011100111" => rgb <= "000000";
					when "00110000011101000" => rgb <= "000000";
					when "00110000011101001" => rgb <= "000000";
					when "00110000011101010" => rgb <= "000000";
					when "00110000011101011" => rgb <= "000000";
					when "00110000011101100" => rgb <= "000000";
					when "00110000011101101" => rgb <= "000000";
					when "00110000011101110" => rgb <= "000000";
					when "00110000011101111" => rgb <= "000000";
					when "00110000011110000" => rgb <= "000000";
					when "00110000011110001" => rgb <= "000000";
					when "00110000011110010" => rgb <= "000000";
					when "00110000011110011" => rgb <= "000000";
					when "00110000011110100" => rgb <= "000000";
					when "00110000011110101" => rgb <= "000000";
					when "00110000011110110" => rgb <= "000000";
					when "00110000011110111" => rgb <= "000000";
					when "00110000011111000" => rgb <= "000000";
					when "00110000011111001" => rgb <= "000000";
					when "00110000011111010" => rgb <= "000000";
					when "00110000011111011" => rgb <= "000000";
					when "00110000011111100" => rgb <= "000000";
					when "00110000011111101" => rgb <= "000000";
					when "00110000011111110" => rgb <= "000000";
					when "00110000011111111" => rgb <= "000000";
					when "00110000100000000" => rgb <= "000000";
					when "00110000100000001" => rgb <= "000000";
					when "00110000100000010" => rgb <= "000000";
					when "00110000100000011" => rgb <= "000000";
					when "00110000100000100" => rgb <= "000000";
					when "00110000100000101" => rgb <= "000000";
					when "00110000100000110" => rgb <= "000000";
					when "00110000100000111" => rgb <= "000000";
					when "00110000100001000" => rgb <= "000000";
					when "00110000100001001" => rgb <= "000000";
					when "00110000100001010" => rgb <= "000000";
					when "00110000100001011" => rgb <= "000000";
					when "00110000100001100" => rgb <= "000000";
					when "00110000100001101" => rgb <= "000000";
					when "00110000100001110" => rgb <= "000000";
					when "00110000100001111" => rgb <= "000000";
					when "00110000100010000" => rgb <= "000000";
					when "00110000100010001" => rgb <= "000000";
					when "00110000100010010" => rgb <= "000000";
					when "00110000100010011" => rgb <= "000000";
					when "00110000100010100" => rgb <= "000000";
					when "00110000100010101" => rgb <= "000000";
					when "00110000100010110" => rgb <= "000000";
					when "00110000100010111" => rgb <= "000000";
					when "00110000100011000" => rgb <= "000000";
					when "00110000100011001" => rgb <= "000000";
					when "00110000100011010" => rgb <= "000000";
					when "00110000100011011" => rgb <= "000000";
					when "00110000100011100" => rgb <= "000000";
					when "00110000100011101" => rgb <= "000000";
					when "00110000100011110" => rgb <= "000000";
					when "00110000100011111" => rgb <= "000000";
					when "00110000100100000" => rgb <= "000000";
					when "00110000100100001" => rgb <= "000000";
					when "00110000100100010" => rgb <= "000000";
					when "00110000100100011" => rgb <= "000000";
					when "00110000100100100" => rgb <= "000000";
					when "00110000100100101" => rgb <= "000000";
					when "00110000100100110" => rgb <= "000000";
					when "00110000100100111" => rgb <= "000000";
					when "00110000100101000" => rgb <= "000000";
					when "00110000100101001" => rgb <= "000000";
					when "00110000100101010" => rgb <= "000000";
					when "00110000100101011" => rgb <= "000000";
					when "00110000100101100" => rgb <= "000000";
					when "00110000100101101" => rgb <= "000000";
					when "00110000100101110" => rgb <= "000000";
					when "00110000100101111" => rgb <= "000000";
					when "00110000100110000" => rgb <= "000000";
					when "00110000100110001" => rgb <= "000000";
					when "00110000100110010" => rgb <= "000000";
					when "00110000100110011" => rgb <= "000000";
					when "00110000100110100" => rgb <= "000000";
					when "00110000100110101" => rgb <= "000000";
					when "00110000100110110" => rgb <= "000000";
					when "00110000100110111" => rgb <= "000000";
					when "00110000100111000" => rgb <= "000000";
					when "00110000100111001" => rgb <= "000000";
					when "00110000100111010" => rgb <= "000000";
					when "00110000100111011" => rgb <= "000000";
					when "00110000100111100" => rgb <= "000000";
					when "00110000100111101" => rgb <= "000000";
					when "00110000100111110" => rgb <= "000000";
					when "00110000100111111" => rgb <= "000000";
					when "00110001000000000" => rgb <= "000000";
					when "00110001000000001" => rgb <= "000000";
					when "00110001000000010" => rgb <= "000000";
					when "00110001000000011" => rgb <= "000000";
					when "00110001000000100" => rgb <= "000000";
					when "00110001000000101" => rgb <= "000000";
					when "00110001000000110" => rgb <= "000000";
					when "00110001000000111" => rgb <= "000000";
					when "00110001000001000" => rgb <= "000000";
					when "00110001000001001" => rgb <= "000000";
					when "00110001000001010" => rgb <= "000000";
					when "00110001000001011" => rgb <= "000000";
					when "00110001000001100" => rgb <= "000000";
					when "00110001000001101" => rgb <= "000000";
					when "00110001000001110" => rgb <= "000000";
					when "00110001000001111" => rgb <= "000000";
					when "00110001000010000" => rgb <= "000000";
					when "00110001000010001" => rgb <= "000000";
					when "00110001000010010" => rgb <= "000000";
					when "00110001000010011" => rgb <= "000000";
					when "00110001000010100" => rgb <= "000000";
					when "00110001000010101" => rgb <= "000000";
					when "00110001000010110" => rgb <= "000000";
					when "00110001000010111" => rgb <= "000000";
					when "00110001000011000" => rgb <= "000000";
					when "00110001000011001" => rgb <= "000000";
					when "00110001000011010" => rgb <= "000000";
					when "00110001000011011" => rgb <= "000000";
					when "00110001000011100" => rgb <= "000000";
					when "00110001000011101" => rgb <= "000000";
					when "00110001000011110" => rgb <= "000000";
					when "00110001000011111" => rgb <= "000000";
					when "00110001000100000" => rgb <= "000000";
					when "00110001000100001" => rgb <= "000000";
					when "00110001000100010" => rgb <= "000000";
					when "00110001000100011" => rgb <= "000000";
					when "00110001000100100" => rgb <= "000000";
					when "00110001000100101" => rgb <= "000000";
					when "00110001000100110" => rgb <= "000000";
					when "00110001000100111" => rgb <= "000000";
					when "00110001000101000" => rgb <= "000000";
					when "00110001000101001" => rgb <= "000000";
					when "00110001000101010" => rgb <= "000000";
					when "00110001000101011" => rgb <= "000000";
					when "00110001000101100" => rgb <= "000000";
					when "00110001000101101" => rgb <= "000000";
					when "00110001000101110" => rgb <= "000000";
					when "00110001000101111" => rgb <= "000000";
					when "00110001000110000" => rgb <= "000000";
					when "00110001000110001" => rgb <= "000000";
					when "00110001000110010" => rgb <= "000000";
					when "00110001000110011" => rgb <= "000000";
					when "00110001000110100" => rgb <= "000000";
					when "00110001000110101" => rgb <= "000000";
					when "00110001000110110" => rgb <= "000000";
					when "00110001000110111" => rgb <= "000000";
					when "00110001000111000" => rgb <= "000000";
					when "00110001000111001" => rgb <= "000000";
					when "00110001000111010" => rgb <= "000000";
					when "00110001000111011" => rgb <= "000000";
					when "00110001000111100" => rgb <= "000000";
					when "00110001000111101" => rgb <= "000000";
					when "00110001000111110" => rgb <= "000000";
					when "00110001000111111" => rgb <= "000000";
					when "00110001001000000" => rgb <= "000000";
					when "00110001001000001" => rgb <= "000000";
					when "00110001001000010" => rgb <= "000000";
					when "00110001001000011" => rgb <= "000000";
					when "00110001001000100" => rgb <= "000000";
					when "00110001001000101" => rgb <= "000000";
					when "00110001001000110" => rgb <= "000000";
					when "00110001001000111" => rgb <= "000000";
					when "00110001001001000" => rgb <= "000000";
					when "00110001001001001" => rgb <= "000000";
					when "00110001001001010" => rgb <= "000000";
					when "00110001001001011" => rgb <= "000000";
					when "00110001001001100" => rgb <= "000000";
					when "00110001001001101" => rgb <= "000000";
					when "00110001001001110" => rgb <= "000000";
					when "00110001001001111" => rgb <= "000000";
					when "00110001001010000" => rgb <= "000000";
					when "00110001001010001" => rgb <= "000000";
					when "00110001001010010" => rgb <= "000000";
					when "00110001001010011" => rgb <= "000000";
					when "00110001001010100" => rgb <= "000000";
					when "00110001001010101" => rgb <= "000000";
					when "00110001001010110" => rgb <= "000000";
					when "00110001001010111" => rgb <= "000000";
					when "00110001001011000" => rgb <= "000000";
					when "00110001001011001" => rgb <= "000000";
					when "00110001001011010" => rgb <= "000000";
					when "00110001001011011" => rgb <= "000000";
					when "00110001001011100" => rgb <= "000000";
					when "00110001001011101" => rgb <= "000000";
					when "00110001001011110" => rgb <= "000000";
					when "00110001001011111" => rgb <= "000000";
					when "00110001001100000" => rgb <= "000000";
					when "00110001001100001" => rgb <= "000000";
					when "00110001001100010" => rgb <= "000000";
					when "00110001001100011" => rgb <= "000000";
					when "00110001001100100" => rgb <= "000000";
					when "00110001001100101" => rgb <= "000000";
					when "00110001001100110" => rgb <= "010100";
					when "00110001001100111" => rgb <= "111000";
					when "00110001001101000" => rgb <= "101000";
					when "00110001001101001" => rgb <= "101000";
					when "00110001001101010" => rgb <= "101000";
					when "00110001001101011" => rgb <= "101000";
					when "00110001001101100" => rgb <= "101000";
					when "00110001001101101" => rgb <= "101000";
					when "00110001001101110" => rgb <= "101000";
					when "00110001001101111" => rgb <= "101000";
					when "00110001001110000" => rgb <= "101000";
					when "00110001001110001" => rgb <= "101000";
					when "00110001001110010" => rgb <= "101000";
					when "00110001001110011" => rgb <= "101000";
					when "00110001001110100" => rgb <= "101000";
					when "00110001001110101" => rgb <= "101000";
					when "00110001001110110" => rgb <= "101000";
					when "00110001001110111" => rgb <= "101000";
					when "00110001001111000" => rgb <= "101000";
					when "00110001001111001" => rgb <= "101000";
					when "00110001001111010" => rgb <= "101000";
					when "00110001001111011" => rgb <= "101000";
					when "00110001001111100" => rgb <= "101000";
					when "00110001001111101" => rgb <= "101000";
					when "00110001001111110" => rgb <= "101000";
					when "00110001001111111" => rgb <= "101000";
					when "00110001010000000" => rgb <= "101000";
					when "00110001010000001" => rgb <= "101000";
					when "00110001010000010" => rgb <= "101000";
					when "00110001010000011" => rgb <= "101000";
					when "00110001010000100" => rgb <= "101000";
					when "00110001010000101" => rgb <= "101000";
					when "00110001010000110" => rgb <= "101000";
					when "00110001010000111" => rgb <= "101000";
					when "00110001010001000" => rgb <= "101001";
					when "00110001010001001" => rgb <= "101001";
					when "00110001010001010" => rgb <= "101001";
					when "00110001010001011" => rgb <= "101001";
					when "00110001010001100" => rgb <= "101001";
					when "00110001010001101" => rgb <= "101001";
					when "00110001010001110" => rgb <= "101001";
					when "00110001010001111" => rgb <= "101001";
					when "00110001010010000" => rgb <= "101001";
					when "00110001010010001" => rgb <= "111010";
					when "00110001010010010" => rgb <= "111001";
					when "00110001010010011" => rgb <= "101001";
					when "00110001010010100" => rgb <= "101001";
					when "00110001010010101" => rgb <= "101000";
					when "00110001010010110" => rgb <= "101000";
					when "00110001010010111" => rgb <= "101000";
					when "00110001010011000" => rgb <= "101000";
					when "00110001010011001" => rgb <= "101000";
					when "00110001010011010" => rgb <= "101000";
					when "00110001010011011" => rgb <= "101000";
					when "00110001010011100" => rgb <= "101000";
					when "00110001010011101" => rgb <= "101000";
					when "00110001010011110" => rgb <= "101000";
					when "00110001010011111" => rgb <= "101000";
					when "00110001010100000" => rgb <= "101000";
					when "00110001010100001" => rgb <= "101000";
					when "00110001010100010" => rgb <= "101000";
					when "00110001010100011" => rgb <= "101000";
					when "00110001010100100" => rgb <= "101000";
					when "00110001010100101" => rgb <= "101000";
					when "00110001010100110" => rgb <= "101000";
					when "00110001010100111" => rgb <= "101000";
					when "00110001010101000" => rgb <= "101000";
					when "00110001010101001" => rgb <= "101000";
					when "00110001010101010" => rgb <= "101000";
					when "00110001010101011" => rgb <= "101000";
					when "00110001010101100" => rgb <= "101000";
					when "00110001010101101" => rgb <= "101000";
					when "00110001010101110" => rgb <= "101000";
					when "00110001010101111" => rgb <= "101000";
					when "00110001010110000" => rgb <= "101000";
					when "00110001010110001" => rgb <= "101000";
					when "00110001010110010" => rgb <= "101000";
					when "00110001010110011" => rgb <= "101000";
					when "00110001010110100" => rgb <= "101000";
					when "00110001010110101" => rgb <= "101000";
					when "00110001010110110" => rgb <= "101000";
					when "00110001010110111" => rgb <= "101000";
					when "00110001010111000" => rgb <= "101000";
					when "00110001010111001" => rgb <= "101000";
					when "00110001010111010" => rgb <= "101000";
					when "00110001010111011" => rgb <= "101000";
					when "00110001010111100" => rgb <= "101000";
					when "00110001010111101" => rgb <= "101000";
					when "00110001010111110" => rgb <= "101000";
					when "00110001010111111" => rgb <= "101000";
					when "00110001011000000" => rgb <= "101000";
					when "00110001011000001" => rgb <= "101001";
					when "00110001011000010" => rgb <= "101000";
					when "00110001011000011" => rgb <= "101000";
					when "00110001011000100" => rgb <= "101000";
					when "00110001011000101" => rgb <= "111001";
					when "00110001011000110" => rgb <= "101000";
					when "00110001011000111" => rgb <= "101000";
					when "00110001011001000" => rgb <= "101001";
					when "00110001011001001" => rgb <= "101000";
					when "00110001011001010" => rgb <= "101000";
					when "00110001011001011" => rgb <= "101000";
					when "00110001011001100" => rgb <= "101000";
					when "00110001011001101" => rgb <= "101000";
					when "00110001011001110" => rgb <= "101000";
					when "00110001011001111" => rgb <= "101000";
					when "00110001011010000" => rgb <= "101000";
					when "00110001011010001" => rgb <= "101000";
					when "00110001011010010" => rgb <= "101000";
					when "00110001011010011" => rgb <= "101000";
					when "00110001011010100" => rgb <= "101000";
					when "00110001011010101" => rgb <= "101000";
					when "00110001011010110" => rgb <= "101000";
					when "00110001011010111" => rgb <= "010100";
					when "00110001011011000" => rgb <= "000000";
					when "00110001011011001" => rgb <= "000000";
					when "00110001011011010" => rgb <= "000000";
					when "00110001011011011" => rgb <= "000000";
					when "00110001011011100" => rgb <= "000000";
					when "00110001011011101" => rgb <= "000000";
					when "00110001011011110" => rgb <= "000000";
					when "00110001011011111" => rgb <= "000000";
					when "00110001011100000" => rgb <= "000000";
					when "00110001011100001" => rgb <= "000000";
					when "00110001011100010" => rgb <= "000000";
					when "00110001011100011" => rgb <= "000000";
					when "00110001011100100" => rgb <= "000000";
					when "00110001011100101" => rgb <= "000000";
					when "00110001011100110" => rgb <= "000000";
					when "00110001011100111" => rgb <= "000000";
					when "00110001011101000" => rgb <= "000000";
					when "00110001011101001" => rgb <= "000000";
					when "00110001011101010" => rgb <= "000000";
					when "00110001011101011" => rgb <= "000000";
					when "00110001011101100" => rgb <= "000000";
					when "00110001011101101" => rgb <= "000000";
					when "00110001011101110" => rgb <= "000000";
					when "00110001011101111" => rgb <= "000000";
					when "00110001011110000" => rgb <= "000000";
					when "00110001011110001" => rgb <= "000000";
					when "00110001011110010" => rgb <= "000000";
					when "00110001011110011" => rgb <= "000000";
					when "00110001011110100" => rgb <= "000000";
					when "00110001011110101" => rgb <= "000000";
					when "00110001011110110" => rgb <= "000000";
					when "00110001011110111" => rgb <= "000000";
					when "00110001011111000" => rgb <= "000000";
					when "00110001011111001" => rgb <= "000000";
					when "00110001011111010" => rgb <= "000000";
					when "00110001011111011" => rgb <= "000000";
					when "00110001011111100" => rgb <= "000000";
					when "00110001011111101" => rgb <= "000000";
					when "00110001011111110" => rgb <= "000000";
					when "00110001011111111" => rgb <= "000000";
					when "00110001100000000" => rgb <= "000000";
					when "00110001100000001" => rgb <= "000000";
					when "00110001100000010" => rgb <= "000000";
					when "00110001100000011" => rgb <= "000000";
					when "00110001100000100" => rgb <= "000000";
					when "00110001100000101" => rgb <= "000000";
					when "00110001100000110" => rgb <= "000000";
					when "00110001100000111" => rgb <= "000000";
					when "00110001100001000" => rgb <= "000000";
					when "00110001100001001" => rgb <= "000000";
					when "00110001100001010" => rgb <= "000000";
					when "00110001100001011" => rgb <= "000000";
					when "00110001100001100" => rgb <= "000000";
					when "00110001100001101" => rgb <= "000000";
					when "00110001100001110" => rgb <= "000000";
					when "00110001100001111" => rgb <= "000000";
					when "00110001100010000" => rgb <= "000000";
					when "00110001100010001" => rgb <= "000000";
					when "00110001100010010" => rgb <= "000000";
					when "00110001100010011" => rgb <= "000000";
					when "00110001100010100" => rgb <= "000000";
					when "00110001100010101" => rgb <= "000000";
					when "00110001100010110" => rgb <= "000000";
					when "00110001100010111" => rgb <= "000000";
					when "00110001100011000" => rgb <= "000000";
					when "00110001100011001" => rgb <= "000000";
					when "00110001100011010" => rgb <= "000000";
					when "00110001100011011" => rgb <= "000000";
					when "00110001100011100" => rgb <= "000000";
					when "00110001100011101" => rgb <= "000000";
					when "00110001100011110" => rgb <= "000000";
					when "00110001100011111" => rgb <= "000000";
					when "00110001100100000" => rgb <= "000000";
					when "00110001100100001" => rgb <= "000000";
					when "00110001100100010" => rgb <= "000000";
					when "00110001100100011" => rgb <= "000000";
					when "00110001100100100" => rgb <= "000000";
					when "00110001100100101" => rgb <= "000000";
					when "00110001100100110" => rgb <= "000000";
					when "00110001100100111" => rgb <= "000000";
					when "00110001100101000" => rgb <= "000000";
					when "00110001100101001" => rgb <= "000000";
					when "00110001100101010" => rgb <= "000000";
					when "00110001100101011" => rgb <= "000000";
					when "00110001100101100" => rgb <= "000000";
					when "00110001100101101" => rgb <= "000000";
					when "00110001100101110" => rgb <= "000000";
					when "00110001100101111" => rgb <= "000000";
					when "00110001100110000" => rgb <= "000000";
					when "00110001100110001" => rgb <= "000000";
					when "00110001100110010" => rgb <= "000000";
					when "00110001100110011" => rgb <= "000000";
					when "00110001100110100" => rgb <= "000000";
					when "00110001100110101" => rgb <= "000000";
					when "00110001100110110" => rgb <= "000000";
					when "00110001100110111" => rgb <= "000000";
					when "00110001100111000" => rgb <= "000000";
					when "00110001100111001" => rgb <= "000000";
					when "00110001100111010" => rgb <= "000000";
					when "00110001100111011" => rgb <= "000000";
					when "00110001100111100" => rgb <= "000000";
					when "00110001100111101" => rgb <= "000000";
					when "00110001100111110" => rgb <= "000000";
					when "00110001100111111" => rgb <= "000000";
					when "00110010000000000" => rgb <= "000000";
					when "00110010000000001" => rgb <= "000000";
					when "00110010000000010" => rgb <= "000000";
					when "00110010000000011" => rgb <= "000000";
					when "00110010000000100" => rgb <= "000000";
					when "00110010000000101" => rgb <= "000000";
					when "00110010000000110" => rgb <= "000000";
					when "00110010000000111" => rgb <= "000000";
					when "00110010000001000" => rgb <= "000000";
					when "00110010000001001" => rgb <= "000000";
					when "00110010000001010" => rgb <= "000000";
					when "00110010000001011" => rgb <= "000000";
					when "00110010000001100" => rgb <= "000000";
					when "00110010000001101" => rgb <= "000000";
					when "00110010000001110" => rgb <= "000000";
					when "00110010000001111" => rgb <= "000000";
					when "00110010000010000" => rgb <= "000000";
					when "00110010000010001" => rgb <= "000000";
					when "00110010000010010" => rgb <= "000000";
					when "00110010000010011" => rgb <= "000000";
					when "00110010000010100" => rgb <= "000000";
					when "00110010000010101" => rgb <= "000000";
					when "00110010000010110" => rgb <= "000000";
					when "00110010000010111" => rgb <= "000000";
					when "00110010000011000" => rgb <= "000000";
					when "00110010000011001" => rgb <= "000000";
					when "00110010000011010" => rgb <= "000000";
					when "00110010000011011" => rgb <= "000000";
					when "00110010000011100" => rgb <= "000000";
					when "00110010000011101" => rgb <= "000000";
					when "00110010000011110" => rgb <= "000000";
					when "00110010000011111" => rgb <= "000000";
					when "00110010000100000" => rgb <= "000000";
					when "00110010000100001" => rgb <= "000000";
					when "00110010000100010" => rgb <= "000000";
					when "00110010000100011" => rgb <= "000000";
					when "00110010000100100" => rgb <= "000000";
					when "00110010000100101" => rgb <= "000000";
					when "00110010000100110" => rgb <= "000000";
					when "00110010000100111" => rgb <= "000000";
					when "00110010000101000" => rgb <= "000000";
					when "00110010000101001" => rgb <= "000000";
					when "00110010000101010" => rgb <= "000000";
					when "00110010000101011" => rgb <= "000000";
					when "00110010000101100" => rgb <= "000000";
					when "00110010000101101" => rgb <= "000000";
					when "00110010000101110" => rgb <= "000000";
					when "00110010000101111" => rgb <= "000000";
					when "00110010000110000" => rgb <= "000000";
					when "00110010000110001" => rgb <= "000000";
					when "00110010000110010" => rgb <= "000000";
					when "00110010000110011" => rgb <= "000000";
					when "00110010000110100" => rgb <= "000000";
					when "00110010000110101" => rgb <= "000000";
					when "00110010000110110" => rgb <= "000000";
					when "00110010000110111" => rgb <= "000000";
					when "00110010000111000" => rgb <= "000000";
					when "00110010000111001" => rgb <= "000000";
					when "00110010000111010" => rgb <= "000000";
					when "00110010000111011" => rgb <= "000000";
					when "00110010000111100" => rgb <= "000000";
					when "00110010000111101" => rgb <= "000000";
					when "00110010000111110" => rgb <= "000000";
					when "00110010000111111" => rgb <= "000000";
					when "00110010001000000" => rgb <= "000000";
					when "00110010001000001" => rgb <= "000000";
					when "00110010001000010" => rgb <= "000000";
					when "00110010001000011" => rgb <= "000000";
					when "00110010001000100" => rgb <= "000000";
					when "00110010001000101" => rgb <= "000000";
					when "00110010001000110" => rgb <= "000000";
					when "00110010001000111" => rgb <= "000000";
					when "00110010001001000" => rgb <= "000000";
					when "00110010001001001" => rgb <= "000000";
					when "00110010001001010" => rgb <= "000000";
					when "00110010001001011" => rgb <= "000000";
					when "00110010001001100" => rgb <= "000000";
					when "00110010001001101" => rgb <= "000000";
					when "00110010001001110" => rgb <= "000000";
					when "00110010001001111" => rgb <= "000000";
					when "00110010001010000" => rgb <= "000000";
					when "00110010001010001" => rgb <= "000000";
					when "00110010001010010" => rgb <= "000000";
					when "00110010001010011" => rgb <= "000000";
					when "00110010001010100" => rgb <= "000000";
					when "00110010001010101" => rgb <= "000000";
					when "00110010001010110" => rgb <= "000000";
					when "00110010001010111" => rgb <= "000000";
					when "00110010001011000" => rgb <= "000000";
					when "00110010001011001" => rgb <= "000000";
					when "00110010001011010" => rgb <= "000000";
					when "00110010001011011" => rgb <= "000000";
					when "00110010001011100" => rgb <= "000000";
					when "00110010001011101" => rgb <= "000000";
					when "00110010001011110" => rgb <= "000000";
					when "00110010001011111" => rgb <= "000000";
					when "00110010001100000" => rgb <= "000000";
					when "00110010001100001" => rgb <= "000000";
					when "00110010001100010" => rgb <= "000000";
					when "00110010001100011" => rgb <= "000000";
					when "00110010001100100" => rgb <= "000000";
					when "00110010001100101" => rgb <= "000000";
					when "00110010001100110" => rgb <= "010100";
					when "00110010001100111" => rgb <= "111000";
					when "00110010001101000" => rgb <= "101000";
					when "00110010001101001" => rgb <= "101000";
					when "00110010001101010" => rgb <= "101000";
					when "00110010001101011" => rgb <= "101000";
					when "00110010001101100" => rgb <= "101000";
					when "00110010001101101" => rgb <= "101000";
					when "00110010001101110" => rgb <= "101000";
					when "00110010001101111" => rgb <= "101000";
					when "00110010001110000" => rgb <= "101000";
					when "00110010001110001" => rgb <= "101000";
					when "00110010001110010" => rgb <= "101000";
					when "00110010001110011" => rgb <= "101000";
					when "00110010001110100" => rgb <= "101000";
					when "00110010001110101" => rgb <= "101000";
					when "00110010001110110" => rgb <= "101000";
					when "00110010001110111" => rgb <= "101000";
					when "00110010001111000" => rgb <= "101000";
					when "00110010001111001" => rgb <= "101000";
					when "00110010001111010" => rgb <= "101000";
					when "00110010001111011" => rgb <= "101000";
					when "00110010001111100" => rgb <= "101000";
					when "00110010001111101" => rgb <= "101000";
					when "00110010001111110" => rgb <= "101000";
					when "00110010001111111" => rgb <= "101000";
					when "00110010010000000" => rgb <= "101000";
					when "00110010010000001" => rgb <= "101000";
					when "00110010010000010" => rgb <= "101000";
					when "00110010010000011" => rgb <= "101000";
					when "00110010010000100" => rgb <= "101000";
					when "00110010010000101" => rgb <= "101000";
					when "00110010010000110" => rgb <= "101000";
					when "00110010010000111" => rgb <= "101000";
					when "00110010010001000" => rgb <= "101001";
					when "00110010010001001" => rgb <= "101001";
					when "00110010010001010" => rgb <= "101001";
					when "00110010010001011" => rgb <= "101001";
					when "00110010010001100" => rgb <= "101001";
					when "00110010010001101" => rgb <= "111001";
					when "00110010010001110" => rgb <= "101001";
					when "00110010010001111" => rgb <= "101001";
					when "00110010010010000" => rgb <= "101001";
					when "00110010010010001" => rgb <= "101001";
					when "00110010010010010" => rgb <= "111001";
					when "00110010010010011" => rgb <= "101001";
					when "00110010010010100" => rgb <= "101000";
					when "00110010010010101" => rgb <= "101000";
					when "00110010010010110" => rgb <= "101000";
					when "00110010010010111" => rgb <= "101000";
					when "00110010010011000" => rgb <= "101000";
					when "00110010010011001" => rgb <= "101000";
					when "00110010010011010" => rgb <= "101000";
					when "00110010010011011" => rgb <= "101000";
					when "00110010010011100" => rgb <= "101000";
					when "00110010010011101" => rgb <= "101000";
					when "00110010010011110" => rgb <= "101000";
					when "00110010010011111" => rgb <= "101000";
					when "00110010010100000" => rgb <= "101000";
					when "00110010010100001" => rgb <= "101000";
					when "00110010010100010" => rgb <= "101000";
					when "00110010010100011" => rgb <= "101000";
					when "00110010010100100" => rgb <= "101000";
					when "00110010010100101" => rgb <= "101000";
					when "00110010010100110" => rgb <= "101000";
					when "00110010010100111" => rgb <= "101000";
					when "00110010010101000" => rgb <= "101000";
					when "00110010010101001" => rgb <= "101000";
					when "00110010010101010" => rgb <= "101000";
					when "00110010010101011" => rgb <= "101000";
					when "00110010010101100" => rgb <= "101000";
					when "00110010010101101" => rgb <= "101000";
					when "00110010010101110" => rgb <= "101000";
					when "00110010010101111" => rgb <= "101000";
					when "00110010010110000" => rgb <= "101000";
					when "00110010010110001" => rgb <= "101000";
					when "00110010010110010" => rgb <= "101000";
					when "00110010010110011" => rgb <= "101000";
					when "00110010010110100" => rgb <= "101000";
					when "00110010010110101" => rgb <= "101000";
					when "00110010010110110" => rgb <= "101000";
					when "00110010010110111" => rgb <= "101000";
					when "00110010010111000" => rgb <= "101000";
					when "00110010010111001" => rgb <= "101000";
					when "00110010010111010" => rgb <= "101000";
					when "00110010010111011" => rgb <= "101000";
					when "00110010010111100" => rgb <= "101000";
					when "00110010010111101" => rgb <= "101000";
					when "00110010010111110" => rgb <= "101000";
					when "00110010010111111" => rgb <= "101000";
					when "00110010011000000" => rgb <= "101000";
					when "00110010011000001" => rgb <= "101000";
					when "00110010011000010" => rgb <= "101001";
					when "00110010011000011" => rgb <= "101000";
					when "00110010011000100" => rgb <= "101000";
					when "00110010011000101" => rgb <= "101000";
					when "00110010011000110" => rgb <= "101000";
					when "00110010011000111" => rgb <= "101000";
					when "00110010011001000" => rgb <= "101000";
					when "00110010011001001" => rgb <= "101000";
					when "00110010011001010" => rgb <= "101000";
					when "00110010011001011" => rgb <= "101000";
					when "00110010011001100" => rgb <= "101000";
					when "00110010011001101" => rgb <= "101000";
					when "00110010011001110" => rgb <= "101000";
					when "00110010011001111" => rgb <= "101000";
					when "00110010011010000" => rgb <= "101000";
					when "00110010011010001" => rgb <= "101000";
					when "00110010011010010" => rgb <= "101000";
					when "00110010011010011" => rgb <= "101000";
					when "00110010011010100" => rgb <= "101000";
					when "00110010011010101" => rgb <= "101000";
					when "00110010011010110" => rgb <= "101000";
					when "00110010011010111" => rgb <= "010100";
					when "00110010011011000" => rgb <= "000000";
					when "00110010011011001" => rgb <= "000000";
					when "00110010011011010" => rgb <= "000000";
					when "00110010011011011" => rgb <= "000000";
					when "00110010011011100" => rgb <= "000000";
					when "00110010011011101" => rgb <= "000000";
					when "00110010011011110" => rgb <= "000000";
					when "00110010011011111" => rgb <= "000000";
					when "00110010011100000" => rgb <= "000000";
					when "00110010011100001" => rgb <= "000000";
					when "00110010011100010" => rgb <= "000000";
					when "00110010011100011" => rgb <= "000000";
					when "00110010011100100" => rgb <= "000000";
					when "00110010011100101" => rgb <= "000000";
					when "00110010011100110" => rgb <= "000000";
					when "00110010011100111" => rgb <= "000000";
					when "00110010011101000" => rgb <= "000000";
					when "00110010011101001" => rgb <= "000000";
					when "00110010011101010" => rgb <= "000000";
					when "00110010011101011" => rgb <= "000000";
					when "00110010011101100" => rgb <= "000000";
					when "00110010011101101" => rgb <= "000000";
					when "00110010011101110" => rgb <= "000000";
					when "00110010011101111" => rgb <= "000000";
					when "00110010011110000" => rgb <= "000000";
					when "00110010011110001" => rgb <= "000000";
					when "00110010011110010" => rgb <= "000000";
					when "00110010011110011" => rgb <= "000000";
					when "00110010011110100" => rgb <= "000000";
					when "00110010011110101" => rgb <= "000000";
					when "00110010011110110" => rgb <= "000000";
					when "00110010011110111" => rgb <= "000000";
					when "00110010011111000" => rgb <= "000000";
					when "00110010011111001" => rgb <= "000000";
					when "00110010011111010" => rgb <= "000000";
					when "00110010011111011" => rgb <= "000000";
					when "00110010011111100" => rgb <= "000000";
					when "00110010011111101" => rgb <= "000000";
					when "00110010011111110" => rgb <= "000000";
					when "00110010011111111" => rgb <= "000000";
					when "00110010100000000" => rgb <= "000000";
					when "00110010100000001" => rgb <= "000000";
					when "00110010100000010" => rgb <= "000000";
					when "00110010100000011" => rgb <= "000000";
					when "00110010100000100" => rgb <= "000000";
					when "00110010100000101" => rgb <= "000000";
					when "00110010100000110" => rgb <= "000000";
					when "00110010100000111" => rgb <= "000000";
					when "00110010100001000" => rgb <= "000000";
					when "00110010100001001" => rgb <= "000000";
					when "00110010100001010" => rgb <= "000000";
					when "00110010100001011" => rgb <= "000000";
					when "00110010100001100" => rgb <= "000000";
					when "00110010100001101" => rgb <= "000000";
					when "00110010100001110" => rgb <= "000000";
					when "00110010100001111" => rgb <= "000000";
					when "00110010100010000" => rgb <= "000000";
					when "00110010100010001" => rgb <= "000000";
					when "00110010100010010" => rgb <= "000000";
					when "00110010100010011" => rgb <= "000000";
					when "00110010100010100" => rgb <= "000000";
					when "00110010100010101" => rgb <= "000000";
					when "00110010100010110" => rgb <= "000000";
					when "00110010100010111" => rgb <= "000000";
					when "00110010100011000" => rgb <= "000000";
					when "00110010100011001" => rgb <= "000000";
					when "00110010100011010" => rgb <= "000000";
					when "00110010100011011" => rgb <= "000000";
					when "00110010100011100" => rgb <= "000000";
					when "00110010100011101" => rgb <= "000000";
					when "00110010100011110" => rgb <= "000000";
					when "00110010100011111" => rgb <= "000000";
					when "00110010100100000" => rgb <= "000000";
					when "00110010100100001" => rgb <= "000000";
					when "00110010100100010" => rgb <= "000000";
					when "00110010100100011" => rgb <= "000000";
					when "00110010100100100" => rgb <= "000000";
					when "00110010100100101" => rgb <= "000000";
					when "00110010100100110" => rgb <= "000000";
					when "00110010100100111" => rgb <= "000000";
					when "00110010100101000" => rgb <= "000000";
					when "00110010100101001" => rgb <= "000000";
					when "00110010100101010" => rgb <= "000000";
					when "00110010100101011" => rgb <= "000000";
					when "00110010100101100" => rgb <= "000000";
					when "00110010100101101" => rgb <= "000000";
					when "00110010100101110" => rgb <= "000000";
					when "00110010100101111" => rgb <= "000000";
					when "00110010100110000" => rgb <= "000000";
					when "00110010100110001" => rgb <= "000000";
					when "00110010100110010" => rgb <= "000000";
					when "00110010100110011" => rgb <= "000000";
					when "00110010100110100" => rgb <= "000000";
					when "00110010100110101" => rgb <= "000000";
					when "00110010100110110" => rgb <= "000000";
					when "00110010100110111" => rgb <= "000000";
					when "00110010100111000" => rgb <= "000000";
					when "00110010100111001" => rgb <= "000000";
					when "00110010100111010" => rgb <= "000000";
					when "00110010100111011" => rgb <= "000000";
					when "00110010100111100" => rgb <= "000000";
					when "00110010100111101" => rgb <= "000000";
					when "00110010100111110" => rgb <= "000000";
					when "00110010100111111" => rgb <= "000000";
					when "00110011000000000" => rgb <= "000000";
					when "00110011000000001" => rgb <= "000000";
					when "00110011000000010" => rgb <= "000000";
					when "00110011000000011" => rgb <= "000000";
					when "00110011000000100" => rgb <= "000000";
					when "00110011000000101" => rgb <= "000000";
					when "00110011000000110" => rgb <= "000000";
					when "00110011000000111" => rgb <= "000000";
					when "00110011000001000" => rgb <= "000000";
					when "00110011000001001" => rgb <= "000000";
					when "00110011000001010" => rgb <= "000000";
					when "00110011000001011" => rgb <= "000000";
					when "00110011000001100" => rgb <= "000000";
					when "00110011000001101" => rgb <= "000000";
					when "00110011000001110" => rgb <= "000000";
					when "00110011000001111" => rgb <= "000000";
					when "00110011000010000" => rgb <= "000000";
					when "00110011000010001" => rgb <= "000000";
					when "00110011000010010" => rgb <= "000000";
					when "00110011000010011" => rgb <= "000000";
					when "00110011000010100" => rgb <= "000000";
					when "00110011000010101" => rgb <= "000000";
					when "00110011000010110" => rgb <= "000000";
					when "00110011000010111" => rgb <= "000000";
					when "00110011000011000" => rgb <= "000000";
					when "00110011000011001" => rgb <= "000000";
					when "00110011000011010" => rgb <= "000000";
					when "00110011000011011" => rgb <= "000000";
					when "00110011000011100" => rgb <= "000000";
					when "00110011000011101" => rgb <= "000000";
					when "00110011000011110" => rgb <= "000000";
					when "00110011000011111" => rgb <= "000000";
					when "00110011000100000" => rgb <= "000000";
					when "00110011000100001" => rgb <= "000000";
					when "00110011000100010" => rgb <= "000000";
					when "00110011000100011" => rgb <= "000000";
					when "00110011000100100" => rgb <= "000000";
					when "00110011000100101" => rgb <= "000000";
					when "00110011000100110" => rgb <= "000000";
					when "00110011000100111" => rgb <= "000000";
					when "00110011000101000" => rgb <= "000000";
					when "00110011000101001" => rgb <= "000000";
					when "00110011000101010" => rgb <= "000000";
					when "00110011000101011" => rgb <= "000000";
					when "00110011000101100" => rgb <= "000000";
					when "00110011000101101" => rgb <= "000000";
					when "00110011000101110" => rgb <= "000000";
					when "00110011000101111" => rgb <= "000000";
					when "00110011000110000" => rgb <= "000000";
					when "00110011000110001" => rgb <= "000000";
					when "00110011000110010" => rgb <= "000000";
					when "00110011000110011" => rgb <= "000000";
					when "00110011000110100" => rgb <= "000000";
					when "00110011000110101" => rgb <= "000000";
					when "00110011000110110" => rgb <= "000000";
					when "00110011000110111" => rgb <= "000000";
					when "00110011000111000" => rgb <= "000000";
					when "00110011000111001" => rgb <= "000000";
					when "00110011000111010" => rgb <= "000000";
					when "00110011000111011" => rgb <= "000000";
					when "00110011000111100" => rgb <= "000000";
					when "00110011000111101" => rgb <= "000000";
					when "00110011000111110" => rgb <= "000000";
					when "00110011000111111" => rgb <= "000000";
					when "00110011001000000" => rgb <= "000000";
					when "00110011001000001" => rgb <= "000000";
					when "00110011001000010" => rgb <= "000000";
					when "00110011001000011" => rgb <= "000000";
					when "00110011001000100" => rgb <= "000000";
					when "00110011001000101" => rgb <= "000000";
					when "00110011001000110" => rgb <= "000000";
					when "00110011001000111" => rgb <= "000000";
					when "00110011001001000" => rgb <= "000000";
					when "00110011001001001" => rgb <= "000000";
					when "00110011001001010" => rgb <= "000000";
					when "00110011001001011" => rgb <= "000000";
					when "00110011001001100" => rgb <= "000000";
					when "00110011001001101" => rgb <= "000000";
					when "00110011001001110" => rgb <= "000000";
					when "00110011001001111" => rgb <= "000000";
					when "00110011001010000" => rgb <= "000000";
					when "00110011001010001" => rgb <= "000000";
					when "00110011001010010" => rgb <= "000000";
					when "00110011001010011" => rgb <= "000000";
					when "00110011001010100" => rgb <= "000000";
					when "00110011001010101" => rgb <= "000000";
					when "00110011001010110" => rgb <= "000000";
					when "00110011001010111" => rgb <= "000000";
					when "00110011001011000" => rgb <= "000000";
					when "00110011001011001" => rgb <= "000000";
					when "00110011001011010" => rgb <= "000000";
					when "00110011001011011" => rgb <= "000000";
					when "00110011001011100" => rgb <= "000000";
					when "00110011001011101" => rgb <= "000000";
					when "00110011001011110" => rgb <= "000000";
					when "00110011001011111" => rgb <= "000000";
					when "00110011001100000" => rgb <= "000000";
					when "00110011001100001" => rgb <= "000000";
					when "00110011001100010" => rgb <= "000000";
					when "00110011001100011" => rgb <= "000000";
					when "00110011001100100" => rgb <= "000000";
					when "00110011001100101" => rgb <= "000000";
					when "00110011001100110" => rgb <= "010100";
					when "00110011001100111" => rgb <= "111000";
					when "00110011001101000" => rgb <= "101000";
					when "00110011001101001" => rgb <= "101000";
					when "00110011001101010" => rgb <= "101000";
					when "00110011001101011" => rgb <= "101000";
					when "00110011001101100" => rgb <= "101000";
					when "00110011001101101" => rgb <= "101000";
					when "00110011001101110" => rgb <= "101000";
					when "00110011001101111" => rgb <= "101000";
					when "00110011001110000" => rgb <= "101000";
					when "00110011001110001" => rgb <= "100100";
					when "00110011001110010" => rgb <= "000000";
					when "00110011001110011" => rgb <= "000000";
					when "00110011001110100" => rgb <= "000000";
					when "00110011001110101" => rgb <= "000000";
					when "00110011001110110" => rgb <= "000000";
					when "00110011001110111" => rgb <= "000000";
					when "00110011001111000" => rgb <= "000000";
					when "00110011001111001" => rgb <= "000000";
					when "00110011001111010" => rgb <= "000000";
					when "00110011001111011" => rgb <= "000000";
					when "00110011001111100" => rgb <= "000000";
					when "00110011001111101" => rgb <= "101000";
					when "00110011001111110" => rgb <= "101000";
					when "00110011001111111" => rgb <= "101000";
					when "00110011010000000" => rgb <= "101000";
					when "00110011010000001" => rgb <= "101000";
					when "00110011010000010" => rgb <= "101000";
					when "00110011010000011" => rgb <= "101000";
					when "00110011010000100" => rgb <= "101000";
					when "00110011010000101" => rgb <= "101000";
					when "00110011010000110" => rgb <= "101000";
					when "00110011010000111" => rgb <= "101000";
					when "00110011010001000" => rgb <= "101000";
					when "00110011010001001" => rgb <= "101001";
					when "00110011010001010" => rgb <= "101001";
					when "00110011010001011" => rgb <= "101001";
					when "00110011010001100" => rgb <= "101001";
					when "00110011010001101" => rgb <= "101001";
					when "00110011010001110" => rgb <= "101001";
					when "00110011010001111" => rgb <= "101001";
					when "00110011010010000" => rgb <= "101000";
					when "00110011010010001" => rgb <= "101001";
					when "00110011010010010" => rgb <= "101001";
					when "00110011010010011" => rgb <= "101000";
					when "00110011010010100" => rgb <= "101000";
					when "00110011010010101" => rgb <= "101000";
					when "00110011010010110" => rgb <= "101000";
					when "00110011010010111" => rgb <= "101000";
					when "00110011010011000" => rgb <= "101000";
					when "00110011010011001" => rgb <= "101000";
					when "00110011010011010" => rgb <= "101000";
					when "00110011010011011" => rgb <= "101000";
					when "00110011010011100" => rgb <= "101000";
					when "00110011010011101" => rgb <= "101000";
					when "00110011010011110" => rgb <= "101000";
					when "00110011010011111" => rgb <= "101000";
					when "00110011010100000" => rgb <= "101000";
					when "00110011010100001" => rgb <= "101000";
					when "00110011010100010" => rgb <= "101000";
					when "00110011010100011" => rgb <= "101000";
					when "00110011010100100" => rgb <= "101000";
					when "00110011010100101" => rgb <= "101000";
					when "00110011010100110" => rgb <= "101000";
					when "00110011010100111" => rgb <= "101000";
					when "00110011010101000" => rgb <= "101000";
					when "00110011010101001" => rgb <= "101000";
					when "00110011010101010" => rgb <= "101000";
					when "00110011010101011" => rgb <= "101000";
					when "00110011010101100" => rgb <= "101000";
					when "00110011010101101" => rgb <= "101000";
					when "00110011010101110" => rgb <= "101000";
					when "00110011010101111" => rgb <= "101000";
					when "00110011010110000" => rgb <= "101000";
					when "00110011010110001" => rgb <= "101000";
					when "00110011010110010" => rgb <= "101000";
					when "00110011010110011" => rgb <= "101000";
					when "00110011010110100" => rgb <= "101000";
					when "00110011010110101" => rgb <= "101000";
					when "00110011010110110" => rgb <= "101000";
					when "00110011010110111" => rgb <= "101000";
					when "00110011010111000" => rgb <= "101000";
					when "00110011010111001" => rgb <= "101000";
					when "00110011010111010" => rgb <= "101000";
					when "00110011010111011" => rgb <= "101000";
					when "00110011010111100" => rgb <= "101000";
					when "00110011010111101" => rgb <= "101000";
					when "00110011010111110" => rgb <= "101000";
					when "00110011010111111" => rgb <= "101000";
					when "00110011011000000" => rgb <= "100100";
					when "00110011011000001" => rgb <= "000000";
					when "00110011011000010" => rgb <= "000000";
					when "00110011011000011" => rgb <= "000000";
					when "00110011011000100" => rgb <= "000000";
					when "00110011011000101" => rgb <= "000000";
					when "00110011011000110" => rgb <= "000000";
					when "00110011011000111" => rgb <= "000000";
					when "00110011011001000" => rgb <= "000000";
					when "00110011011001001" => rgb <= "000000";
					when "00110011011001010" => rgb <= "000000";
					when "00110011011001011" => rgb <= "000000";
					when "00110011011001100" => rgb <= "100100";
					when "00110011011001101" => rgb <= "101000";
					when "00110011011001110" => rgb <= "101000";
					when "00110011011001111" => rgb <= "101000";
					when "00110011011010000" => rgb <= "101000";
					when "00110011011010001" => rgb <= "101000";
					when "00110011011010010" => rgb <= "101000";
					when "00110011011010011" => rgb <= "101000";
					when "00110011011010100" => rgb <= "101000";
					when "00110011011010101" => rgb <= "101000";
					when "00110011011010110" => rgb <= "101000";
					when "00110011011010111" => rgb <= "010100";
					when "00110011011011000" => rgb <= "000000";
					when "00110011011011001" => rgb <= "000000";
					when "00110011011011010" => rgb <= "000000";
					when "00110011011011011" => rgb <= "000000";
					when "00110011011011100" => rgb <= "000000";
					when "00110011011011101" => rgb <= "000000";
					when "00110011011011110" => rgb <= "000000";
					when "00110011011011111" => rgb <= "000000";
					when "00110011011100000" => rgb <= "000000";
					when "00110011011100001" => rgb <= "000000";
					when "00110011011100010" => rgb <= "000000";
					when "00110011011100011" => rgb <= "000000";
					when "00110011011100100" => rgb <= "000000";
					when "00110011011100101" => rgb <= "000000";
					when "00110011011100110" => rgb <= "000000";
					when "00110011011100111" => rgb <= "000000";
					when "00110011011101000" => rgb <= "000000";
					when "00110011011101001" => rgb <= "000000";
					when "00110011011101010" => rgb <= "000000";
					when "00110011011101011" => rgb <= "000000";
					when "00110011011101100" => rgb <= "000000";
					when "00110011011101101" => rgb <= "000000";
					when "00110011011101110" => rgb <= "000000";
					when "00110011011101111" => rgb <= "000000";
					when "00110011011110000" => rgb <= "000000";
					when "00110011011110001" => rgb <= "000000";
					when "00110011011110010" => rgb <= "000000";
					when "00110011011110011" => rgb <= "000000";
					when "00110011011110100" => rgb <= "000000";
					when "00110011011110101" => rgb <= "000000";
					when "00110011011110110" => rgb <= "000000";
					when "00110011011110111" => rgb <= "000000";
					when "00110011011111000" => rgb <= "000000";
					when "00110011011111001" => rgb <= "000000";
					when "00110011011111010" => rgb <= "000000";
					when "00110011011111011" => rgb <= "000000";
					when "00110011011111100" => rgb <= "000000";
					when "00110011011111101" => rgb <= "000000";
					when "00110011011111110" => rgb <= "000000";
					when "00110011011111111" => rgb <= "000000";
					when "00110011100000000" => rgb <= "000000";
					when "00110011100000001" => rgb <= "000000";
					when "00110011100000010" => rgb <= "000000";
					when "00110011100000011" => rgb <= "000000";
					when "00110011100000100" => rgb <= "000000";
					when "00110011100000101" => rgb <= "000000";
					when "00110011100000110" => rgb <= "000000";
					when "00110011100000111" => rgb <= "000000";
					when "00110011100001000" => rgb <= "000000";
					when "00110011100001001" => rgb <= "000000";
					when "00110011100001010" => rgb <= "000000";
					when "00110011100001011" => rgb <= "000000";
					when "00110011100001100" => rgb <= "000000";
					when "00110011100001101" => rgb <= "000000";
					when "00110011100001110" => rgb <= "000000";
					when "00110011100001111" => rgb <= "000000";
					when "00110011100010000" => rgb <= "000000";
					when "00110011100010001" => rgb <= "000000";
					when "00110011100010010" => rgb <= "000000";
					when "00110011100010011" => rgb <= "000000";
					when "00110011100010100" => rgb <= "000000";
					when "00110011100010101" => rgb <= "000000";
					when "00110011100010110" => rgb <= "000000";
					when "00110011100010111" => rgb <= "000000";
					when "00110011100011000" => rgb <= "000000";
					when "00110011100011001" => rgb <= "000000";
					when "00110011100011010" => rgb <= "000000";
					when "00110011100011011" => rgb <= "000000";
					when "00110011100011100" => rgb <= "000000";
					when "00110011100011101" => rgb <= "000000";
					when "00110011100011110" => rgb <= "000000";
					when "00110011100011111" => rgb <= "000000";
					when "00110011100100000" => rgb <= "000000";
					when "00110011100100001" => rgb <= "000000";
					when "00110011100100010" => rgb <= "000000";
					when "00110011100100011" => rgb <= "000000";
					when "00110011100100100" => rgb <= "000000";
					when "00110011100100101" => rgb <= "000000";
					when "00110011100100110" => rgb <= "000000";
					when "00110011100100111" => rgb <= "000000";
					when "00110011100101000" => rgb <= "000000";
					when "00110011100101001" => rgb <= "000000";
					when "00110011100101010" => rgb <= "000000";
					when "00110011100101011" => rgb <= "000000";
					when "00110011100101100" => rgb <= "000000";
					when "00110011100101101" => rgb <= "000000";
					when "00110011100101110" => rgb <= "000000";
					when "00110011100101111" => rgb <= "000000";
					when "00110011100110000" => rgb <= "000000";
					when "00110011100110001" => rgb <= "000000";
					when "00110011100110010" => rgb <= "000000";
					when "00110011100110011" => rgb <= "000000";
					when "00110011100110100" => rgb <= "000000";
					when "00110011100110101" => rgb <= "000000";
					when "00110011100110110" => rgb <= "000000";
					when "00110011100110111" => rgb <= "000000";
					when "00110011100111000" => rgb <= "000000";
					when "00110011100111001" => rgb <= "000000";
					when "00110011100111010" => rgb <= "000000";
					when "00110011100111011" => rgb <= "000000";
					when "00110011100111100" => rgb <= "000000";
					when "00110011100111101" => rgb <= "000000";
					when "00110011100111110" => rgb <= "000000";
					when "00110011100111111" => rgb <= "000000";
					when "00110100000000000" => rgb <= "000000";
					when "00110100000000001" => rgb <= "000000";
					when "00110100000000010" => rgb <= "000000";
					when "00110100000000011" => rgb <= "000000";
					when "00110100000000100" => rgb <= "000000";
					when "00110100000000101" => rgb <= "000000";
					when "00110100000000110" => rgb <= "000000";
					when "00110100000000111" => rgb <= "000000";
					when "00110100000001000" => rgb <= "000000";
					when "00110100000001001" => rgb <= "000000";
					when "00110100000001010" => rgb <= "000000";
					when "00110100000001011" => rgb <= "000000";
					when "00110100000001100" => rgb <= "000000";
					when "00110100000001101" => rgb <= "000000";
					when "00110100000001110" => rgb <= "000000";
					when "00110100000001111" => rgb <= "000000";
					when "00110100000010000" => rgb <= "000000";
					when "00110100000010001" => rgb <= "000000";
					when "00110100000010010" => rgb <= "000000";
					when "00110100000010011" => rgb <= "000000";
					when "00110100000010100" => rgb <= "000000";
					when "00110100000010101" => rgb <= "000000";
					when "00110100000010110" => rgb <= "000000";
					when "00110100000010111" => rgb <= "000000";
					when "00110100000011000" => rgb <= "000000";
					when "00110100000011001" => rgb <= "000000";
					when "00110100000011010" => rgb <= "000000";
					when "00110100000011011" => rgb <= "000000";
					when "00110100000011100" => rgb <= "000000";
					when "00110100000011101" => rgb <= "000000";
					when "00110100000011110" => rgb <= "000000";
					when "00110100000011111" => rgb <= "000000";
					when "00110100000100000" => rgb <= "000000";
					when "00110100000100001" => rgb <= "000000";
					when "00110100000100010" => rgb <= "000000";
					when "00110100000100011" => rgb <= "000000";
					when "00110100000100100" => rgb <= "000000";
					when "00110100000100101" => rgb <= "000000";
					when "00110100000100110" => rgb <= "000000";
					when "00110100000100111" => rgb <= "000000";
					when "00110100000101000" => rgb <= "000000";
					when "00110100000101001" => rgb <= "000000";
					when "00110100000101010" => rgb <= "000000";
					when "00110100000101011" => rgb <= "000000";
					when "00110100000101100" => rgb <= "000000";
					when "00110100000101101" => rgb <= "000000";
					when "00110100000101110" => rgb <= "000000";
					when "00110100000101111" => rgb <= "000000";
					when "00110100000110000" => rgb <= "000000";
					when "00110100000110001" => rgb <= "000000";
					when "00110100000110010" => rgb <= "000000";
					when "00110100000110011" => rgb <= "000000";
					when "00110100000110100" => rgb <= "000000";
					when "00110100000110101" => rgb <= "000000";
					when "00110100000110110" => rgb <= "000000";
					when "00110100000110111" => rgb <= "000000";
					when "00110100000111000" => rgb <= "000000";
					when "00110100000111001" => rgb <= "000000";
					when "00110100000111010" => rgb <= "000000";
					when "00110100000111011" => rgb <= "000000";
					when "00110100000111100" => rgb <= "000000";
					when "00110100000111101" => rgb <= "000000";
					when "00110100000111110" => rgb <= "000000";
					when "00110100000111111" => rgb <= "000000";
					when "00110100001000000" => rgb <= "000000";
					when "00110100001000001" => rgb <= "000000";
					when "00110100001000010" => rgb <= "000000";
					when "00110100001000011" => rgb <= "000000";
					when "00110100001000100" => rgb <= "000000";
					when "00110100001000101" => rgb <= "000000";
					when "00110100001000110" => rgb <= "000000";
					when "00110100001000111" => rgb <= "000000";
					when "00110100001001000" => rgb <= "000000";
					when "00110100001001001" => rgb <= "000000";
					when "00110100001001010" => rgb <= "000000";
					when "00110100001001011" => rgb <= "000000";
					when "00110100001001100" => rgb <= "000000";
					when "00110100001001101" => rgb <= "000000";
					when "00110100001001110" => rgb <= "000000";
					when "00110100001001111" => rgb <= "000000";
					when "00110100001010000" => rgb <= "000000";
					when "00110100001010001" => rgb <= "000000";
					when "00110100001010010" => rgb <= "000000";
					when "00110100001010011" => rgb <= "000000";
					when "00110100001010100" => rgb <= "000000";
					when "00110100001010101" => rgb <= "000000";
					when "00110100001010110" => rgb <= "000000";
					when "00110100001010111" => rgb <= "000000";
					when "00110100001011000" => rgb <= "000000";
					when "00110100001011001" => rgb <= "000000";
					when "00110100001011010" => rgb <= "000000";
					when "00110100001011011" => rgb <= "000000";
					when "00110100001011100" => rgb <= "000000";
					when "00110100001011101" => rgb <= "000000";
					when "00110100001011110" => rgb <= "000000";
					when "00110100001011111" => rgb <= "000000";
					when "00110100001100000" => rgb <= "000000";
					when "00110100001100001" => rgb <= "000000";
					when "00110100001100010" => rgb <= "000000";
					when "00110100001100011" => rgb <= "000000";
					when "00110100001100100" => rgb <= "000000";
					when "00110100001100101" => rgb <= "000000";
					when "00110100001100110" => rgb <= "010100";
					when "00110100001100111" => rgb <= "111000";
					when "00110100001101000" => rgb <= "101000";
					when "00110100001101001" => rgb <= "101000";
					when "00110100001101010" => rgb <= "101000";
					when "00110100001101011" => rgb <= "101000";
					when "00110100001101100" => rgb <= "101000";
					when "00110100001101101" => rgb <= "101000";
					when "00110100001101110" => rgb <= "101000";
					when "00110100001101111" => rgb <= "101000";
					when "00110100001110000" => rgb <= "101000";
					when "00110100001110001" => rgb <= "100100";
					when "00110100001110010" => rgb <= "000000";
					when "00110100001110011" => rgb <= "000000";
					when "00110100001110100" => rgb <= "000000";
					when "00110100001110101" => rgb <= "000000";
					when "00110100001110110" => rgb <= "000000";
					when "00110100001110111" => rgb <= "000000";
					when "00110100001111000" => rgb <= "000000";
					when "00110100001111001" => rgb <= "000000";
					when "00110100001111010" => rgb <= "000000";
					when "00110100001111011" => rgb <= "000000";
					when "00110100001111100" => rgb <= "000000";
					when "00110100001111101" => rgb <= "101000";
					when "00110100001111110" => rgb <= "101000";
					when "00110100001111111" => rgb <= "101000";
					when "00110100010000000" => rgb <= "101000";
					when "00110100010000001" => rgb <= "101000";
					when "00110100010000010" => rgb <= "101000";
					when "00110100010000011" => rgb <= "101000";
					when "00110100010000100" => rgb <= "101000";
					when "00110100010000101" => rgb <= "101000";
					when "00110100010000110" => rgb <= "101000";
					when "00110100010000111" => rgb <= "101000";
					when "00110100010001000" => rgb <= "101000";
					when "00110100010001001" => rgb <= "101000";
					when "00110100010001010" => rgb <= "101000";
					when "00110100010001011" => rgb <= "101000";
					when "00110100010001100" => rgb <= "101000";
					when "00110100010001101" => rgb <= "101000";
					when "00110100010001110" => rgb <= "101000";
					when "00110100010001111" => rgb <= "101000";
					when "00110100010010000" => rgb <= "101000";
					when "00110100010010001" => rgb <= "101000";
					when "00110100010010010" => rgb <= "101000";
					when "00110100010010011" => rgb <= "101000";
					when "00110100010010100" => rgb <= "101000";
					when "00110100010010101" => rgb <= "101000";
					when "00110100010010110" => rgb <= "101000";
					when "00110100010010111" => rgb <= "101000";
					when "00110100010011000" => rgb <= "101000";
					when "00110100010011001" => rgb <= "101000";
					when "00110100010011010" => rgb <= "101000";
					when "00110100010011011" => rgb <= "101000";
					when "00110100010011100" => rgb <= "101000";
					when "00110100010011101" => rgb <= "101000";
					when "00110100010011110" => rgb <= "101000";
					when "00110100010011111" => rgb <= "101000";
					when "00110100010100000" => rgb <= "101000";
					when "00110100010100001" => rgb <= "101000";
					when "00110100010100010" => rgb <= "101000";
					when "00110100010100011" => rgb <= "101000";
					when "00110100010100100" => rgb <= "101000";
					when "00110100010100101" => rgb <= "101000";
					when "00110100010100110" => rgb <= "101000";
					when "00110100010100111" => rgb <= "101000";
					when "00110100010101000" => rgb <= "101000";
					when "00110100010101001" => rgb <= "101000";
					when "00110100010101010" => rgb <= "101000";
					when "00110100010101011" => rgb <= "101000";
					when "00110100010101100" => rgb <= "101000";
					when "00110100010101101" => rgb <= "101000";
					when "00110100010101110" => rgb <= "101000";
					when "00110100010101111" => rgb <= "101000";
					when "00110100010110000" => rgb <= "101000";
					when "00110100010110001" => rgb <= "101000";
					when "00110100010110010" => rgb <= "101000";
					when "00110100010110011" => rgb <= "101000";
					when "00110100010110100" => rgb <= "101000";
					when "00110100010110101" => rgb <= "101000";
					when "00110100010110110" => rgb <= "101000";
					when "00110100010110111" => rgb <= "101000";
					when "00110100010111000" => rgb <= "101000";
					when "00110100010111001" => rgb <= "101000";
					when "00110100010111010" => rgb <= "101000";
					when "00110100010111011" => rgb <= "101000";
					when "00110100010111100" => rgb <= "101000";
					when "00110100010111101" => rgb <= "101000";
					when "00110100010111110" => rgb <= "101000";
					when "00110100010111111" => rgb <= "101000";
					when "00110100011000000" => rgb <= "100100";
					when "00110100011000001" => rgb <= "000000";
					when "00110100011000010" => rgb <= "000000";
					when "00110100011000011" => rgb <= "000000";
					when "00110100011000100" => rgb <= "000000";
					when "00110100011000101" => rgb <= "000000";
					when "00110100011000110" => rgb <= "000000";
					when "00110100011000111" => rgb <= "000000";
					when "00110100011001000" => rgb <= "000000";
					when "00110100011001001" => rgb <= "000000";
					when "00110100011001010" => rgb <= "000000";
					when "00110100011001011" => rgb <= "000000";
					when "00110100011001100" => rgb <= "100100";
					when "00110100011001101" => rgb <= "101000";
					when "00110100011001110" => rgb <= "101000";
					when "00110100011001111" => rgb <= "101000";
					when "00110100011010000" => rgb <= "101000";
					when "00110100011010001" => rgb <= "101000";
					when "00110100011010010" => rgb <= "101000";
					when "00110100011010011" => rgb <= "101000";
					when "00110100011010100" => rgb <= "101000";
					when "00110100011010101" => rgb <= "101000";
					when "00110100011010110" => rgb <= "101000";
					when "00110100011010111" => rgb <= "010100";
					when "00110100011011000" => rgb <= "000000";
					when "00110100011011001" => rgb <= "000000";
					when "00110100011011010" => rgb <= "000000";
					when "00110100011011011" => rgb <= "000000";
					when "00110100011011100" => rgb <= "000000";
					when "00110100011011101" => rgb <= "000000";
					when "00110100011011110" => rgb <= "000000";
					when "00110100011011111" => rgb <= "000000";
					when "00110100011100000" => rgb <= "000000";
					when "00110100011100001" => rgb <= "000000";
					when "00110100011100010" => rgb <= "000000";
					when "00110100011100011" => rgb <= "000000";
					when "00110100011100100" => rgb <= "000000";
					when "00110100011100101" => rgb <= "000000";
					when "00110100011100110" => rgb <= "000000";
					when "00110100011100111" => rgb <= "000000";
					when "00110100011101000" => rgb <= "000000";
					when "00110100011101001" => rgb <= "000000";
					when "00110100011101010" => rgb <= "000000";
					when "00110100011101011" => rgb <= "000000";
					when "00110100011101100" => rgb <= "000000";
					when "00110100011101101" => rgb <= "000000";
					when "00110100011101110" => rgb <= "000000";
					when "00110100011101111" => rgb <= "000000";
					when "00110100011110000" => rgb <= "000000";
					when "00110100011110001" => rgb <= "000000";
					when "00110100011110010" => rgb <= "000000";
					when "00110100011110011" => rgb <= "000000";
					when "00110100011110100" => rgb <= "000000";
					when "00110100011110101" => rgb <= "000000";
					when "00110100011110110" => rgb <= "000000";
					when "00110100011110111" => rgb <= "000000";
					when "00110100011111000" => rgb <= "000000";
					when "00110100011111001" => rgb <= "000000";
					when "00110100011111010" => rgb <= "000000";
					when "00110100011111011" => rgb <= "000000";
					when "00110100011111100" => rgb <= "000000";
					when "00110100011111101" => rgb <= "000000";
					when "00110100011111110" => rgb <= "000000";
					when "00110100011111111" => rgb <= "000000";
					when "00110100100000000" => rgb <= "000000";
					when "00110100100000001" => rgb <= "000000";
					when "00110100100000010" => rgb <= "000000";
					when "00110100100000011" => rgb <= "000000";
					when "00110100100000100" => rgb <= "000000";
					when "00110100100000101" => rgb <= "000000";
					when "00110100100000110" => rgb <= "000000";
					when "00110100100000111" => rgb <= "000000";
					when "00110100100001000" => rgb <= "000000";
					when "00110100100001001" => rgb <= "000000";
					when "00110100100001010" => rgb <= "000000";
					when "00110100100001011" => rgb <= "000000";
					when "00110100100001100" => rgb <= "000000";
					when "00110100100001101" => rgb <= "000000";
					when "00110100100001110" => rgb <= "000000";
					when "00110100100001111" => rgb <= "000000";
					when "00110100100010000" => rgb <= "000000";
					when "00110100100010001" => rgb <= "000000";
					when "00110100100010010" => rgb <= "000000";
					when "00110100100010011" => rgb <= "000000";
					when "00110100100010100" => rgb <= "000000";
					when "00110100100010101" => rgb <= "000000";
					when "00110100100010110" => rgb <= "000000";
					when "00110100100010111" => rgb <= "000000";
					when "00110100100011000" => rgb <= "000000";
					when "00110100100011001" => rgb <= "000000";
					when "00110100100011010" => rgb <= "000000";
					when "00110100100011011" => rgb <= "000000";
					when "00110100100011100" => rgb <= "000000";
					when "00110100100011101" => rgb <= "000000";
					when "00110100100011110" => rgb <= "000000";
					when "00110100100011111" => rgb <= "000000";
					when "00110100100100000" => rgb <= "000000";
					when "00110100100100001" => rgb <= "000000";
					when "00110100100100010" => rgb <= "000000";
					when "00110100100100011" => rgb <= "000000";
					when "00110100100100100" => rgb <= "000000";
					when "00110100100100101" => rgb <= "000000";
					when "00110100100100110" => rgb <= "000000";
					when "00110100100100111" => rgb <= "000000";
					when "00110100100101000" => rgb <= "000000";
					when "00110100100101001" => rgb <= "000000";
					when "00110100100101010" => rgb <= "000000";
					when "00110100100101011" => rgb <= "000000";
					when "00110100100101100" => rgb <= "000000";
					when "00110100100101101" => rgb <= "000000";
					when "00110100100101110" => rgb <= "000000";
					when "00110100100101111" => rgb <= "000000";
					when "00110100100110000" => rgb <= "000000";
					when "00110100100110001" => rgb <= "000000";
					when "00110100100110010" => rgb <= "000000";
					when "00110100100110011" => rgb <= "000000";
					when "00110100100110100" => rgb <= "000000";
					when "00110100100110101" => rgb <= "000000";
					when "00110100100110110" => rgb <= "000000";
					when "00110100100110111" => rgb <= "000000";
					when "00110100100111000" => rgb <= "000000";
					when "00110100100111001" => rgb <= "000000";
					when "00110100100111010" => rgb <= "000000";
					when "00110100100111011" => rgb <= "000000";
					when "00110100100111100" => rgb <= "000000";
					when "00110100100111101" => rgb <= "000000";
					when "00110100100111110" => rgb <= "000000";
					when "00110100100111111" => rgb <= "000000";
					when "00110101000000000" => rgb <= "000000";
					when "00110101000000001" => rgb <= "000000";
					when "00110101000000010" => rgb <= "000000";
					when "00110101000000011" => rgb <= "000000";
					when "00110101000000100" => rgb <= "000000";
					when "00110101000000101" => rgb <= "000000";
					when "00110101000000110" => rgb <= "000000";
					when "00110101000000111" => rgb <= "000000";
					when "00110101000001000" => rgb <= "000000";
					when "00110101000001001" => rgb <= "000000";
					when "00110101000001010" => rgb <= "000000";
					when "00110101000001011" => rgb <= "000000";
					when "00110101000001100" => rgb <= "000000";
					when "00110101000001101" => rgb <= "000000";
					when "00110101000001110" => rgb <= "000000";
					when "00110101000001111" => rgb <= "000000";
					when "00110101000010000" => rgb <= "000000";
					when "00110101000010001" => rgb <= "000000";
					when "00110101000010010" => rgb <= "000000";
					when "00110101000010011" => rgb <= "000000";
					when "00110101000010100" => rgb <= "000000";
					when "00110101000010101" => rgb <= "000000";
					when "00110101000010110" => rgb <= "000000";
					when "00110101000010111" => rgb <= "000000";
					when "00110101000011000" => rgb <= "000000";
					when "00110101000011001" => rgb <= "000000";
					when "00110101000011010" => rgb <= "000000";
					when "00110101000011011" => rgb <= "000000";
					when "00110101000011100" => rgb <= "000000";
					when "00110101000011101" => rgb <= "000000";
					when "00110101000011110" => rgb <= "000000";
					when "00110101000011111" => rgb <= "000000";
					when "00110101000100000" => rgb <= "000000";
					when "00110101000100001" => rgb <= "000000";
					when "00110101000100010" => rgb <= "000000";
					when "00110101000100011" => rgb <= "000000";
					when "00110101000100100" => rgb <= "000000";
					when "00110101000100101" => rgb <= "000000";
					when "00110101000100110" => rgb <= "000000";
					when "00110101000100111" => rgb <= "000000";
					when "00110101000101000" => rgb <= "000000";
					when "00110101000101001" => rgb <= "000000";
					when "00110101000101010" => rgb <= "000000";
					when "00110101000101011" => rgb <= "000000";
					when "00110101000101100" => rgb <= "000000";
					when "00110101000101101" => rgb <= "000000";
					when "00110101000101110" => rgb <= "000000";
					when "00110101000101111" => rgb <= "000000";
					when "00110101000110000" => rgb <= "000000";
					when "00110101000110001" => rgb <= "000000";
					when "00110101000110010" => rgb <= "000000";
					when "00110101000110011" => rgb <= "000000";
					when "00110101000110100" => rgb <= "000000";
					when "00110101000110101" => rgb <= "000000";
					when "00110101000110110" => rgb <= "000000";
					when "00110101000110111" => rgb <= "000000";
					when "00110101000111000" => rgb <= "000000";
					when "00110101000111001" => rgb <= "000000";
					when "00110101000111010" => rgb <= "000000";
					when "00110101000111011" => rgb <= "000000";
					when "00110101000111100" => rgb <= "000000";
					when "00110101000111101" => rgb <= "000000";
					when "00110101000111110" => rgb <= "000000";
					when "00110101000111111" => rgb <= "000000";
					when "00110101001000000" => rgb <= "000000";
					when "00110101001000001" => rgb <= "000000";
					when "00110101001000010" => rgb <= "000000";
					when "00110101001000011" => rgb <= "000000";
					when "00110101001000100" => rgb <= "000000";
					when "00110101001000101" => rgb <= "000000";
					when "00110101001000110" => rgb <= "000000";
					when "00110101001000111" => rgb <= "000000";
					when "00110101001001000" => rgb <= "000000";
					when "00110101001001001" => rgb <= "000000";
					when "00110101001001010" => rgb <= "000000";
					when "00110101001001011" => rgb <= "000000";
					when "00110101001001100" => rgb <= "000000";
					when "00110101001001101" => rgb <= "000000";
					when "00110101001001110" => rgb <= "000000";
					when "00110101001001111" => rgb <= "000000";
					when "00110101001010000" => rgb <= "000000";
					when "00110101001010001" => rgb <= "000000";
					when "00110101001010010" => rgb <= "000000";
					when "00110101001010011" => rgb <= "000000";
					when "00110101001010100" => rgb <= "000000";
					when "00110101001010101" => rgb <= "000000";
					when "00110101001010110" => rgb <= "000000";
					when "00110101001010111" => rgb <= "000000";
					when "00110101001011000" => rgb <= "000000";
					when "00110101001011001" => rgb <= "000000";
					when "00110101001011010" => rgb <= "000000";
					when "00110101001011011" => rgb <= "000000";
					when "00110101001011100" => rgb <= "000000";
					when "00110101001011101" => rgb <= "000000";
					when "00110101001011110" => rgb <= "000000";
					when "00110101001011111" => rgb <= "000000";
					when "00110101001100000" => rgb <= "000000";
					when "00110101001100001" => rgb <= "000000";
					when "00110101001100010" => rgb <= "000000";
					when "00110101001100011" => rgb <= "000000";
					when "00110101001100100" => rgb <= "000000";
					when "00110101001100101" => rgb <= "000000";
					when "00110101001100110" => rgb <= "010100";
					when "00110101001100111" => rgb <= "111000";
					when "00110101001101000" => rgb <= "101000";
					when "00110101001101001" => rgb <= "101000";
					when "00110101001101010" => rgb <= "101000";
					when "00110101001101011" => rgb <= "101000";
					when "00110101001101100" => rgb <= "101000";
					when "00110101001101101" => rgb <= "101000";
					when "00110101001101110" => rgb <= "101000";
					when "00110101001101111" => rgb <= "101000";
					when "00110101001110000" => rgb <= "111000";
					when "00110101001110001" => rgb <= "100100";
					when "00110101001110010" => rgb <= "000000";
					when "00110101001110011" => rgb <= "000000";
					when "00110101001110100" => rgb <= "000000";
					when "00110101001110101" => rgb <= "000000";
					when "00110101001110110" => rgb <= "000000";
					when "00110101001110111" => rgb <= "000000";
					when "00110101001111000" => rgb <= "000000";
					when "00110101001111001" => rgb <= "000000";
					when "00110101001111010" => rgb <= "000000";
					when "00110101001111011" => rgb <= "000000";
					when "00110101001111100" => rgb <= "000000";
					when "00110101001111101" => rgb <= "101000";
					when "00110101001111110" => rgb <= "101000";
					when "00110101001111111" => rgb <= "101000";
					when "00110101010000000" => rgb <= "101000";
					when "00110101010000001" => rgb <= "101000";
					when "00110101010000010" => rgb <= "101000";
					when "00110101010000011" => rgb <= "101000";
					when "00110101010000100" => rgb <= "101000";
					when "00110101010000101" => rgb <= "101000";
					when "00110101010000110" => rgb <= "101000";
					when "00110101010000111" => rgb <= "101000";
					when "00110101010001000" => rgb <= "101000";
					when "00110101010001001" => rgb <= "101000";
					when "00110101010001010" => rgb <= "101000";
					when "00110101010001011" => rgb <= "101000";
					when "00110101010001100" => rgb <= "101000";
					when "00110101010001101" => rgb <= "101000";
					when "00110101010001110" => rgb <= "101000";
					when "00110101010001111" => rgb <= "101000";
					when "00110101010010000" => rgb <= "101000";
					when "00110101010010001" => rgb <= "101000";
					when "00110101010010010" => rgb <= "101000";
					when "00110101010010011" => rgb <= "101000";
					when "00110101010010100" => rgb <= "101000";
					when "00110101010010101" => rgb <= "101000";
					when "00110101010010110" => rgb <= "101000";
					when "00110101010010111" => rgb <= "101000";
					when "00110101010011000" => rgb <= "101000";
					when "00110101010011001" => rgb <= "101000";
					when "00110101010011010" => rgb <= "101000";
					when "00110101010011011" => rgb <= "101000";
					when "00110101010011100" => rgb <= "101000";
					when "00110101010011101" => rgb <= "101000";
					when "00110101010011110" => rgb <= "101000";
					when "00110101010011111" => rgb <= "101000";
					when "00110101010100000" => rgb <= "101000";
					when "00110101010100001" => rgb <= "101000";
					when "00110101010100010" => rgb <= "101000";
					when "00110101010100011" => rgb <= "101000";
					when "00110101010100100" => rgb <= "101000";
					when "00110101010100101" => rgb <= "101000";
					when "00110101010100110" => rgb <= "101000";
					when "00110101010100111" => rgb <= "101000";
					when "00110101010101000" => rgb <= "101000";
					when "00110101010101001" => rgb <= "101000";
					when "00110101010101010" => rgb <= "101000";
					when "00110101010101011" => rgb <= "101000";
					when "00110101010101100" => rgb <= "101000";
					when "00110101010101101" => rgb <= "101000";
					when "00110101010101110" => rgb <= "101000";
					when "00110101010101111" => rgb <= "101000";
					when "00110101010110000" => rgb <= "101000";
					when "00110101010110001" => rgb <= "101000";
					when "00110101010110010" => rgb <= "101000";
					when "00110101010110011" => rgb <= "101000";
					when "00110101010110100" => rgb <= "101000";
					when "00110101010110101" => rgb <= "101000";
					when "00110101010110110" => rgb <= "101000";
					when "00110101010110111" => rgb <= "101000";
					when "00110101010111000" => rgb <= "101000";
					when "00110101010111001" => rgb <= "101000";
					when "00110101010111010" => rgb <= "101000";
					when "00110101010111011" => rgb <= "101000";
					when "00110101010111100" => rgb <= "101000";
					when "00110101010111101" => rgb <= "101000";
					when "00110101010111110" => rgb <= "101000";
					when "00110101010111111" => rgb <= "101000";
					when "00110101011000000" => rgb <= "101000";
					when "00110101011000001" => rgb <= "000000";
					when "00110101011000010" => rgb <= "000000";
					when "00110101011000011" => rgb <= "000000";
					when "00110101011000100" => rgb <= "000000";
					when "00110101011000101" => rgb <= "000000";
					when "00110101011000110" => rgb <= "000000";
					when "00110101011000111" => rgb <= "000000";
					when "00110101011001000" => rgb <= "000000";
					when "00110101011001001" => rgb <= "000000";
					when "00110101011001010" => rgb <= "000000";
					when "00110101011001011" => rgb <= "000000";
					when "00110101011001100" => rgb <= "100100";
					when "00110101011001101" => rgb <= "101000";
					when "00110101011001110" => rgb <= "101000";
					when "00110101011001111" => rgb <= "101000";
					when "00110101011010000" => rgb <= "101000";
					when "00110101011010001" => rgb <= "101000";
					when "00110101011010010" => rgb <= "101000";
					when "00110101011010011" => rgb <= "101000";
					when "00110101011010100" => rgb <= "101000";
					when "00110101011010101" => rgb <= "101000";
					when "00110101011010110" => rgb <= "101000";
					when "00110101011010111" => rgb <= "010100";
					when "00110101011011000" => rgb <= "000000";
					when "00110101011011001" => rgb <= "000000";
					when "00110101011011010" => rgb <= "000000";
					when "00110101011011011" => rgb <= "000000";
					when "00110101011011100" => rgb <= "000000";
					when "00110101011011101" => rgb <= "000000";
					when "00110101011011110" => rgb <= "000000";
					when "00110101011011111" => rgb <= "000000";
					when "00110101011100000" => rgb <= "000000";
					when "00110101011100001" => rgb <= "000000";
					when "00110101011100010" => rgb <= "000000";
					when "00110101011100011" => rgb <= "000000";
					when "00110101011100100" => rgb <= "000000";
					when "00110101011100101" => rgb <= "000000";
					when "00110101011100110" => rgb <= "000000";
					when "00110101011100111" => rgb <= "000000";
					when "00110101011101000" => rgb <= "000000";
					when "00110101011101001" => rgb <= "000000";
					when "00110101011101010" => rgb <= "000000";
					when "00110101011101011" => rgb <= "000000";
					when "00110101011101100" => rgb <= "000000";
					when "00110101011101101" => rgb <= "000000";
					when "00110101011101110" => rgb <= "000000";
					when "00110101011101111" => rgb <= "000000";
					when "00110101011110000" => rgb <= "000000";
					when "00110101011110001" => rgb <= "000000";
					when "00110101011110010" => rgb <= "000000";
					when "00110101011110011" => rgb <= "000000";
					when "00110101011110100" => rgb <= "000000";
					when "00110101011110101" => rgb <= "000000";
					when "00110101011110110" => rgb <= "000000";
					when "00110101011110111" => rgb <= "000000";
					when "00110101011111000" => rgb <= "000000";
					when "00110101011111001" => rgb <= "000000";
					when "00110101011111010" => rgb <= "000000";
					when "00110101011111011" => rgb <= "000000";
					when "00110101011111100" => rgb <= "000000";
					when "00110101011111101" => rgb <= "000000";
					when "00110101011111110" => rgb <= "000000";
					when "00110101011111111" => rgb <= "000000";
					when "00110101100000000" => rgb <= "000000";
					when "00110101100000001" => rgb <= "000000";
					when "00110101100000010" => rgb <= "000000";
					when "00110101100000011" => rgb <= "000000";
					when "00110101100000100" => rgb <= "000000";
					when "00110101100000101" => rgb <= "000000";
					when "00110101100000110" => rgb <= "000000";
					when "00110101100000111" => rgb <= "000000";
					when "00110101100001000" => rgb <= "000000";
					when "00110101100001001" => rgb <= "000000";
					when "00110101100001010" => rgb <= "000000";
					when "00110101100001011" => rgb <= "000000";
					when "00110101100001100" => rgb <= "000000";
					when "00110101100001101" => rgb <= "000000";
					when "00110101100001110" => rgb <= "000000";
					when "00110101100001111" => rgb <= "000000";
					when "00110101100010000" => rgb <= "000000";
					when "00110101100010001" => rgb <= "000000";
					when "00110101100010010" => rgb <= "000000";
					when "00110101100010011" => rgb <= "000000";
					when "00110101100010100" => rgb <= "000000";
					when "00110101100010101" => rgb <= "000000";
					when "00110101100010110" => rgb <= "000000";
					when "00110101100010111" => rgb <= "000000";
					when "00110101100011000" => rgb <= "000000";
					when "00110101100011001" => rgb <= "000000";
					when "00110101100011010" => rgb <= "000000";
					when "00110101100011011" => rgb <= "000000";
					when "00110101100011100" => rgb <= "000000";
					when "00110101100011101" => rgb <= "000000";
					when "00110101100011110" => rgb <= "000000";
					when "00110101100011111" => rgb <= "000000";
					when "00110101100100000" => rgb <= "000000";
					when "00110101100100001" => rgb <= "000000";
					when "00110101100100010" => rgb <= "000000";
					when "00110101100100011" => rgb <= "000000";
					when "00110101100100100" => rgb <= "000000";
					when "00110101100100101" => rgb <= "000000";
					when "00110101100100110" => rgb <= "000000";
					when "00110101100100111" => rgb <= "000000";
					when "00110101100101000" => rgb <= "000000";
					when "00110101100101001" => rgb <= "000000";
					when "00110101100101010" => rgb <= "000000";
					when "00110101100101011" => rgb <= "000000";
					when "00110101100101100" => rgb <= "000000";
					when "00110101100101101" => rgb <= "000000";
					when "00110101100101110" => rgb <= "000000";
					when "00110101100101111" => rgb <= "000000";
					when "00110101100110000" => rgb <= "000000";
					when "00110101100110001" => rgb <= "000000";
					when "00110101100110010" => rgb <= "000000";
					when "00110101100110011" => rgb <= "000000";
					when "00110101100110100" => rgb <= "000000";
					when "00110101100110101" => rgb <= "000000";
					when "00110101100110110" => rgb <= "000000";
					when "00110101100110111" => rgb <= "000000";
					when "00110101100111000" => rgb <= "000000";
					when "00110101100111001" => rgb <= "000000";
					when "00110101100111010" => rgb <= "000000";
					when "00110101100111011" => rgb <= "000000";
					when "00110101100111100" => rgb <= "000000";
					when "00110101100111101" => rgb <= "000000";
					when "00110101100111110" => rgb <= "000000";
					when "00110101100111111" => rgb <= "000000";
					when "00110110000000000" => rgb <= "000000";
					when "00110110000000001" => rgb <= "000000";
					when "00110110000000010" => rgb <= "000000";
					when "00110110000000011" => rgb <= "000000";
					when "00110110000000100" => rgb <= "000000";
					when "00110110000000101" => rgb <= "000000";
					when "00110110000000110" => rgb <= "000000";
					when "00110110000000111" => rgb <= "000000";
					when "00110110000001000" => rgb <= "000000";
					when "00110110000001001" => rgb <= "000000";
					when "00110110000001010" => rgb <= "000000";
					when "00110110000001011" => rgb <= "000000";
					when "00110110000001100" => rgb <= "000000";
					when "00110110000001101" => rgb <= "000000";
					when "00110110000001110" => rgb <= "000000";
					when "00110110000001111" => rgb <= "000000";
					when "00110110000010000" => rgb <= "000000";
					when "00110110000010001" => rgb <= "000000";
					when "00110110000010010" => rgb <= "000000";
					when "00110110000010011" => rgb <= "000000";
					when "00110110000010100" => rgb <= "000000";
					when "00110110000010101" => rgb <= "000000";
					when "00110110000010110" => rgb <= "000000";
					when "00110110000010111" => rgb <= "000000";
					when "00110110000011000" => rgb <= "000000";
					when "00110110000011001" => rgb <= "000000";
					when "00110110000011010" => rgb <= "000000";
					when "00110110000011011" => rgb <= "000000";
					when "00110110000011100" => rgb <= "000000";
					when "00110110000011101" => rgb <= "000000";
					when "00110110000011110" => rgb <= "000000";
					when "00110110000011111" => rgb <= "000000";
					when "00110110000100000" => rgb <= "000000";
					when "00110110000100001" => rgb <= "000000";
					when "00110110000100010" => rgb <= "000000";
					when "00110110000100011" => rgb <= "000000";
					when "00110110000100100" => rgb <= "000000";
					when "00110110000100101" => rgb <= "000000";
					when "00110110000100110" => rgb <= "000000";
					when "00110110000100111" => rgb <= "000000";
					when "00110110000101000" => rgb <= "000000";
					when "00110110000101001" => rgb <= "000000";
					when "00110110000101010" => rgb <= "000000";
					when "00110110000101011" => rgb <= "000000";
					when "00110110000101100" => rgb <= "000000";
					when "00110110000101101" => rgb <= "000000";
					when "00110110000101110" => rgb <= "000000";
					when "00110110000101111" => rgb <= "000000";
					when "00110110000110000" => rgb <= "000000";
					when "00110110000110001" => rgb <= "000000";
					when "00110110000110010" => rgb <= "000000";
					when "00110110000110011" => rgb <= "000000";
					when "00110110000110100" => rgb <= "000000";
					when "00110110000110101" => rgb <= "000000";
					when "00110110000110110" => rgb <= "000000";
					when "00110110000110111" => rgb <= "000000";
					when "00110110000111000" => rgb <= "000000";
					when "00110110000111001" => rgb <= "000000";
					when "00110110000111010" => rgb <= "000000";
					when "00110110000111011" => rgb <= "000000";
					when "00110110000111100" => rgb <= "000000";
					when "00110110000111101" => rgb <= "000000";
					when "00110110000111110" => rgb <= "000000";
					when "00110110000111111" => rgb <= "000000";
					when "00110110001000000" => rgb <= "000000";
					when "00110110001000001" => rgb <= "000000";
					when "00110110001000010" => rgb <= "000000";
					when "00110110001000011" => rgb <= "000000";
					when "00110110001000100" => rgb <= "000000";
					when "00110110001000101" => rgb <= "000000";
					when "00110110001000110" => rgb <= "000000";
					when "00110110001000111" => rgb <= "000000";
					when "00110110001001000" => rgb <= "000000";
					when "00110110001001001" => rgb <= "000000";
					when "00110110001001010" => rgb <= "000000";
					when "00110110001001011" => rgb <= "000000";
					when "00110110001001100" => rgb <= "000000";
					when "00110110001001101" => rgb <= "000000";
					when "00110110001001110" => rgb <= "000000";
					when "00110110001001111" => rgb <= "000000";
					when "00110110001010000" => rgb <= "000000";
					when "00110110001010001" => rgb <= "000000";
					when "00110110001010010" => rgb <= "000000";
					when "00110110001010011" => rgb <= "000000";
					when "00110110001010100" => rgb <= "000000";
					when "00110110001010101" => rgb <= "000000";
					when "00110110001010110" => rgb <= "000000";
					when "00110110001010111" => rgb <= "000000";
					when "00110110001011000" => rgb <= "000000";
					when "00110110001011001" => rgb <= "000000";
					when "00110110001011010" => rgb <= "000000";
					when "00110110001011011" => rgb <= "000000";
					when "00110110001011100" => rgb <= "000000";
					when "00110110001011101" => rgb <= "000000";
					when "00110110001011110" => rgb <= "000000";
					when "00110110001011111" => rgb <= "000000";
					when "00110110001100000" => rgb <= "000000";
					when "00110110001100001" => rgb <= "000000";
					when "00110110001100010" => rgb <= "000000";
					when "00110110001100011" => rgb <= "000000";
					when "00110110001100100" => rgb <= "000000";
					when "00110110001100101" => rgb <= "000000";
					when "00110110001100110" => rgb <= "010100";
					when "00110110001100111" => rgb <= "111000";
					when "00110110001101000" => rgb <= "101000";
					when "00110110001101001" => rgb <= "101000";
					when "00110110001101010" => rgb <= "101000";
					when "00110110001101011" => rgb <= "101000";
					when "00110110001101100" => rgb <= "101000";
					when "00110110001101101" => rgb <= "101000";
					when "00110110001101110" => rgb <= "101000";
					when "00110110001101111" => rgb <= "101000";
					when "00110110001110000" => rgb <= "111000";
					when "00110110001110001" => rgb <= "100100";
					when "00110110001110010" => rgb <= "000000";
					when "00110110001110011" => rgb <= "000000";
					when "00110110001110100" => rgb <= "000000";
					when "00110110001110101" => rgb <= "000000";
					when "00110110001110110" => rgb <= "000000";
					when "00110110001110111" => rgb <= "000000";
					when "00110110001111000" => rgb <= "000000";
					when "00110110001111001" => rgb <= "000000";
					when "00110110001111010" => rgb <= "000000";
					when "00110110001111011" => rgb <= "000000";
					when "00110110001111100" => rgb <= "000000";
					when "00110110001111101" => rgb <= "101000";
					when "00110110001111110" => rgb <= "101000";
					when "00110110001111111" => rgb <= "101000";
					when "00110110010000000" => rgb <= "101000";
					when "00110110010000001" => rgb <= "101000";
					when "00110110010000010" => rgb <= "101000";
					when "00110110010000011" => rgb <= "101000";
					when "00110110010000100" => rgb <= "101000";
					when "00110110010000101" => rgb <= "101000";
					when "00110110010000110" => rgb <= "101000";
					when "00110110010000111" => rgb <= "101000";
					when "00110110010001000" => rgb <= "101000";
					when "00110110010001001" => rgb <= "101000";
					when "00110110010001010" => rgb <= "101000";
					when "00110110010001011" => rgb <= "101000";
					when "00110110010001100" => rgb <= "101000";
					when "00110110010001101" => rgb <= "101000";
					when "00110110010001110" => rgb <= "101000";
					when "00110110010001111" => rgb <= "101000";
					when "00110110010010000" => rgb <= "101000";
					when "00110110010010001" => rgb <= "101000";
					when "00110110010010010" => rgb <= "101000";
					when "00110110010010011" => rgb <= "101000";
					when "00110110010010100" => rgb <= "101000";
					when "00110110010010101" => rgb <= "101000";
					when "00110110010010110" => rgb <= "101000";
					when "00110110010010111" => rgb <= "101000";
					when "00110110010011000" => rgb <= "101000";
					when "00110110010011001" => rgb <= "101000";
					when "00110110010011010" => rgb <= "101000";
					when "00110110010011011" => rgb <= "101000";
					when "00110110010011100" => rgb <= "101000";
					when "00110110010011101" => rgb <= "101000";
					when "00110110010011110" => rgb <= "101000";
					when "00110110010011111" => rgb <= "101000";
					when "00110110010100000" => rgb <= "101000";
					when "00110110010100001" => rgb <= "101000";
					when "00110110010100010" => rgb <= "101000";
					when "00110110010100011" => rgb <= "101000";
					when "00110110010100100" => rgb <= "101000";
					when "00110110010100101" => rgb <= "101000";
					when "00110110010100110" => rgb <= "101000";
					when "00110110010100111" => rgb <= "101000";
					when "00110110010101000" => rgb <= "101000";
					when "00110110010101001" => rgb <= "101000";
					when "00110110010101010" => rgb <= "101000";
					when "00110110010101011" => rgb <= "101000";
					when "00110110010101100" => rgb <= "101000";
					when "00110110010101101" => rgb <= "101000";
					when "00110110010101110" => rgb <= "101000";
					when "00110110010101111" => rgb <= "101000";
					when "00110110010110000" => rgb <= "101000";
					when "00110110010110001" => rgb <= "101000";
					when "00110110010110010" => rgb <= "101000";
					when "00110110010110011" => rgb <= "101000";
					when "00110110010110100" => rgb <= "101000";
					when "00110110010110101" => rgb <= "101000";
					when "00110110010110110" => rgb <= "101000";
					when "00110110010110111" => rgb <= "101000";
					when "00110110010111000" => rgb <= "101000";
					when "00110110010111001" => rgb <= "101000";
					when "00110110010111010" => rgb <= "101000";
					when "00110110010111011" => rgb <= "101000";
					when "00110110010111100" => rgb <= "101000";
					when "00110110010111101" => rgb <= "101000";
					when "00110110010111110" => rgb <= "101000";
					when "00110110010111111" => rgb <= "101000";
					when "00110110011000000" => rgb <= "100100";
					when "00110110011000001" => rgb <= "000000";
					when "00110110011000010" => rgb <= "000000";
					when "00110110011000011" => rgb <= "000000";
					when "00110110011000100" => rgb <= "000000";
					when "00110110011000101" => rgb <= "000000";
					when "00110110011000110" => rgb <= "000000";
					when "00110110011000111" => rgb <= "000000";
					when "00110110011001000" => rgb <= "000000";
					when "00110110011001001" => rgb <= "000000";
					when "00110110011001010" => rgb <= "000000";
					when "00110110011001011" => rgb <= "000000";
					when "00110110011001100" => rgb <= "100100";
					when "00110110011001101" => rgb <= "101000";
					when "00110110011001110" => rgb <= "101000";
					when "00110110011001111" => rgb <= "101000";
					when "00110110011010000" => rgb <= "101000";
					when "00110110011010001" => rgb <= "101000";
					when "00110110011010010" => rgb <= "101000";
					when "00110110011010011" => rgb <= "101000";
					when "00110110011010100" => rgb <= "101000";
					when "00110110011010101" => rgb <= "101000";
					when "00110110011010110" => rgb <= "101000";
					when "00110110011010111" => rgb <= "010100";
					when "00110110011011000" => rgb <= "000000";
					when "00110110011011001" => rgb <= "000000";
					when "00110110011011010" => rgb <= "000000";
					when "00110110011011011" => rgb <= "000000";
					when "00110110011011100" => rgb <= "000000";
					when "00110110011011101" => rgb <= "000000";
					when "00110110011011110" => rgb <= "000000";
					when "00110110011011111" => rgb <= "000000";
					when "00110110011100000" => rgb <= "000000";
					when "00110110011100001" => rgb <= "000000";
					when "00110110011100010" => rgb <= "000000";
					when "00110110011100011" => rgb <= "000000";
					when "00110110011100100" => rgb <= "000000";
					when "00110110011100101" => rgb <= "000000";
					when "00110110011100110" => rgb <= "000000";
					when "00110110011100111" => rgb <= "000000";
					when "00110110011101000" => rgb <= "000000";
					when "00110110011101001" => rgb <= "000000";
					when "00110110011101010" => rgb <= "000000";
					when "00110110011101011" => rgb <= "000000";
					when "00110110011101100" => rgb <= "000000";
					when "00110110011101101" => rgb <= "000000";
					when "00110110011101110" => rgb <= "000000";
					when "00110110011101111" => rgb <= "000000";
					when "00110110011110000" => rgb <= "000000";
					when "00110110011110001" => rgb <= "000000";
					when "00110110011110010" => rgb <= "000000";
					when "00110110011110011" => rgb <= "000000";
					when "00110110011110100" => rgb <= "000000";
					when "00110110011110101" => rgb <= "000000";
					when "00110110011110110" => rgb <= "000000";
					when "00110110011110111" => rgb <= "000000";
					when "00110110011111000" => rgb <= "000000";
					when "00110110011111001" => rgb <= "000000";
					when "00110110011111010" => rgb <= "000000";
					when "00110110011111011" => rgb <= "000000";
					when "00110110011111100" => rgb <= "000000";
					when "00110110011111101" => rgb <= "000000";
					when "00110110011111110" => rgb <= "000000";
					when "00110110011111111" => rgb <= "000000";
					when "00110110100000000" => rgb <= "000000";
					when "00110110100000001" => rgb <= "000000";
					when "00110110100000010" => rgb <= "000000";
					when "00110110100000011" => rgb <= "000000";
					when "00110110100000100" => rgb <= "000000";
					when "00110110100000101" => rgb <= "000000";
					when "00110110100000110" => rgb <= "000000";
					when "00110110100000111" => rgb <= "000000";
					when "00110110100001000" => rgb <= "000000";
					when "00110110100001001" => rgb <= "000000";
					when "00110110100001010" => rgb <= "000000";
					when "00110110100001011" => rgb <= "000000";
					when "00110110100001100" => rgb <= "000000";
					when "00110110100001101" => rgb <= "000000";
					when "00110110100001110" => rgb <= "000000";
					when "00110110100001111" => rgb <= "000000";
					when "00110110100010000" => rgb <= "000000";
					when "00110110100010001" => rgb <= "000000";
					when "00110110100010010" => rgb <= "000000";
					when "00110110100010011" => rgb <= "000000";
					when "00110110100010100" => rgb <= "000000";
					when "00110110100010101" => rgb <= "000000";
					when "00110110100010110" => rgb <= "000000";
					when "00110110100010111" => rgb <= "000000";
					when "00110110100011000" => rgb <= "000000";
					when "00110110100011001" => rgb <= "000000";
					when "00110110100011010" => rgb <= "000000";
					when "00110110100011011" => rgb <= "000000";
					when "00110110100011100" => rgb <= "000000";
					when "00110110100011101" => rgb <= "000000";
					when "00110110100011110" => rgb <= "000000";
					when "00110110100011111" => rgb <= "000000";
					when "00110110100100000" => rgb <= "000000";
					when "00110110100100001" => rgb <= "000000";
					when "00110110100100010" => rgb <= "000000";
					when "00110110100100011" => rgb <= "000000";
					when "00110110100100100" => rgb <= "000000";
					when "00110110100100101" => rgb <= "000000";
					when "00110110100100110" => rgb <= "000000";
					when "00110110100100111" => rgb <= "000000";
					when "00110110100101000" => rgb <= "000000";
					when "00110110100101001" => rgb <= "000000";
					when "00110110100101010" => rgb <= "000000";
					when "00110110100101011" => rgb <= "000000";
					when "00110110100101100" => rgb <= "000000";
					when "00110110100101101" => rgb <= "000000";
					when "00110110100101110" => rgb <= "000000";
					when "00110110100101111" => rgb <= "000000";
					when "00110110100110000" => rgb <= "000000";
					when "00110110100110001" => rgb <= "000000";
					when "00110110100110010" => rgb <= "000000";
					when "00110110100110011" => rgb <= "000000";
					when "00110110100110100" => rgb <= "000000";
					when "00110110100110101" => rgb <= "000000";
					when "00110110100110110" => rgb <= "000000";
					when "00110110100110111" => rgb <= "000000";
					when "00110110100111000" => rgb <= "000000";
					when "00110110100111001" => rgb <= "000000";
					when "00110110100111010" => rgb <= "000000";
					when "00110110100111011" => rgb <= "000000";
					when "00110110100111100" => rgb <= "000000";
					when "00110110100111101" => rgb <= "000000";
					when "00110110100111110" => rgb <= "000000";
					when "00110110100111111" => rgb <= "000000";
					when "00110111000000000" => rgb <= "000000";
					when "00110111000000001" => rgb <= "000000";
					when "00110111000000010" => rgb <= "000000";
					when "00110111000000011" => rgb <= "000000";
					when "00110111000000100" => rgb <= "000000";
					when "00110111000000101" => rgb <= "000000";
					when "00110111000000110" => rgb <= "000000";
					when "00110111000000111" => rgb <= "000000";
					when "00110111000001000" => rgb <= "000000";
					when "00110111000001001" => rgb <= "000000";
					when "00110111000001010" => rgb <= "000000";
					when "00110111000001011" => rgb <= "000000";
					when "00110111000001100" => rgb <= "000000";
					when "00110111000001101" => rgb <= "000000";
					when "00110111000001110" => rgb <= "000000";
					when "00110111000001111" => rgb <= "000000";
					when "00110111000010000" => rgb <= "000000";
					when "00110111000010001" => rgb <= "000000";
					when "00110111000010010" => rgb <= "000000";
					when "00110111000010011" => rgb <= "000000";
					when "00110111000010100" => rgb <= "000000";
					when "00110111000010101" => rgb <= "000000";
					when "00110111000010110" => rgb <= "000000";
					when "00110111000010111" => rgb <= "000000";
					when "00110111000011000" => rgb <= "000000";
					when "00110111000011001" => rgb <= "000000";
					when "00110111000011010" => rgb <= "000000";
					when "00110111000011011" => rgb <= "000000";
					when "00110111000011100" => rgb <= "000000";
					when "00110111000011101" => rgb <= "000000";
					when "00110111000011110" => rgb <= "000000";
					when "00110111000011111" => rgb <= "000000";
					when "00110111000100000" => rgb <= "000000";
					when "00110111000100001" => rgb <= "000000";
					when "00110111000100010" => rgb <= "000000";
					when "00110111000100011" => rgb <= "000000";
					when "00110111000100100" => rgb <= "000000";
					when "00110111000100101" => rgb <= "000000";
					when "00110111000100110" => rgb <= "000000";
					when "00110111000100111" => rgb <= "000000";
					when "00110111000101000" => rgb <= "000000";
					when "00110111000101001" => rgb <= "000000";
					when "00110111000101010" => rgb <= "000000";
					when "00110111000101011" => rgb <= "000000";
					when "00110111000101100" => rgb <= "000000";
					when "00110111000101101" => rgb <= "000000";
					when "00110111000101110" => rgb <= "000000";
					when "00110111000101111" => rgb <= "000000";
					when "00110111000110000" => rgb <= "000000";
					when "00110111000110001" => rgb <= "000000";
					when "00110111000110010" => rgb <= "000000";
					when "00110111000110011" => rgb <= "000000";
					when "00110111000110100" => rgb <= "000000";
					when "00110111000110101" => rgb <= "000000";
					when "00110111000110110" => rgb <= "000000";
					when "00110111000110111" => rgb <= "000000";
					when "00110111000111000" => rgb <= "000000";
					when "00110111000111001" => rgb <= "000000";
					when "00110111000111010" => rgb <= "000000";
					when "00110111000111011" => rgb <= "000000";
					when "00110111000111100" => rgb <= "000000";
					when "00110111000111101" => rgb <= "000000";
					when "00110111000111110" => rgb <= "000000";
					when "00110111000111111" => rgb <= "000000";
					when "00110111001000000" => rgb <= "000000";
					when "00110111001000001" => rgb <= "000000";
					when "00110111001000010" => rgb <= "000000";
					when "00110111001000011" => rgb <= "000000";
					when "00110111001000100" => rgb <= "000000";
					when "00110111001000101" => rgb <= "000000";
					when "00110111001000110" => rgb <= "000000";
					when "00110111001000111" => rgb <= "000000";
					when "00110111001001000" => rgb <= "000000";
					when "00110111001001001" => rgb <= "000000";
					when "00110111001001010" => rgb <= "000000";
					when "00110111001001011" => rgb <= "000000";
					when "00110111001001100" => rgb <= "000000";
					when "00110111001001101" => rgb <= "000000";
					when "00110111001001110" => rgb <= "000000";
					when "00110111001001111" => rgb <= "000000";
					when "00110111001010000" => rgb <= "000000";
					when "00110111001010001" => rgb <= "000000";
					when "00110111001010010" => rgb <= "000000";
					when "00110111001010011" => rgb <= "000000";
					when "00110111001010100" => rgb <= "000000";
					when "00110111001010101" => rgb <= "000000";
					when "00110111001010110" => rgb <= "000000";
					when "00110111001010111" => rgb <= "000000";
					when "00110111001011000" => rgb <= "000000";
					when "00110111001011001" => rgb <= "000000";
					when "00110111001011010" => rgb <= "000000";
					when "00110111001011011" => rgb <= "000000";
					when "00110111001011100" => rgb <= "000000";
					when "00110111001011101" => rgb <= "000000";
					when "00110111001011110" => rgb <= "000000";
					when "00110111001011111" => rgb <= "000000";
					when "00110111001100000" => rgb <= "000000";
					when "00110111001100001" => rgb <= "000000";
					when "00110111001100010" => rgb <= "000000";
					when "00110111001100011" => rgb <= "000000";
					when "00110111001100100" => rgb <= "000000";
					when "00110111001100101" => rgb <= "000000";
					when "00110111001100110" => rgb <= "010100";
					when "00110111001100111" => rgb <= "111000";
					when "00110111001101000" => rgb <= "101000";
					when "00110111001101001" => rgb <= "101000";
					when "00110111001101010" => rgb <= "101000";
					when "00110111001101011" => rgb <= "101000";
					when "00110111001101100" => rgb <= "101000";
					when "00110111001101101" => rgb <= "101000";
					when "00110111001101110" => rgb <= "101000";
					when "00110111001101111" => rgb <= "101000";
					when "00110111001110000" => rgb <= "101000";
					when "00110111001110001" => rgb <= "100100";
					when "00110111001110010" => rgb <= "000000";
					when "00110111001110011" => rgb <= "000000";
					when "00110111001110100" => rgb <= "000000";
					when "00110111001110101" => rgb <= "000000";
					when "00110111001110110" => rgb <= "000000";
					when "00110111001110111" => rgb <= "000000";
					when "00110111001111000" => rgb <= "000000";
					when "00110111001111001" => rgb <= "000000";
					when "00110111001111010" => rgb <= "000000";
					when "00110111001111011" => rgb <= "000000";
					when "00110111001111100" => rgb <= "000000";
					when "00110111001111101" => rgb <= "101000";
					when "00110111001111110" => rgb <= "101000";
					when "00110111001111111" => rgb <= "101000";
					when "00110111010000000" => rgb <= "101000";
					when "00110111010000001" => rgb <= "101000";
					when "00110111010000010" => rgb <= "101000";
					when "00110111010000011" => rgb <= "101000";
					when "00110111010000100" => rgb <= "101000";
					when "00110111010000101" => rgb <= "101000";
					when "00110111010000110" => rgb <= "101000";
					when "00110111010000111" => rgb <= "101000";
					when "00110111010001000" => rgb <= "101000";
					when "00110111010001001" => rgb <= "101000";
					when "00110111010001010" => rgb <= "101000";
					when "00110111010001011" => rgb <= "101000";
					when "00110111010001100" => rgb <= "101000";
					when "00110111010001101" => rgb <= "101000";
					when "00110111010001110" => rgb <= "101000";
					when "00110111010001111" => rgb <= "101000";
					when "00110111010010000" => rgb <= "101000";
					when "00110111010010001" => rgb <= "101000";
					when "00110111010010010" => rgb <= "101000";
					when "00110111010010011" => rgb <= "101000";
					when "00110111010010100" => rgb <= "101000";
					when "00110111010010101" => rgb <= "101000";
					when "00110111010010110" => rgb <= "101000";
					when "00110111010010111" => rgb <= "101000";
					when "00110111010011000" => rgb <= "101000";
					when "00110111010011001" => rgb <= "101000";
					when "00110111010011010" => rgb <= "101000";
					when "00110111010011011" => rgb <= "101000";
					when "00110111010011100" => rgb <= "101000";
					when "00110111010011101" => rgb <= "101000";
					when "00110111010011110" => rgb <= "101000";
					when "00110111010011111" => rgb <= "101000";
					when "00110111010100000" => rgb <= "101000";
					when "00110111010100001" => rgb <= "101000";
					when "00110111010100010" => rgb <= "101000";
					when "00110111010100011" => rgb <= "101000";
					when "00110111010100100" => rgb <= "101000";
					when "00110111010100101" => rgb <= "101000";
					when "00110111010100110" => rgb <= "101000";
					when "00110111010100111" => rgb <= "101000";
					when "00110111010101000" => rgb <= "101000";
					when "00110111010101001" => rgb <= "101000";
					when "00110111010101010" => rgb <= "101000";
					when "00110111010101011" => rgb <= "101000";
					when "00110111010101100" => rgb <= "101000";
					when "00110111010101101" => rgb <= "101000";
					when "00110111010101110" => rgb <= "101000";
					when "00110111010101111" => rgb <= "101000";
					when "00110111010110000" => rgb <= "101000";
					when "00110111010110001" => rgb <= "101000";
					when "00110111010110010" => rgb <= "101000";
					when "00110111010110011" => rgb <= "101000";
					when "00110111010110100" => rgb <= "101000";
					when "00110111010110101" => rgb <= "101000";
					when "00110111010110110" => rgb <= "101000";
					when "00110111010110111" => rgb <= "101000";
					when "00110111010111000" => rgb <= "101000";
					when "00110111010111001" => rgb <= "101000";
					when "00110111010111010" => rgb <= "101000";
					when "00110111010111011" => rgb <= "101000";
					when "00110111010111100" => rgb <= "101000";
					when "00110111010111101" => rgb <= "101000";
					when "00110111010111110" => rgb <= "101000";
					when "00110111010111111" => rgb <= "101000";
					when "00110111011000000" => rgb <= "100100";
					when "00110111011000001" => rgb <= "000000";
					when "00110111011000010" => rgb <= "000000";
					when "00110111011000011" => rgb <= "000000";
					when "00110111011000100" => rgb <= "000000";
					when "00110111011000101" => rgb <= "000000";
					when "00110111011000110" => rgb <= "000000";
					when "00110111011000111" => rgb <= "000000";
					when "00110111011001000" => rgb <= "000000";
					when "00110111011001001" => rgb <= "000000";
					when "00110111011001010" => rgb <= "000000";
					when "00110111011001011" => rgb <= "000000";
					when "00110111011001100" => rgb <= "010100";
					when "00110111011001101" => rgb <= "101000";
					when "00110111011001110" => rgb <= "101000";
					when "00110111011001111" => rgb <= "101000";
					when "00110111011010000" => rgb <= "101000";
					when "00110111011010001" => rgb <= "101000";
					when "00110111011010010" => rgb <= "101000";
					when "00110111011010011" => rgb <= "101000";
					when "00110111011010100" => rgb <= "101000";
					when "00110111011010101" => rgb <= "101000";
					when "00110111011010110" => rgb <= "101000";
					when "00110111011010111" => rgb <= "010100";
					when "00110111011011000" => rgb <= "000000";
					when "00110111011011001" => rgb <= "000000";
					when "00110111011011010" => rgb <= "000000";
					when "00110111011011011" => rgb <= "000000";
					when "00110111011011100" => rgb <= "000000";
					when "00110111011011101" => rgb <= "000000";
					when "00110111011011110" => rgb <= "000000";
					when "00110111011011111" => rgb <= "000000";
					when "00110111011100000" => rgb <= "000000";
					when "00110111011100001" => rgb <= "000000";
					when "00110111011100010" => rgb <= "000000";
					when "00110111011100011" => rgb <= "000000";
					when "00110111011100100" => rgb <= "000000";
					when "00110111011100101" => rgb <= "000000";
					when "00110111011100110" => rgb <= "000000";
					when "00110111011100111" => rgb <= "000000";
					when "00110111011101000" => rgb <= "000000";
					when "00110111011101001" => rgb <= "000000";
					when "00110111011101010" => rgb <= "000000";
					when "00110111011101011" => rgb <= "000000";
					when "00110111011101100" => rgb <= "000000";
					when "00110111011101101" => rgb <= "000000";
					when "00110111011101110" => rgb <= "000000";
					when "00110111011101111" => rgb <= "000000";
					when "00110111011110000" => rgb <= "000000";
					when "00110111011110001" => rgb <= "000000";
					when "00110111011110010" => rgb <= "000000";
					when "00110111011110011" => rgb <= "000000";
					when "00110111011110100" => rgb <= "000000";
					when "00110111011110101" => rgb <= "000000";
					when "00110111011110110" => rgb <= "000000";
					when "00110111011110111" => rgb <= "000000";
					when "00110111011111000" => rgb <= "000000";
					when "00110111011111001" => rgb <= "000000";
					when "00110111011111010" => rgb <= "000000";
					when "00110111011111011" => rgb <= "000000";
					when "00110111011111100" => rgb <= "000000";
					when "00110111011111101" => rgb <= "000000";
					when "00110111011111110" => rgb <= "000000";
					when "00110111011111111" => rgb <= "000000";
					when "00110111100000000" => rgb <= "000000";
					when "00110111100000001" => rgb <= "000000";
					when "00110111100000010" => rgb <= "000000";
					when "00110111100000011" => rgb <= "000000";
					when "00110111100000100" => rgb <= "000000";
					when "00110111100000101" => rgb <= "000000";
					when "00110111100000110" => rgb <= "000000";
					when "00110111100000111" => rgb <= "000000";
					when "00110111100001000" => rgb <= "000000";
					when "00110111100001001" => rgb <= "000000";
					when "00110111100001010" => rgb <= "000000";
					when "00110111100001011" => rgb <= "000000";
					when "00110111100001100" => rgb <= "000000";
					when "00110111100001101" => rgb <= "000000";
					when "00110111100001110" => rgb <= "000000";
					when "00110111100001111" => rgb <= "000000";
					when "00110111100010000" => rgb <= "000000";
					when "00110111100010001" => rgb <= "000000";
					when "00110111100010010" => rgb <= "000000";
					when "00110111100010011" => rgb <= "000000";
					when "00110111100010100" => rgb <= "000000";
					when "00110111100010101" => rgb <= "000000";
					when "00110111100010110" => rgb <= "000000";
					when "00110111100010111" => rgb <= "000000";
					when "00110111100011000" => rgb <= "000000";
					when "00110111100011001" => rgb <= "000000";
					when "00110111100011010" => rgb <= "000000";
					when "00110111100011011" => rgb <= "000000";
					when "00110111100011100" => rgb <= "000000";
					when "00110111100011101" => rgb <= "000000";
					when "00110111100011110" => rgb <= "000000";
					when "00110111100011111" => rgb <= "000000";
					when "00110111100100000" => rgb <= "000000";
					when "00110111100100001" => rgb <= "000000";
					when "00110111100100010" => rgb <= "000000";
					when "00110111100100011" => rgb <= "000000";
					when "00110111100100100" => rgb <= "000000";
					when "00110111100100101" => rgb <= "000000";
					when "00110111100100110" => rgb <= "000000";
					when "00110111100100111" => rgb <= "000000";
					when "00110111100101000" => rgb <= "000000";
					when "00110111100101001" => rgb <= "000000";
					when "00110111100101010" => rgb <= "000000";
					when "00110111100101011" => rgb <= "000000";
					when "00110111100101100" => rgb <= "000000";
					when "00110111100101101" => rgb <= "000000";
					when "00110111100101110" => rgb <= "000000";
					when "00110111100101111" => rgb <= "000000";
					when "00110111100110000" => rgb <= "000000";
					when "00110111100110001" => rgb <= "000000";
					when "00110111100110010" => rgb <= "000000";
					when "00110111100110011" => rgb <= "000000";
					when "00110111100110100" => rgb <= "000000";
					when "00110111100110101" => rgb <= "000000";
					when "00110111100110110" => rgb <= "000000";
					when "00110111100110111" => rgb <= "000000";
					when "00110111100111000" => rgb <= "000000";
					when "00110111100111001" => rgb <= "000000";
					when "00110111100111010" => rgb <= "000000";
					when "00110111100111011" => rgb <= "000000";
					when "00110111100111100" => rgb <= "000000";
					when "00110111100111101" => rgb <= "000000";
					when "00110111100111110" => rgb <= "000000";
					when "00110111100111111" => rgb <= "000000";
					when "00111000000000000" => rgb <= "000000";
					when "00111000000000001" => rgb <= "000000";
					when "00111000000000010" => rgb <= "000000";
					when "00111000000000011" => rgb <= "000000";
					when "00111000000000100" => rgb <= "000000";
					when "00111000000000101" => rgb <= "000000";
					when "00111000000000110" => rgb <= "000000";
					when "00111000000000111" => rgb <= "000000";
					when "00111000000001000" => rgb <= "000000";
					when "00111000000001001" => rgb <= "000000";
					when "00111000000001010" => rgb <= "000000";
					when "00111000000001011" => rgb <= "000000";
					when "00111000000001100" => rgb <= "000000";
					when "00111000000001101" => rgb <= "000000";
					when "00111000000001110" => rgb <= "000000";
					when "00111000000001111" => rgb <= "000000";
					when "00111000000010000" => rgb <= "000000";
					when "00111000000010001" => rgb <= "000000";
					when "00111000000010010" => rgb <= "000000";
					when "00111000000010011" => rgb <= "000000";
					when "00111000000010100" => rgb <= "000000";
					when "00111000000010101" => rgb <= "000000";
					when "00111000000010110" => rgb <= "000000";
					when "00111000000010111" => rgb <= "000000";
					when "00111000000011000" => rgb <= "000000";
					when "00111000000011001" => rgb <= "000000";
					when "00111000000011010" => rgb <= "000000";
					when "00111000000011011" => rgb <= "000000";
					when "00111000000011100" => rgb <= "000000";
					when "00111000000011101" => rgb <= "000000";
					when "00111000000011110" => rgb <= "000000";
					when "00111000000011111" => rgb <= "000000";
					when "00111000000100000" => rgb <= "000000";
					when "00111000000100001" => rgb <= "000000";
					when "00111000000100010" => rgb <= "000000";
					when "00111000000100011" => rgb <= "000000";
					when "00111000000100100" => rgb <= "000000";
					when "00111000000100101" => rgb <= "000000";
					when "00111000000100110" => rgb <= "000000";
					when "00111000000100111" => rgb <= "000000";
					when "00111000000101000" => rgb <= "000000";
					when "00111000000101001" => rgb <= "000000";
					when "00111000000101010" => rgb <= "000000";
					when "00111000000101011" => rgb <= "000000";
					when "00111000000101100" => rgb <= "000000";
					when "00111000000101101" => rgb <= "000000";
					when "00111000000101110" => rgb <= "000000";
					when "00111000000101111" => rgb <= "000000";
					when "00111000000110000" => rgb <= "000000";
					when "00111000000110001" => rgb <= "000000";
					when "00111000000110010" => rgb <= "000000";
					when "00111000000110011" => rgb <= "000000";
					when "00111000000110100" => rgb <= "000000";
					when "00111000000110101" => rgb <= "000000";
					when "00111000000110110" => rgb <= "000000";
					when "00111000000110111" => rgb <= "000000";
					when "00111000000111000" => rgb <= "000000";
					when "00111000000111001" => rgb <= "000000";
					when "00111000000111010" => rgb <= "000000";
					when "00111000000111011" => rgb <= "000000";
					when "00111000000111100" => rgb <= "000000";
					when "00111000000111101" => rgb <= "000000";
					when "00111000000111110" => rgb <= "000000";
					when "00111000000111111" => rgb <= "000000";
					when "00111000001000000" => rgb <= "000000";
					when "00111000001000001" => rgb <= "000000";
					when "00111000001000010" => rgb <= "000000";
					when "00111000001000011" => rgb <= "000000";
					when "00111000001000100" => rgb <= "000000";
					when "00111000001000101" => rgb <= "000000";
					when "00111000001000110" => rgb <= "000000";
					when "00111000001000111" => rgb <= "000000";
					when "00111000001001000" => rgb <= "000000";
					when "00111000001001001" => rgb <= "000000";
					when "00111000001001010" => rgb <= "000000";
					when "00111000001001011" => rgb <= "000000";
					when "00111000001001100" => rgb <= "000000";
					when "00111000001001101" => rgb <= "000000";
					when "00111000001001110" => rgb <= "000000";
					when "00111000001001111" => rgb <= "000000";
					when "00111000001010000" => rgb <= "000000";
					when "00111000001010001" => rgb <= "000000";
					when "00111000001010010" => rgb <= "000000";
					when "00111000001010011" => rgb <= "000000";
					when "00111000001010100" => rgb <= "000000";
					when "00111000001010101" => rgb <= "000000";
					when "00111000001010110" => rgb <= "000000";
					when "00111000001010111" => rgb <= "000000";
					when "00111000001011000" => rgb <= "000000";
					when "00111000001011001" => rgb <= "000000";
					when "00111000001011010" => rgb <= "000000";
					when "00111000001011011" => rgb <= "000000";
					when "00111000001011100" => rgb <= "000000";
					when "00111000001011101" => rgb <= "000000";
					when "00111000001011110" => rgb <= "000000";
					when "00111000001011111" => rgb <= "000000";
					when "00111000001100000" => rgb <= "000000";
					when "00111000001100001" => rgb <= "000000";
					when "00111000001100010" => rgb <= "000000";
					when "00111000001100011" => rgb <= "000000";
					when "00111000001100100" => rgb <= "000000";
					when "00111000001100101" => rgb <= "000000";
					when "00111000001100110" => rgb <= "010100";
					when "00111000001100111" => rgb <= "101000";
					when "00111000001101000" => rgb <= "101000";
					when "00111000001101001" => rgb <= "101000";
					when "00111000001101010" => rgb <= "101000";
					when "00111000001101011" => rgb <= "101000";
					when "00111000001101100" => rgb <= "101000";
					when "00111000001101101" => rgb <= "101000";
					when "00111000001101110" => rgb <= "101000";
					when "00111000001101111" => rgb <= "101000";
					when "00111000001110000" => rgb <= "111000";
					when "00111000001110001" => rgb <= "100100";
					when "00111000001110010" => rgb <= "000000";
					when "00111000001110011" => rgb <= "000000";
					when "00111000001110100" => rgb <= "000000";
					when "00111000001110101" => rgb <= "000000";
					when "00111000001110110" => rgb <= "000000";
					when "00111000001110111" => rgb <= "000000";
					when "00111000001111000" => rgb <= "000000";
					when "00111000001111001" => rgb <= "000000";
					when "00111000001111010" => rgb <= "000000";
					when "00111000001111011" => rgb <= "000000";
					when "00111000001111100" => rgb <= "000000";
					when "00111000001111101" => rgb <= "101000";
					when "00111000001111110" => rgb <= "101000";
					when "00111000001111111" => rgb <= "101000";
					when "00111000010000000" => rgb <= "101000";
					when "00111000010000001" => rgb <= "101000";
					when "00111000010000010" => rgb <= "101000";
					when "00111000010000011" => rgb <= "101000";
					when "00111000010000100" => rgb <= "101000";
					when "00111000010000101" => rgb <= "101000";
					when "00111000010000110" => rgb <= "101000";
					when "00111000010000111" => rgb <= "101000";
					when "00111000010001000" => rgb <= "101000";
					when "00111000010001001" => rgb <= "101000";
					when "00111000010001010" => rgb <= "101000";
					when "00111000010001011" => rgb <= "101000";
					when "00111000010001100" => rgb <= "101000";
					when "00111000010001101" => rgb <= "101000";
					when "00111000010001110" => rgb <= "101000";
					when "00111000010001111" => rgb <= "101000";
					when "00111000010010000" => rgb <= "101000";
					when "00111000010010001" => rgb <= "101000";
					when "00111000010010010" => rgb <= "101000";
					when "00111000010010011" => rgb <= "101000";
					when "00111000010010100" => rgb <= "101000";
					when "00111000010010101" => rgb <= "101000";
					when "00111000010010110" => rgb <= "101000";
					when "00111000010010111" => rgb <= "101000";
					when "00111000010011000" => rgb <= "101000";
					when "00111000010011001" => rgb <= "101000";
					when "00111000010011010" => rgb <= "101000";
					when "00111000010011011" => rgb <= "101000";
					when "00111000010011100" => rgb <= "101000";
					when "00111000010011101" => rgb <= "101000";
					when "00111000010011110" => rgb <= "101000";
					when "00111000010011111" => rgb <= "101000";
					when "00111000010100000" => rgb <= "101000";
					when "00111000010100001" => rgb <= "101000";
					when "00111000010100010" => rgb <= "101000";
					when "00111000010100011" => rgb <= "101000";
					when "00111000010100100" => rgb <= "101000";
					when "00111000010100101" => rgb <= "101000";
					when "00111000010100110" => rgb <= "101000";
					when "00111000010100111" => rgb <= "101000";
					when "00111000010101000" => rgb <= "101000";
					when "00111000010101001" => rgb <= "101000";
					when "00111000010101010" => rgb <= "101000";
					when "00111000010101011" => rgb <= "101000";
					when "00111000010101100" => rgb <= "101000";
					when "00111000010101101" => rgb <= "101000";
					when "00111000010101110" => rgb <= "101000";
					when "00111000010101111" => rgb <= "101000";
					when "00111000010110000" => rgb <= "101000";
					when "00111000010110001" => rgb <= "101000";
					when "00111000010110010" => rgb <= "101000";
					when "00111000010110011" => rgb <= "101000";
					when "00111000010110100" => rgb <= "101000";
					when "00111000010110101" => rgb <= "101000";
					when "00111000010110110" => rgb <= "101000";
					when "00111000010110111" => rgb <= "101000";
					when "00111000010111000" => rgb <= "101000";
					when "00111000010111001" => rgb <= "101000";
					when "00111000010111010" => rgb <= "101000";
					when "00111000010111011" => rgb <= "101000";
					when "00111000010111100" => rgb <= "101000";
					when "00111000010111101" => rgb <= "101000";
					when "00111000010111110" => rgb <= "101000";
					when "00111000010111111" => rgb <= "101000";
					when "00111000011000000" => rgb <= "100100";
					when "00111000011000001" => rgb <= "000000";
					when "00111000011000010" => rgb <= "000000";
					when "00111000011000011" => rgb <= "000000";
					when "00111000011000100" => rgb <= "000000";
					when "00111000011000101" => rgb <= "000000";
					when "00111000011000110" => rgb <= "000000";
					when "00111000011000111" => rgb <= "000000";
					when "00111000011001000" => rgb <= "000000";
					when "00111000011001001" => rgb <= "000000";
					when "00111000011001010" => rgb <= "000000";
					when "00111000011001011" => rgb <= "000000";
					when "00111000011001100" => rgb <= "010100";
					when "00111000011001101" => rgb <= "101000";
					when "00111000011001110" => rgb <= "101000";
					when "00111000011001111" => rgb <= "101000";
					when "00111000011010000" => rgb <= "101000";
					when "00111000011010001" => rgb <= "101000";
					when "00111000011010010" => rgb <= "101000";
					when "00111000011010011" => rgb <= "101000";
					when "00111000011010100" => rgb <= "101000";
					when "00111000011010101" => rgb <= "101000";
					when "00111000011010110" => rgb <= "101000";
					when "00111000011010111" => rgb <= "010100";
					when "00111000011011000" => rgb <= "000000";
					when "00111000011011001" => rgb <= "000000";
					when "00111000011011010" => rgb <= "000000";
					when "00111000011011011" => rgb <= "000000";
					when "00111000011011100" => rgb <= "000000";
					when "00111000011011101" => rgb <= "000000";
					when "00111000011011110" => rgb <= "000000";
					when "00111000011011111" => rgb <= "000000";
					when "00111000011100000" => rgb <= "000000";
					when "00111000011100001" => rgb <= "000000";
					when "00111000011100010" => rgb <= "000000";
					when "00111000011100011" => rgb <= "000000";
					when "00111000011100100" => rgb <= "000000";
					when "00111000011100101" => rgb <= "000000";
					when "00111000011100110" => rgb <= "000000";
					when "00111000011100111" => rgb <= "000000";
					when "00111000011101000" => rgb <= "000000";
					when "00111000011101001" => rgb <= "000000";
					when "00111000011101010" => rgb <= "000000";
					when "00111000011101011" => rgb <= "000000";
					when "00111000011101100" => rgb <= "000000";
					when "00111000011101101" => rgb <= "000000";
					when "00111000011101110" => rgb <= "000000";
					when "00111000011101111" => rgb <= "000000";
					when "00111000011110000" => rgb <= "000000";
					when "00111000011110001" => rgb <= "000000";
					when "00111000011110010" => rgb <= "000000";
					when "00111000011110011" => rgb <= "000000";
					when "00111000011110100" => rgb <= "000000";
					when "00111000011110101" => rgb <= "000000";
					when "00111000011110110" => rgb <= "000000";
					when "00111000011110111" => rgb <= "000000";
					when "00111000011111000" => rgb <= "000000";
					when "00111000011111001" => rgb <= "000000";
					when "00111000011111010" => rgb <= "000000";
					when "00111000011111011" => rgb <= "000000";
					when "00111000011111100" => rgb <= "000000";
					when "00111000011111101" => rgb <= "000000";
					when "00111000011111110" => rgb <= "000000";
					when "00111000011111111" => rgb <= "000000";
					when "00111000100000000" => rgb <= "000000";
					when "00111000100000001" => rgb <= "000000";
					when "00111000100000010" => rgb <= "000000";
					when "00111000100000011" => rgb <= "000000";
					when "00111000100000100" => rgb <= "000000";
					when "00111000100000101" => rgb <= "000000";
					when "00111000100000110" => rgb <= "000000";
					when "00111000100000111" => rgb <= "000000";
					when "00111000100001000" => rgb <= "000000";
					when "00111000100001001" => rgb <= "000000";
					when "00111000100001010" => rgb <= "000000";
					when "00111000100001011" => rgb <= "000000";
					when "00111000100001100" => rgb <= "000000";
					when "00111000100001101" => rgb <= "000000";
					when "00111000100001110" => rgb <= "000000";
					when "00111000100001111" => rgb <= "000000";
					when "00111000100010000" => rgb <= "000000";
					when "00111000100010001" => rgb <= "000000";
					when "00111000100010010" => rgb <= "000000";
					when "00111000100010011" => rgb <= "000000";
					when "00111000100010100" => rgb <= "000000";
					when "00111000100010101" => rgb <= "000000";
					when "00111000100010110" => rgb <= "000000";
					when "00111000100010111" => rgb <= "000000";
					when "00111000100011000" => rgb <= "000000";
					when "00111000100011001" => rgb <= "000000";
					when "00111000100011010" => rgb <= "000000";
					when "00111000100011011" => rgb <= "000000";
					when "00111000100011100" => rgb <= "000000";
					when "00111000100011101" => rgb <= "000000";
					when "00111000100011110" => rgb <= "000000";
					when "00111000100011111" => rgb <= "000000";
					when "00111000100100000" => rgb <= "000000";
					when "00111000100100001" => rgb <= "000000";
					when "00111000100100010" => rgb <= "000000";
					when "00111000100100011" => rgb <= "000000";
					when "00111000100100100" => rgb <= "000000";
					when "00111000100100101" => rgb <= "000000";
					when "00111000100100110" => rgb <= "000000";
					when "00111000100100111" => rgb <= "000000";
					when "00111000100101000" => rgb <= "000000";
					when "00111000100101001" => rgb <= "000000";
					when "00111000100101010" => rgb <= "000000";
					when "00111000100101011" => rgb <= "000000";
					when "00111000100101100" => rgb <= "000000";
					when "00111000100101101" => rgb <= "000000";
					when "00111000100101110" => rgb <= "000000";
					when "00111000100101111" => rgb <= "000000";
					when "00111000100110000" => rgb <= "000000";
					when "00111000100110001" => rgb <= "000000";
					when "00111000100110010" => rgb <= "000000";
					when "00111000100110011" => rgb <= "000000";
					when "00111000100110100" => rgb <= "000000";
					when "00111000100110101" => rgb <= "000000";
					when "00111000100110110" => rgb <= "000000";
					when "00111000100110111" => rgb <= "000000";
					when "00111000100111000" => rgb <= "000000";
					when "00111000100111001" => rgb <= "000000";
					when "00111000100111010" => rgb <= "000000";
					when "00111000100111011" => rgb <= "000000";
					when "00111000100111100" => rgb <= "000000";
					when "00111000100111101" => rgb <= "000000";
					when "00111000100111110" => rgb <= "000000";
					when "00111000100111111" => rgb <= "000000";
					when "00111001000000000" => rgb <= "000000";
					when "00111001000000001" => rgb <= "000000";
					when "00111001000000010" => rgb <= "000000";
					when "00111001000000011" => rgb <= "000000";
					when "00111001000000100" => rgb <= "000000";
					when "00111001000000101" => rgb <= "000000";
					when "00111001000000110" => rgb <= "000000";
					when "00111001000000111" => rgb <= "000000";
					when "00111001000001000" => rgb <= "000000";
					when "00111001000001001" => rgb <= "000000";
					when "00111001000001010" => rgb <= "000000";
					when "00111001000001011" => rgb <= "000000";
					when "00111001000001100" => rgb <= "000000";
					when "00111001000001101" => rgb <= "000000";
					when "00111001000001110" => rgb <= "000000";
					when "00111001000001111" => rgb <= "000000";
					when "00111001000010000" => rgb <= "000000";
					when "00111001000010001" => rgb <= "000000";
					when "00111001000010010" => rgb <= "000000";
					when "00111001000010011" => rgb <= "000000";
					when "00111001000010100" => rgb <= "000000";
					when "00111001000010101" => rgb <= "000000";
					when "00111001000010110" => rgb <= "000000";
					when "00111001000010111" => rgb <= "000000";
					when "00111001000011000" => rgb <= "000000";
					when "00111001000011001" => rgb <= "000000";
					when "00111001000011010" => rgb <= "000000";
					when "00111001000011011" => rgb <= "000000";
					when "00111001000011100" => rgb <= "000000";
					when "00111001000011101" => rgb <= "000000";
					when "00111001000011110" => rgb <= "000000";
					when "00111001000011111" => rgb <= "000000";
					when "00111001000100000" => rgb <= "000000";
					when "00111001000100001" => rgb <= "000000";
					when "00111001000100010" => rgb <= "000000";
					when "00111001000100011" => rgb <= "000000";
					when "00111001000100100" => rgb <= "000000";
					when "00111001000100101" => rgb <= "000000";
					when "00111001000100110" => rgb <= "000000";
					when "00111001000100111" => rgb <= "000000";
					when "00111001000101000" => rgb <= "000000";
					when "00111001000101001" => rgb <= "000000";
					when "00111001000101010" => rgb <= "000000";
					when "00111001000101011" => rgb <= "000000";
					when "00111001000101100" => rgb <= "000000";
					when "00111001000101101" => rgb <= "000000";
					when "00111001000101110" => rgb <= "000000";
					when "00111001000101111" => rgb <= "000000";
					when "00111001000110000" => rgb <= "000000";
					when "00111001000110001" => rgb <= "000000";
					when "00111001000110010" => rgb <= "000000";
					when "00111001000110011" => rgb <= "000000";
					when "00111001000110100" => rgb <= "000000";
					when "00111001000110101" => rgb <= "000000";
					when "00111001000110110" => rgb <= "000000";
					when "00111001000110111" => rgb <= "000000";
					when "00111001000111000" => rgb <= "000000";
					when "00111001000111001" => rgb <= "000000";
					when "00111001000111010" => rgb <= "000000";
					when "00111001000111011" => rgb <= "000000";
					when "00111001000111100" => rgb <= "000000";
					when "00111001000111101" => rgb <= "000000";
					when "00111001000111110" => rgb <= "000000";
					when "00111001000111111" => rgb <= "000000";
					when "00111001001000000" => rgb <= "000000";
					when "00111001001000001" => rgb <= "000000";
					when "00111001001000010" => rgb <= "000000";
					when "00111001001000011" => rgb <= "000000";
					when "00111001001000100" => rgb <= "000000";
					when "00111001001000101" => rgb <= "000000";
					when "00111001001000110" => rgb <= "000000";
					when "00111001001000111" => rgb <= "000000";
					when "00111001001001000" => rgb <= "000000";
					when "00111001001001001" => rgb <= "000000";
					when "00111001001001010" => rgb <= "000000";
					when "00111001001001011" => rgb <= "000000";
					when "00111001001001100" => rgb <= "000000";
					when "00111001001001101" => rgb <= "000000";
					when "00111001001001110" => rgb <= "000000";
					when "00111001001001111" => rgb <= "000000";
					when "00111001001010000" => rgb <= "000000";
					when "00111001001010001" => rgb <= "000000";
					when "00111001001010010" => rgb <= "000000";
					when "00111001001010011" => rgb <= "000000";
					when "00111001001010100" => rgb <= "000000";
					when "00111001001010101" => rgb <= "000000";
					when "00111001001010110" => rgb <= "000000";
					when "00111001001010111" => rgb <= "000000";
					when "00111001001011000" => rgb <= "000000";
					when "00111001001011001" => rgb <= "000000";
					when "00111001001011010" => rgb <= "000000";
					when "00111001001011011" => rgb <= "000000";
					when "00111001001011100" => rgb <= "000000";
					when "00111001001011101" => rgb <= "000000";
					when "00111001001011110" => rgb <= "000000";
					when "00111001001011111" => rgb <= "000000";
					when "00111001001100000" => rgb <= "000000";
					when "00111001001100001" => rgb <= "000000";
					when "00111001001100010" => rgb <= "000000";
					when "00111001001100011" => rgb <= "000000";
					when "00111001001100100" => rgb <= "000000";
					when "00111001001100101" => rgb <= "000000";
					when "00111001001100110" => rgb <= "010100";
					when "00111001001100111" => rgb <= "111000";
					when "00111001001101000" => rgb <= "101000";
					when "00111001001101001" => rgb <= "101000";
					when "00111001001101010" => rgb <= "101000";
					when "00111001001101011" => rgb <= "101000";
					when "00111001001101100" => rgb <= "101000";
					when "00111001001101101" => rgb <= "101000";
					when "00111001001101110" => rgb <= "101000";
					when "00111001001101111" => rgb <= "101000";
					when "00111001001110000" => rgb <= "101000";
					when "00111001001110001" => rgb <= "100100";
					when "00111001001110010" => rgb <= "000000";
					when "00111001001110011" => rgb <= "000000";
					when "00111001001110100" => rgb <= "000000";
					when "00111001001110101" => rgb <= "000000";
					when "00111001001110110" => rgb <= "000000";
					when "00111001001110111" => rgb <= "000000";
					when "00111001001111000" => rgb <= "000000";
					when "00111001001111001" => rgb <= "000000";
					when "00111001001111010" => rgb <= "000000";
					when "00111001001111011" => rgb <= "000000";
					when "00111001001111100" => rgb <= "000000";
					when "00111001001111101" => rgb <= "101000";
					when "00111001001111110" => rgb <= "101000";
					when "00111001001111111" => rgb <= "101000";
					when "00111001010000000" => rgb <= "101000";
					when "00111001010000001" => rgb <= "101000";
					when "00111001010000010" => rgb <= "101000";
					when "00111001010000011" => rgb <= "101000";
					when "00111001010000100" => rgb <= "101000";
					when "00111001010000101" => rgb <= "101000";
					when "00111001010000110" => rgb <= "101000";
					when "00111001010000111" => rgb <= "101000";
					when "00111001010001000" => rgb <= "101000";
					when "00111001010001001" => rgb <= "101000";
					when "00111001010001010" => rgb <= "101000";
					when "00111001010001011" => rgb <= "101000";
					when "00111001010001100" => rgb <= "101000";
					when "00111001010001101" => rgb <= "101000";
					when "00111001010001110" => rgb <= "101000";
					when "00111001010001111" => rgb <= "101000";
					when "00111001010010000" => rgb <= "101000";
					when "00111001010010001" => rgb <= "101000";
					when "00111001010010010" => rgb <= "101000";
					when "00111001010010011" => rgb <= "101000";
					when "00111001010010100" => rgb <= "101000";
					when "00111001010010101" => rgb <= "101000";
					when "00111001010010110" => rgb <= "101000";
					when "00111001010010111" => rgb <= "101000";
					when "00111001010011000" => rgb <= "101000";
					when "00111001010011001" => rgb <= "101000";
					when "00111001010011010" => rgb <= "101000";
					when "00111001010011011" => rgb <= "101000";
					when "00111001010011100" => rgb <= "101000";
					when "00111001010011101" => rgb <= "101000";
					when "00111001010011110" => rgb <= "101000";
					when "00111001010011111" => rgb <= "101000";
					when "00111001010100000" => rgb <= "101000";
					when "00111001010100001" => rgb <= "101000";
					when "00111001010100010" => rgb <= "101000";
					when "00111001010100011" => rgb <= "101000";
					when "00111001010100100" => rgb <= "101000";
					when "00111001010100101" => rgb <= "101000";
					when "00111001010100110" => rgb <= "101000";
					when "00111001010100111" => rgb <= "101000";
					when "00111001010101000" => rgb <= "101000";
					when "00111001010101001" => rgb <= "101000";
					when "00111001010101010" => rgb <= "101000";
					when "00111001010101011" => rgb <= "101000";
					when "00111001010101100" => rgb <= "101000";
					when "00111001010101101" => rgb <= "101000";
					when "00111001010101110" => rgb <= "101000";
					when "00111001010101111" => rgb <= "101000";
					when "00111001010110000" => rgb <= "101000";
					when "00111001010110001" => rgb <= "101000";
					when "00111001010110010" => rgb <= "101000";
					when "00111001010110011" => rgb <= "101000";
					when "00111001010110100" => rgb <= "101000";
					when "00111001010110101" => rgb <= "101000";
					when "00111001010110110" => rgb <= "101000";
					when "00111001010110111" => rgb <= "101000";
					when "00111001010111000" => rgb <= "101000";
					when "00111001010111001" => rgb <= "101000";
					when "00111001010111010" => rgb <= "101000";
					when "00111001010111011" => rgb <= "101000";
					when "00111001010111100" => rgb <= "101000";
					when "00111001010111101" => rgb <= "101000";
					when "00111001010111110" => rgb <= "101000";
					when "00111001010111111" => rgb <= "101000";
					when "00111001011000000" => rgb <= "100100";
					when "00111001011000001" => rgb <= "000000";
					when "00111001011000010" => rgb <= "000000";
					when "00111001011000011" => rgb <= "000000";
					when "00111001011000100" => rgb <= "000000";
					when "00111001011000101" => rgb <= "000000";
					when "00111001011000110" => rgb <= "000000";
					when "00111001011000111" => rgb <= "000000";
					when "00111001011001000" => rgb <= "000000";
					when "00111001011001001" => rgb <= "000000";
					when "00111001011001010" => rgb <= "000000";
					when "00111001011001011" => rgb <= "000000";
					when "00111001011001100" => rgb <= "010100";
					when "00111001011001101" => rgb <= "101000";
					when "00111001011001110" => rgb <= "101000";
					when "00111001011001111" => rgb <= "101000";
					when "00111001011010000" => rgb <= "101000";
					when "00111001011010001" => rgb <= "101000";
					when "00111001011010010" => rgb <= "101000";
					when "00111001011010011" => rgb <= "101000";
					when "00111001011010100" => rgb <= "101000";
					when "00111001011010101" => rgb <= "101000";
					when "00111001011010110" => rgb <= "101000";
					when "00111001011010111" => rgb <= "010100";
					when "00111001011011000" => rgb <= "000000";
					when "00111001011011001" => rgb <= "000000";
					when "00111001011011010" => rgb <= "000000";
					when "00111001011011011" => rgb <= "000000";
					when "00111001011011100" => rgb <= "000000";
					when "00111001011011101" => rgb <= "000000";
					when "00111001011011110" => rgb <= "000000";
					when "00111001011011111" => rgb <= "000000";
					when "00111001011100000" => rgb <= "000000";
					when "00111001011100001" => rgb <= "000000";
					when "00111001011100010" => rgb <= "000000";
					when "00111001011100011" => rgb <= "000000";
					when "00111001011100100" => rgb <= "000000";
					when "00111001011100101" => rgb <= "000000";
					when "00111001011100110" => rgb <= "000000";
					when "00111001011100111" => rgb <= "000000";
					when "00111001011101000" => rgb <= "000000";
					when "00111001011101001" => rgb <= "000000";
					when "00111001011101010" => rgb <= "000000";
					when "00111001011101011" => rgb <= "000000";
					when "00111001011101100" => rgb <= "000000";
					when "00111001011101101" => rgb <= "000000";
					when "00111001011101110" => rgb <= "000000";
					when "00111001011101111" => rgb <= "000000";
					when "00111001011110000" => rgb <= "000000";
					when "00111001011110001" => rgb <= "000000";
					when "00111001011110010" => rgb <= "000000";
					when "00111001011110011" => rgb <= "000000";
					when "00111001011110100" => rgb <= "000000";
					when "00111001011110101" => rgb <= "000000";
					when "00111001011110110" => rgb <= "000000";
					when "00111001011110111" => rgb <= "000000";
					when "00111001011111000" => rgb <= "000000";
					when "00111001011111001" => rgb <= "000000";
					when "00111001011111010" => rgb <= "000000";
					when "00111001011111011" => rgb <= "000000";
					when "00111001011111100" => rgb <= "000000";
					when "00111001011111101" => rgb <= "000000";
					when "00111001011111110" => rgb <= "000000";
					when "00111001011111111" => rgb <= "000000";
					when "00111001100000000" => rgb <= "000000";
					when "00111001100000001" => rgb <= "000000";
					when "00111001100000010" => rgb <= "000000";
					when "00111001100000011" => rgb <= "000000";
					when "00111001100000100" => rgb <= "000000";
					when "00111001100000101" => rgb <= "000000";
					when "00111001100000110" => rgb <= "000000";
					when "00111001100000111" => rgb <= "000000";
					when "00111001100001000" => rgb <= "000000";
					when "00111001100001001" => rgb <= "000000";
					when "00111001100001010" => rgb <= "000000";
					when "00111001100001011" => rgb <= "000000";
					when "00111001100001100" => rgb <= "000000";
					when "00111001100001101" => rgb <= "000000";
					when "00111001100001110" => rgb <= "000000";
					when "00111001100001111" => rgb <= "000000";
					when "00111001100010000" => rgb <= "000000";
					when "00111001100010001" => rgb <= "000000";
					when "00111001100010010" => rgb <= "000000";
					when "00111001100010011" => rgb <= "000000";
					when "00111001100010100" => rgb <= "000000";
					when "00111001100010101" => rgb <= "000000";
					when "00111001100010110" => rgb <= "000000";
					when "00111001100010111" => rgb <= "000000";
					when "00111001100011000" => rgb <= "000000";
					when "00111001100011001" => rgb <= "000000";
					when "00111001100011010" => rgb <= "000000";
					when "00111001100011011" => rgb <= "000000";
					when "00111001100011100" => rgb <= "000000";
					when "00111001100011101" => rgb <= "000000";
					when "00111001100011110" => rgb <= "000000";
					when "00111001100011111" => rgb <= "000000";
					when "00111001100100000" => rgb <= "000000";
					when "00111001100100001" => rgb <= "000000";
					when "00111001100100010" => rgb <= "000000";
					when "00111001100100011" => rgb <= "000000";
					when "00111001100100100" => rgb <= "000000";
					when "00111001100100101" => rgb <= "000000";
					when "00111001100100110" => rgb <= "000000";
					when "00111001100100111" => rgb <= "000000";
					when "00111001100101000" => rgb <= "000000";
					when "00111001100101001" => rgb <= "000000";
					when "00111001100101010" => rgb <= "000000";
					when "00111001100101011" => rgb <= "000000";
					when "00111001100101100" => rgb <= "000000";
					when "00111001100101101" => rgb <= "000000";
					when "00111001100101110" => rgb <= "000000";
					when "00111001100101111" => rgb <= "000000";
					when "00111001100110000" => rgb <= "000000";
					when "00111001100110001" => rgb <= "000000";
					when "00111001100110010" => rgb <= "000000";
					when "00111001100110011" => rgb <= "000000";
					when "00111001100110100" => rgb <= "000000";
					when "00111001100110101" => rgb <= "000000";
					when "00111001100110110" => rgb <= "000000";
					when "00111001100110111" => rgb <= "000000";
					when "00111001100111000" => rgb <= "000000";
					when "00111001100111001" => rgb <= "000000";
					when "00111001100111010" => rgb <= "000000";
					when "00111001100111011" => rgb <= "000000";
					when "00111001100111100" => rgb <= "000000";
					when "00111001100111101" => rgb <= "000000";
					when "00111001100111110" => rgb <= "000000";
					when "00111001100111111" => rgb <= "000000";
					when "00111010000000000" => rgb <= "000000";
					when "00111010000000001" => rgb <= "000000";
					when "00111010000000010" => rgb <= "000000";
					when "00111010000000011" => rgb <= "000000";
					when "00111010000000100" => rgb <= "000000";
					when "00111010000000101" => rgb <= "000000";
					when "00111010000000110" => rgb <= "000000";
					when "00111010000000111" => rgb <= "000000";
					when "00111010000001000" => rgb <= "000000";
					when "00111010000001001" => rgb <= "000000";
					when "00111010000001010" => rgb <= "000000";
					when "00111010000001011" => rgb <= "000000";
					when "00111010000001100" => rgb <= "000000";
					when "00111010000001101" => rgb <= "000000";
					when "00111010000001110" => rgb <= "000000";
					when "00111010000001111" => rgb <= "000000";
					when "00111010000010000" => rgb <= "000000";
					when "00111010000010001" => rgb <= "000000";
					when "00111010000010010" => rgb <= "000000";
					when "00111010000010011" => rgb <= "000000";
					when "00111010000010100" => rgb <= "000000";
					when "00111010000010101" => rgb <= "000000";
					when "00111010000010110" => rgb <= "000000";
					when "00111010000010111" => rgb <= "000000";
					when "00111010000011000" => rgb <= "000000";
					when "00111010000011001" => rgb <= "000000";
					when "00111010000011010" => rgb <= "000000";
					when "00111010000011011" => rgb <= "000000";
					when "00111010000011100" => rgb <= "000000";
					when "00111010000011101" => rgb <= "000000";
					when "00111010000011110" => rgb <= "000000";
					when "00111010000011111" => rgb <= "000000";
					when "00111010000100000" => rgb <= "000000";
					when "00111010000100001" => rgb <= "000000";
					when "00111010000100010" => rgb <= "000000";
					when "00111010000100011" => rgb <= "000000";
					when "00111010000100100" => rgb <= "000000";
					when "00111010000100101" => rgb <= "000000";
					when "00111010000100110" => rgb <= "000000";
					when "00111010000100111" => rgb <= "000000";
					when "00111010000101000" => rgb <= "000000";
					when "00111010000101001" => rgb <= "000000";
					when "00111010000101010" => rgb <= "000000";
					when "00111010000101011" => rgb <= "000000";
					when "00111010000101100" => rgb <= "000000";
					when "00111010000101101" => rgb <= "000000";
					when "00111010000101110" => rgb <= "000000";
					when "00111010000101111" => rgb <= "000000";
					when "00111010000110000" => rgb <= "000000";
					when "00111010000110001" => rgb <= "000000";
					when "00111010000110010" => rgb <= "000000";
					when "00111010000110011" => rgb <= "000000";
					when "00111010000110100" => rgb <= "000000";
					when "00111010000110101" => rgb <= "000000";
					when "00111010000110110" => rgb <= "000000";
					when "00111010000110111" => rgb <= "000000";
					when "00111010000111000" => rgb <= "000000";
					when "00111010000111001" => rgb <= "000000";
					when "00111010000111010" => rgb <= "000000";
					when "00111010000111011" => rgb <= "000000";
					when "00111010000111100" => rgb <= "000000";
					when "00111010000111101" => rgb <= "000000";
					when "00111010000111110" => rgb <= "000000";
					when "00111010000111111" => rgb <= "000000";
					when "00111010001000000" => rgb <= "000000";
					when "00111010001000001" => rgb <= "000000";
					when "00111010001000010" => rgb <= "000000";
					when "00111010001000011" => rgb <= "000000";
					when "00111010001000100" => rgb <= "000000";
					when "00111010001000101" => rgb <= "000000";
					when "00111010001000110" => rgb <= "000000";
					when "00111010001000111" => rgb <= "000000";
					when "00111010001001000" => rgb <= "000000";
					when "00111010001001001" => rgb <= "000000";
					when "00111010001001010" => rgb <= "000000";
					when "00111010001001011" => rgb <= "000000";
					when "00111010001001100" => rgb <= "000000";
					when "00111010001001101" => rgb <= "000000";
					when "00111010001001110" => rgb <= "000000";
					when "00111010001001111" => rgb <= "000000";
					when "00111010001010000" => rgb <= "000000";
					when "00111010001010001" => rgb <= "000000";
					when "00111010001010010" => rgb <= "000000";
					when "00111010001010011" => rgb <= "000000";
					when "00111010001010100" => rgb <= "000000";
					when "00111010001010101" => rgb <= "000000";
					when "00111010001010110" => rgb <= "000000";
					when "00111010001010111" => rgb <= "000000";
					when "00111010001011000" => rgb <= "000000";
					when "00111010001011001" => rgb <= "000000";
					when "00111010001011010" => rgb <= "000000";
					when "00111010001011011" => rgb <= "000000";
					when "00111010001011100" => rgb <= "000000";
					when "00111010001011101" => rgb <= "000000";
					when "00111010001011110" => rgb <= "000000";
					when "00111010001011111" => rgb <= "000000";
					when "00111010001100000" => rgb <= "000000";
					when "00111010001100001" => rgb <= "000000";
					when "00111010001100010" => rgb <= "000000";
					when "00111010001100011" => rgb <= "000000";
					when "00111010001100100" => rgb <= "000000";
					when "00111010001100101" => rgb <= "000000";
					when "00111010001100110" => rgb <= "010100";
					when "00111010001100111" => rgb <= "111000";
					when "00111010001101000" => rgb <= "101000";
					when "00111010001101001" => rgb <= "101000";
					when "00111010001101010" => rgb <= "101000";
					when "00111010001101011" => rgb <= "101000";
					when "00111010001101100" => rgb <= "101000";
					when "00111010001101101" => rgb <= "101000";
					when "00111010001101110" => rgb <= "101000";
					when "00111010001101111" => rgb <= "101000";
					when "00111010001110000" => rgb <= "101000";
					when "00111010001110001" => rgb <= "100100";
					when "00111010001110010" => rgb <= "000000";
					when "00111010001110011" => rgb <= "000000";
					when "00111010001110100" => rgb <= "000000";
					when "00111010001110101" => rgb <= "000000";
					when "00111010001110110" => rgb <= "000000";
					when "00111010001110111" => rgb <= "000000";
					when "00111010001111000" => rgb <= "000000";
					when "00111010001111001" => rgb <= "000000";
					when "00111010001111010" => rgb <= "000000";
					when "00111010001111011" => rgb <= "000000";
					when "00111010001111100" => rgb <= "000000";
					when "00111010001111101" => rgb <= "101000";
					when "00111010001111110" => rgb <= "101000";
					when "00111010001111111" => rgb <= "101000";
					when "00111010010000000" => rgb <= "101000";
					when "00111010010000001" => rgb <= "101000";
					when "00111010010000010" => rgb <= "101000";
					when "00111010010000011" => rgb <= "101000";
					when "00111010010000100" => rgb <= "101000";
					when "00111010010000101" => rgb <= "101000";
					when "00111010010000110" => rgb <= "101000";
					when "00111010010000111" => rgb <= "101000";
					when "00111010010001000" => rgb <= "101000";
					when "00111010010001001" => rgb <= "101000";
					when "00111010010001010" => rgb <= "101000";
					when "00111010010001011" => rgb <= "101000";
					when "00111010010001100" => rgb <= "101000";
					when "00111010010001101" => rgb <= "101000";
					when "00111010010001110" => rgb <= "101000";
					when "00111010010001111" => rgb <= "101000";
					when "00111010010010000" => rgb <= "101000";
					when "00111010010010001" => rgb <= "101000";
					when "00111010010010010" => rgb <= "101000";
					when "00111010010010011" => rgb <= "101000";
					when "00111010010010100" => rgb <= "101000";
					when "00111010010010101" => rgb <= "101000";
					when "00111010010010110" => rgb <= "101000";
					when "00111010010010111" => rgb <= "101000";
					when "00111010010011000" => rgb <= "101000";
					when "00111010010011001" => rgb <= "101000";
					when "00111010010011010" => rgb <= "101000";
					when "00111010010011011" => rgb <= "101000";
					when "00111010010011100" => rgb <= "101000";
					when "00111010010011101" => rgb <= "101000";
					when "00111010010011110" => rgb <= "101000";
					when "00111010010011111" => rgb <= "101000";
					when "00111010010100000" => rgb <= "101000";
					when "00111010010100001" => rgb <= "101000";
					when "00111010010100010" => rgb <= "101000";
					when "00111010010100011" => rgb <= "101000";
					when "00111010010100100" => rgb <= "101000";
					when "00111010010100101" => rgb <= "101000";
					when "00111010010100110" => rgb <= "101000";
					when "00111010010100111" => rgb <= "101000";
					when "00111010010101000" => rgb <= "101000";
					when "00111010010101001" => rgb <= "101000";
					when "00111010010101010" => rgb <= "101000";
					when "00111010010101011" => rgb <= "101000";
					when "00111010010101100" => rgb <= "101000";
					when "00111010010101101" => rgb <= "101000";
					when "00111010010101110" => rgb <= "101000";
					when "00111010010101111" => rgb <= "101000";
					when "00111010010110000" => rgb <= "101000";
					when "00111010010110001" => rgb <= "101000";
					when "00111010010110010" => rgb <= "101000";
					when "00111010010110011" => rgb <= "101000";
					when "00111010010110100" => rgb <= "101000";
					when "00111010010110101" => rgb <= "101000";
					when "00111010010110110" => rgb <= "101000";
					when "00111010010110111" => rgb <= "101000";
					when "00111010010111000" => rgb <= "101000";
					when "00111010010111001" => rgb <= "101000";
					when "00111010010111010" => rgb <= "101000";
					when "00111010010111011" => rgb <= "101000";
					when "00111010010111100" => rgb <= "101000";
					when "00111010010111101" => rgb <= "101000";
					when "00111010010111110" => rgb <= "101000";
					when "00111010010111111" => rgb <= "101000";
					when "00111010011000000" => rgb <= "100100";
					when "00111010011000001" => rgb <= "000000";
					when "00111010011000010" => rgb <= "000000";
					when "00111010011000011" => rgb <= "000000";
					when "00111010011000100" => rgb <= "000000";
					when "00111010011000101" => rgb <= "000000";
					when "00111010011000110" => rgb <= "000000";
					when "00111010011000111" => rgb <= "000000";
					when "00111010011001000" => rgb <= "000000";
					when "00111010011001001" => rgb <= "000000";
					when "00111010011001010" => rgb <= "000000";
					when "00111010011001011" => rgb <= "000000";
					when "00111010011001100" => rgb <= "100100";
					when "00111010011001101" => rgb <= "101000";
					when "00111010011001110" => rgb <= "101000";
					when "00111010011001111" => rgb <= "101000";
					when "00111010011010000" => rgb <= "101000";
					when "00111010011010001" => rgb <= "101000";
					when "00111010011010010" => rgb <= "101000";
					when "00111010011010011" => rgb <= "101000";
					when "00111010011010100" => rgb <= "101000";
					when "00111010011010101" => rgb <= "101000";
					when "00111010011010110" => rgb <= "101000";
					when "00111010011010111" => rgb <= "010100";
					when "00111010011011000" => rgb <= "000000";
					when "00111010011011001" => rgb <= "000000";
					when "00111010011011010" => rgb <= "000000";
					when "00111010011011011" => rgb <= "000000";
					when "00111010011011100" => rgb <= "000000";
					when "00111010011011101" => rgb <= "000000";
					when "00111010011011110" => rgb <= "000000";
					when "00111010011011111" => rgb <= "000000";
					when "00111010011100000" => rgb <= "000000";
					when "00111010011100001" => rgb <= "000000";
					when "00111010011100010" => rgb <= "000000";
					when "00111010011100011" => rgb <= "000000";
					when "00111010011100100" => rgb <= "000000";
					when "00111010011100101" => rgb <= "000000";
					when "00111010011100110" => rgb <= "000000";
					when "00111010011100111" => rgb <= "000000";
					when "00111010011101000" => rgb <= "000000";
					when "00111010011101001" => rgb <= "000000";
					when "00111010011101010" => rgb <= "000000";
					when "00111010011101011" => rgb <= "000000";
					when "00111010011101100" => rgb <= "000000";
					when "00111010011101101" => rgb <= "000000";
					when "00111010011101110" => rgb <= "000000";
					when "00111010011101111" => rgb <= "000000";
					when "00111010011110000" => rgb <= "000000";
					when "00111010011110001" => rgb <= "000000";
					when "00111010011110010" => rgb <= "000000";
					when "00111010011110011" => rgb <= "000000";
					when "00111010011110100" => rgb <= "000000";
					when "00111010011110101" => rgb <= "000000";
					when "00111010011110110" => rgb <= "000000";
					when "00111010011110111" => rgb <= "000000";
					when "00111010011111000" => rgb <= "000000";
					when "00111010011111001" => rgb <= "000000";
					when "00111010011111010" => rgb <= "000000";
					when "00111010011111011" => rgb <= "000000";
					when "00111010011111100" => rgb <= "000000";
					when "00111010011111101" => rgb <= "000000";
					when "00111010011111110" => rgb <= "000000";
					when "00111010011111111" => rgb <= "000000";
					when "00111010100000000" => rgb <= "000000";
					when "00111010100000001" => rgb <= "000000";
					when "00111010100000010" => rgb <= "000000";
					when "00111010100000011" => rgb <= "000000";
					when "00111010100000100" => rgb <= "000000";
					when "00111010100000101" => rgb <= "000000";
					when "00111010100000110" => rgb <= "000000";
					when "00111010100000111" => rgb <= "000000";
					when "00111010100001000" => rgb <= "000000";
					when "00111010100001001" => rgb <= "000000";
					when "00111010100001010" => rgb <= "000000";
					when "00111010100001011" => rgb <= "000000";
					when "00111010100001100" => rgb <= "000000";
					when "00111010100001101" => rgb <= "000000";
					when "00111010100001110" => rgb <= "000000";
					when "00111010100001111" => rgb <= "000000";
					when "00111010100010000" => rgb <= "000000";
					when "00111010100010001" => rgb <= "000000";
					when "00111010100010010" => rgb <= "000000";
					when "00111010100010011" => rgb <= "000000";
					when "00111010100010100" => rgb <= "000000";
					when "00111010100010101" => rgb <= "000000";
					when "00111010100010110" => rgb <= "000000";
					when "00111010100010111" => rgb <= "000000";
					when "00111010100011000" => rgb <= "000000";
					when "00111010100011001" => rgb <= "000000";
					when "00111010100011010" => rgb <= "000000";
					when "00111010100011011" => rgb <= "000000";
					when "00111010100011100" => rgb <= "000000";
					when "00111010100011101" => rgb <= "000000";
					when "00111010100011110" => rgb <= "000000";
					when "00111010100011111" => rgb <= "000000";
					when "00111010100100000" => rgb <= "000000";
					when "00111010100100001" => rgb <= "000000";
					when "00111010100100010" => rgb <= "000000";
					when "00111010100100011" => rgb <= "000000";
					when "00111010100100100" => rgb <= "000000";
					when "00111010100100101" => rgb <= "000000";
					when "00111010100100110" => rgb <= "000000";
					when "00111010100100111" => rgb <= "000000";
					when "00111010100101000" => rgb <= "000000";
					when "00111010100101001" => rgb <= "000000";
					when "00111010100101010" => rgb <= "000000";
					when "00111010100101011" => rgb <= "000000";
					when "00111010100101100" => rgb <= "000000";
					when "00111010100101101" => rgb <= "000000";
					when "00111010100101110" => rgb <= "000000";
					when "00111010100101111" => rgb <= "000000";
					when "00111010100110000" => rgb <= "000000";
					when "00111010100110001" => rgb <= "000000";
					when "00111010100110010" => rgb <= "000000";
					when "00111010100110011" => rgb <= "000000";
					when "00111010100110100" => rgb <= "000000";
					when "00111010100110101" => rgb <= "000000";
					when "00111010100110110" => rgb <= "000000";
					when "00111010100110111" => rgb <= "000000";
					when "00111010100111000" => rgb <= "000000";
					when "00111010100111001" => rgb <= "000000";
					when "00111010100111010" => rgb <= "000000";
					when "00111010100111011" => rgb <= "000000";
					when "00111010100111100" => rgb <= "000000";
					when "00111010100111101" => rgb <= "000000";
					when "00111010100111110" => rgb <= "000000";
					when "00111010100111111" => rgb <= "000000";
					when "00111011000000000" => rgb <= "000000";
					when "00111011000000001" => rgb <= "000000";
					when "00111011000000010" => rgb <= "000000";
					when "00111011000000011" => rgb <= "000000";
					when "00111011000000100" => rgb <= "000000";
					when "00111011000000101" => rgb <= "000000";
					when "00111011000000110" => rgb <= "000000";
					when "00111011000000111" => rgb <= "000000";
					when "00111011000001000" => rgb <= "000000";
					when "00111011000001001" => rgb <= "000000";
					when "00111011000001010" => rgb <= "000000";
					when "00111011000001011" => rgb <= "000000";
					when "00111011000001100" => rgb <= "000000";
					when "00111011000001101" => rgb <= "000000";
					when "00111011000001110" => rgb <= "000000";
					when "00111011000001111" => rgb <= "000000";
					when "00111011000010000" => rgb <= "000000";
					when "00111011000010001" => rgb <= "000000";
					when "00111011000010010" => rgb <= "000000";
					when "00111011000010011" => rgb <= "000000";
					when "00111011000010100" => rgb <= "000000";
					when "00111011000010101" => rgb <= "000000";
					when "00111011000010110" => rgb <= "000000";
					when "00111011000010111" => rgb <= "000000";
					when "00111011000011000" => rgb <= "000000";
					when "00111011000011001" => rgb <= "000000";
					when "00111011000011010" => rgb <= "000000";
					when "00111011000011011" => rgb <= "000000";
					when "00111011000011100" => rgb <= "000000";
					when "00111011000011101" => rgb <= "000000";
					when "00111011000011110" => rgb <= "000000";
					when "00111011000011111" => rgb <= "000000";
					when "00111011000100000" => rgb <= "000000";
					when "00111011000100001" => rgb <= "000000";
					when "00111011000100010" => rgb <= "000000";
					when "00111011000100011" => rgb <= "000000";
					when "00111011000100100" => rgb <= "000000";
					when "00111011000100101" => rgb <= "000000";
					when "00111011000100110" => rgb <= "000000";
					when "00111011000100111" => rgb <= "000000";
					when "00111011000101000" => rgb <= "000000";
					when "00111011000101001" => rgb <= "000000";
					when "00111011000101010" => rgb <= "000000";
					when "00111011000101011" => rgb <= "000000";
					when "00111011000101100" => rgb <= "000000";
					when "00111011000101101" => rgb <= "000000";
					when "00111011000101110" => rgb <= "000000";
					when "00111011000101111" => rgb <= "000000";
					when "00111011000110000" => rgb <= "000000";
					when "00111011000110001" => rgb <= "000000";
					when "00111011000110010" => rgb <= "000000";
					when "00111011000110011" => rgb <= "000000";
					when "00111011000110100" => rgb <= "000000";
					when "00111011000110101" => rgb <= "000000";
					when "00111011000110110" => rgb <= "000000";
					when "00111011000110111" => rgb <= "000000";
					when "00111011000111000" => rgb <= "000000";
					when "00111011000111001" => rgb <= "000000";
					when "00111011000111010" => rgb <= "000000";
					when "00111011000111011" => rgb <= "000000";
					when "00111011000111100" => rgb <= "000000";
					when "00111011000111101" => rgb <= "000000";
					when "00111011000111110" => rgb <= "000000";
					when "00111011000111111" => rgb <= "000000";
					when "00111011001000000" => rgb <= "000000";
					when "00111011001000001" => rgb <= "000000";
					when "00111011001000010" => rgb <= "000000";
					when "00111011001000011" => rgb <= "000000";
					when "00111011001000100" => rgb <= "000000";
					when "00111011001000101" => rgb <= "000000";
					when "00111011001000110" => rgb <= "000000";
					when "00111011001000111" => rgb <= "000000";
					when "00111011001001000" => rgb <= "000000";
					when "00111011001001001" => rgb <= "000000";
					when "00111011001001010" => rgb <= "000000";
					when "00111011001001011" => rgb <= "000000";
					when "00111011001001100" => rgb <= "000000";
					when "00111011001001101" => rgb <= "000000";
					when "00111011001001110" => rgb <= "000000";
					when "00111011001001111" => rgb <= "000000";
					when "00111011001010000" => rgb <= "000000";
					when "00111011001010001" => rgb <= "000000";
					when "00111011001010010" => rgb <= "000000";
					when "00111011001010011" => rgb <= "000000";
					when "00111011001010100" => rgb <= "000000";
					when "00111011001010101" => rgb <= "000000";
					when "00111011001010110" => rgb <= "000000";
					when "00111011001010111" => rgb <= "000000";
					when "00111011001011000" => rgb <= "000000";
					when "00111011001011001" => rgb <= "000000";
					when "00111011001011010" => rgb <= "000000";
					when "00111011001011011" => rgb <= "000000";
					when "00111011001011100" => rgb <= "000000";
					when "00111011001011101" => rgb <= "000000";
					when "00111011001011110" => rgb <= "000000";
					when "00111011001011111" => rgb <= "000000";
					when "00111011001100000" => rgb <= "000000";
					when "00111011001100001" => rgb <= "000000";
					when "00111011001100010" => rgb <= "000000";
					when "00111011001100011" => rgb <= "000000";
					when "00111011001100100" => rgb <= "000000";
					when "00111011001100101" => rgb <= "000000";
					when "00111011001100110" => rgb <= "010100";
					when "00111011001100111" => rgb <= "111000";
					when "00111011001101000" => rgb <= "101000";
					when "00111011001101001" => rgb <= "101000";
					when "00111011001101010" => rgb <= "101000";
					when "00111011001101011" => rgb <= "101000";
					when "00111011001101100" => rgb <= "101000";
					when "00111011001101101" => rgb <= "101000";
					when "00111011001101110" => rgb <= "101000";
					when "00111011001101111" => rgb <= "101000";
					when "00111011001110000" => rgb <= "101000";
					when "00111011001110001" => rgb <= "100100";
					when "00111011001110010" => rgb <= "000000";
					when "00111011001110011" => rgb <= "000000";
					when "00111011001110100" => rgb <= "000000";
					when "00111011001110101" => rgb <= "000000";
					when "00111011001110110" => rgb <= "000000";
					when "00111011001110111" => rgb <= "000000";
					when "00111011001111000" => rgb <= "000000";
					when "00111011001111001" => rgb <= "000000";
					when "00111011001111010" => rgb <= "000000";
					when "00111011001111011" => rgb <= "000000";
					when "00111011001111100" => rgb <= "000000";
					when "00111011001111101" => rgb <= "101000";
					when "00111011001111110" => rgb <= "101000";
					when "00111011001111111" => rgb <= "101000";
					when "00111011010000000" => rgb <= "101000";
					when "00111011010000001" => rgb <= "101000";
					when "00111011010000010" => rgb <= "101000";
					when "00111011010000011" => rgb <= "101000";
					when "00111011010000100" => rgb <= "101000";
					when "00111011010000101" => rgb <= "101000";
					when "00111011010000110" => rgb <= "101000";
					when "00111011010000111" => rgb <= "101000";
					when "00111011010001000" => rgb <= "101000";
					when "00111011010001001" => rgb <= "101000";
					when "00111011010001010" => rgb <= "101000";
					when "00111011010001011" => rgb <= "101000";
					when "00111011010001100" => rgb <= "101000";
					when "00111011010001101" => rgb <= "101000";
					when "00111011010001110" => rgb <= "101000";
					when "00111011010001111" => rgb <= "101000";
					when "00111011010010000" => rgb <= "101000";
					when "00111011010010001" => rgb <= "101000";
					when "00111011010010010" => rgb <= "101000";
					when "00111011010010011" => rgb <= "101000";
					when "00111011010010100" => rgb <= "101000";
					when "00111011010010101" => rgb <= "101000";
					when "00111011010010110" => rgb <= "101000";
					when "00111011010010111" => rgb <= "101000";
					when "00111011010011000" => rgb <= "101000";
					when "00111011010011001" => rgb <= "101000";
					when "00111011010011010" => rgb <= "101000";
					when "00111011010011011" => rgb <= "101000";
					when "00111011010011100" => rgb <= "101000";
					when "00111011010011101" => rgb <= "101000";
					when "00111011010011110" => rgb <= "101000";
					when "00111011010011111" => rgb <= "101000";
					when "00111011010100000" => rgb <= "101000";
					when "00111011010100001" => rgb <= "101000";
					when "00111011010100010" => rgb <= "101000";
					when "00111011010100011" => rgb <= "101000";
					when "00111011010100100" => rgb <= "101000";
					when "00111011010100101" => rgb <= "101000";
					when "00111011010100110" => rgb <= "101000";
					when "00111011010100111" => rgb <= "101000";
					when "00111011010101000" => rgb <= "101000";
					when "00111011010101001" => rgb <= "101000";
					when "00111011010101010" => rgb <= "101000";
					when "00111011010101011" => rgb <= "101000";
					when "00111011010101100" => rgb <= "101000";
					when "00111011010101101" => rgb <= "101000";
					when "00111011010101110" => rgb <= "101000";
					when "00111011010101111" => rgb <= "101000";
					when "00111011010110000" => rgb <= "101000";
					when "00111011010110001" => rgb <= "101000";
					when "00111011010110010" => rgb <= "101000";
					when "00111011010110011" => rgb <= "101000";
					when "00111011010110100" => rgb <= "101000";
					when "00111011010110101" => rgb <= "101000";
					when "00111011010110110" => rgb <= "101000";
					when "00111011010110111" => rgb <= "101000";
					when "00111011010111000" => rgb <= "101000";
					when "00111011010111001" => rgb <= "101000";
					when "00111011010111010" => rgb <= "101000";
					when "00111011010111011" => rgb <= "101000";
					when "00111011010111100" => rgb <= "101000";
					when "00111011010111101" => rgb <= "101000";
					when "00111011010111110" => rgb <= "101000";
					when "00111011010111111" => rgb <= "101000";
					when "00111011011000000" => rgb <= "100100";
					when "00111011011000001" => rgb <= "000000";
					when "00111011011000010" => rgb <= "000000";
					when "00111011011000011" => rgb <= "000000";
					when "00111011011000100" => rgb <= "000000";
					when "00111011011000101" => rgb <= "000000";
					when "00111011011000110" => rgb <= "000000";
					when "00111011011000111" => rgb <= "000000";
					when "00111011011001000" => rgb <= "000000";
					when "00111011011001001" => rgb <= "000000";
					when "00111011011001010" => rgb <= "000000";
					when "00111011011001011" => rgb <= "000000";
					when "00111011011001100" => rgb <= "010100";
					when "00111011011001101" => rgb <= "101000";
					when "00111011011001110" => rgb <= "101000";
					when "00111011011001111" => rgb <= "101000";
					when "00111011011010000" => rgb <= "101000";
					when "00111011011010001" => rgb <= "101000";
					when "00111011011010010" => rgb <= "101000";
					when "00111011011010011" => rgb <= "101000";
					when "00111011011010100" => rgb <= "101000";
					when "00111011011010101" => rgb <= "101000";
					when "00111011011010110" => rgb <= "101000";
					when "00111011011010111" => rgb <= "010100";
					when "00111011011011000" => rgb <= "000000";
					when "00111011011011001" => rgb <= "000000";
					when "00111011011011010" => rgb <= "000000";
					when "00111011011011011" => rgb <= "000000";
					when "00111011011011100" => rgb <= "000000";
					when "00111011011011101" => rgb <= "000000";
					when "00111011011011110" => rgb <= "000000";
					when "00111011011011111" => rgb <= "000000";
					when "00111011011100000" => rgb <= "000000";
					when "00111011011100001" => rgb <= "000000";
					when "00111011011100010" => rgb <= "000000";
					when "00111011011100011" => rgb <= "000000";
					when "00111011011100100" => rgb <= "000000";
					when "00111011011100101" => rgb <= "000000";
					when "00111011011100110" => rgb <= "000000";
					when "00111011011100111" => rgb <= "000000";
					when "00111011011101000" => rgb <= "000000";
					when "00111011011101001" => rgb <= "000000";
					when "00111011011101010" => rgb <= "000000";
					when "00111011011101011" => rgb <= "000000";
					when "00111011011101100" => rgb <= "000000";
					when "00111011011101101" => rgb <= "000000";
					when "00111011011101110" => rgb <= "000000";
					when "00111011011101111" => rgb <= "000000";
					when "00111011011110000" => rgb <= "000000";
					when "00111011011110001" => rgb <= "000000";
					when "00111011011110010" => rgb <= "000000";
					when "00111011011110011" => rgb <= "000000";
					when "00111011011110100" => rgb <= "000000";
					when "00111011011110101" => rgb <= "000000";
					when "00111011011110110" => rgb <= "000000";
					when "00111011011110111" => rgb <= "000000";
					when "00111011011111000" => rgb <= "000000";
					when "00111011011111001" => rgb <= "000000";
					when "00111011011111010" => rgb <= "000000";
					when "00111011011111011" => rgb <= "000000";
					when "00111011011111100" => rgb <= "000000";
					when "00111011011111101" => rgb <= "000000";
					when "00111011011111110" => rgb <= "000000";
					when "00111011011111111" => rgb <= "000000";
					when "00111011100000000" => rgb <= "000000";
					when "00111011100000001" => rgb <= "000000";
					when "00111011100000010" => rgb <= "000000";
					when "00111011100000011" => rgb <= "000000";
					when "00111011100000100" => rgb <= "000000";
					when "00111011100000101" => rgb <= "000000";
					when "00111011100000110" => rgb <= "000000";
					when "00111011100000111" => rgb <= "000000";
					when "00111011100001000" => rgb <= "000000";
					when "00111011100001001" => rgb <= "000000";
					when "00111011100001010" => rgb <= "000000";
					when "00111011100001011" => rgb <= "000000";
					when "00111011100001100" => rgb <= "000000";
					when "00111011100001101" => rgb <= "000000";
					when "00111011100001110" => rgb <= "000000";
					when "00111011100001111" => rgb <= "000000";
					when "00111011100010000" => rgb <= "000000";
					when "00111011100010001" => rgb <= "000000";
					when "00111011100010010" => rgb <= "000000";
					when "00111011100010011" => rgb <= "000000";
					when "00111011100010100" => rgb <= "000000";
					when "00111011100010101" => rgb <= "000000";
					when "00111011100010110" => rgb <= "000000";
					when "00111011100010111" => rgb <= "000000";
					when "00111011100011000" => rgb <= "000000";
					when "00111011100011001" => rgb <= "000000";
					when "00111011100011010" => rgb <= "000000";
					when "00111011100011011" => rgb <= "000000";
					when "00111011100011100" => rgb <= "000000";
					when "00111011100011101" => rgb <= "000000";
					when "00111011100011110" => rgb <= "000000";
					when "00111011100011111" => rgb <= "000000";
					when "00111011100100000" => rgb <= "000000";
					when "00111011100100001" => rgb <= "000000";
					when "00111011100100010" => rgb <= "000000";
					when "00111011100100011" => rgb <= "000000";
					when "00111011100100100" => rgb <= "000000";
					when "00111011100100101" => rgb <= "000000";
					when "00111011100100110" => rgb <= "000000";
					when "00111011100100111" => rgb <= "000000";
					when "00111011100101000" => rgb <= "000000";
					when "00111011100101001" => rgb <= "000000";
					when "00111011100101010" => rgb <= "000000";
					when "00111011100101011" => rgb <= "000000";
					when "00111011100101100" => rgb <= "000000";
					when "00111011100101101" => rgb <= "000000";
					when "00111011100101110" => rgb <= "000000";
					when "00111011100101111" => rgb <= "000000";
					when "00111011100110000" => rgb <= "000000";
					when "00111011100110001" => rgb <= "000000";
					when "00111011100110010" => rgb <= "000000";
					when "00111011100110011" => rgb <= "000000";
					when "00111011100110100" => rgb <= "000000";
					when "00111011100110101" => rgb <= "000000";
					when "00111011100110110" => rgb <= "000000";
					when "00111011100110111" => rgb <= "000000";
					when "00111011100111000" => rgb <= "000000";
					when "00111011100111001" => rgb <= "000000";
					when "00111011100111010" => rgb <= "000000";
					when "00111011100111011" => rgb <= "000000";
					when "00111011100111100" => rgb <= "000000";
					when "00111011100111101" => rgb <= "000000";
					when "00111011100111110" => rgb <= "000000";
					when "00111011100111111" => rgb <= "000000";
					when "00111100000000000" => rgb <= "000000";
					when "00111100000000001" => rgb <= "000000";
					when "00111100000000010" => rgb <= "000000";
					when "00111100000000011" => rgb <= "000000";
					when "00111100000000100" => rgb <= "000000";
					when "00111100000000101" => rgb <= "000000";
					when "00111100000000110" => rgb <= "000000";
					when "00111100000000111" => rgb <= "000000";
					when "00111100000001000" => rgb <= "000000";
					when "00111100000001001" => rgb <= "000000";
					when "00111100000001010" => rgb <= "000000";
					when "00111100000001011" => rgb <= "000000";
					when "00111100000001100" => rgb <= "000000";
					when "00111100000001101" => rgb <= "000000";
					when "00111100000001110" => rgb <= "000000";
					when "00111100000001111" => rgb <= "000000";
					when "00111100000010000" => rgb <= "000000";
					when "00111100000010001" => rgb <= "000000";
					when "00111100000010010" => rgb <= "000000";
					when "00111100000010011" => rgb <= "000000";
					when "00111100000010100" => rgb <= "000000";
					when "00111100000010101" => rgb <= "000000";
					when "00111100000010110" => rgb <= "000000";
					when "00111100000010111" => rgb <= "000000";
					when "00111100000011000" => rgb <= "000000";
					when "00111100000011001" => rgb <= "000000";
					when "00111100000011010" => rgb <= "000000";
					when "00111100000011011" => rgb <= "000000";
					when "00111100000011100" => rgb <= "000000";
					when "00111100000011101" => rgb <= "000000";
					when "00111100000011110" => rgb <= "000000";
					when "00111100000011111" => rgb <= "000000";
					when "00111100000100000" => rgb <= "000000";
					when "00111100000100001" => rgb <= "000000";
					when "00111100000100010" => rgb <= "000000";
					when "00111100000100011" => rgb <= "000000";
					when "00111100000100100" => rgb <= "000000";
					when "00111100000100101" => rgb <= "000000";
					when "00111100000100110" => rgb <= "000000";
					when "00111100000100111" => rgb <= "000000";
					when "00111100000101000" => rgb <= "000000";
					when "00111100000101001" => rgb <= "000000";
					when "00111100000101010" => rgb <= "000000";
					when "00111100000101011" => rgb <= "000000";
					when "00111100000101100" => rgb <= "000000";
					when "00111100000101101" => rgb <= "000000";
					when "00111100000101110" => rgb <= "000000";
					when "00111100000101111" => rgb <= "000000";
					when "00111100000110000" => rgb <= "000000";
					when "00111100000110001" => rgb <= "000000";
					when "00111100000110010" => rgb <= "000000";
					when "00111100000110011" => rgb <= "000000";
					when "00111100000110100" => rgb <= "000000";
					when "00111100000110101" => rgb <= "000000";
					when "00111100000110110" => rgb <= "000000";
					when "00111100000110111" => rgb <= "000000";
					when "00111100000111000" => rgb <= "000000";
					when "00111100000111001" => rgb <= "000000";
					when "00111100000111010" => rgb <= "000000";
					when "00111100000111011" => rgb <= "000000";
					when "00111100000111100" => rgb <= "000000";
					when "00111100000111101" => rgb <= "000000";
					when "00111100000111110" => rgb <= "000000";
					when "00111100000111111" => rgb <= "000000";
					when "00111100001000000" => rgb <= "000000";
					when "00111100001000001" => rgb <= "000000";
					when "00111100001000010" => rgb <= "000000";
					when "00111100001000011" => rgb <= "000000";
					when "00111100001000100" => rgb <= "000000";
					when "00111100001000101" => rgb <= "000000";
					when "00111100001000110" => rgb <= "000000";
					when "00111100001000111" => rgb <= "000000";
					when "00111100001001000" => rgb <= "000000";
					when "00111100001001001" => rgb <= "000000";
					when "00111100001001010" => rgb <= "000000";
					when "00111100001001011" => rgb <= "000000";
					when "00111100001001100" => rgb <= "000000";
					when "00111100001001101" => rgb <= "000000";
					when "00111100001001110" => rgb <= "000000";
					when "00111100001001111" => rgb <= "000000";
					when "00111100001010000" => rgb <= "000000";
					when "00111100001010001" => rgb <= "000000";
					when "00111100001010010" => rgb <= "000000";
					when "00111100001010011" => rgb <= "000000";
					when "00111100001010100" => rgb <= "000000";
					when "00111100001010101" => rgb <= "000000";
					when "00111100001010110" => rgb <= "000000";
					when "00111100001010111" => rgb <= "000000";
					when "00111100001011000" => rgb <= "000000";
					when "00111100001011001" => rgb <= "000000";
					when "00111100001011010" => rgb <= "000000";
					when "00111100001011011" => rgb <= "000000";
					when "00111100001011100" => rgb <= "000000";
					when "00111100001011101" => rgb <= "000000";
					when "00111100001011110" => rgb <= "000000";
					when "00111100001011111" => rgb <= "000000";
					when "00111100001100000" => rgb <= "000000";
					when "00111100001100001" => rgb <= "000000";
					when "00111100001100010" => rgb <= "000000";
					when "00111100001100011" => rgb <= "000000";
					when "00111100001100100" => rgb <= "000000";
					when "00111100001100101" => rgb <= "000000";
					when "00111100001100110" => rgb <= "010100";
					when "00111100001100111" => rgb <= "111000";
					when "00111100001101000" => rgb <= "101000";
					when "00111100001101001" => rgb <= "101000";
					when "00111100001101010" => rgb <= "101000";
					when "00111100001101011" => rgb <= "101000";
					when "00111100001101100" => rgb <= "101000";
					when "00111100001101101" => rgb <= "101000";
					when "00111100001101110" => rgb <= "101000";
					when "00111100001101111" => rgb <= "101000";
					when "00111100001110000" => rgb <= "101000";
					when "00111100001110001" => rgb <= "100100";
					when "00111100001110010" => rgb <= "000000";
					when "00111100001110011" => rgb <= "000000";
					when "00111100001110100" => rgb <= "000000";
					when "00111100001110101" => rgb <= "000000";
					when "00111100001110110" => rgb <= "000000";
					when "00111100001110111" => rgb <= "000000";
					when "00111100001111000" => rgb <= "000000";
					when "00111100001111001" => rgb <= "000000";
					when "00111100001111010" => rgb <= "000000";
					when "00111100001111011" => rgb <= "000000";
					when "00111100001111100" => rgb <= "000000";
					when "00111100001111101" => rgb <= "101000";
					when "00111100001111110" => rgb <= "101000";
					when "00111100001111111" => rgb <= "101000";
					when "00111100010000000" => rgb <= "101000";
					when "00111100010000001" => rgb <= "101000";
					when "00111100010000010" => rgb <= "101000";
					when "00111100010000011" => rgb <= "101000";
					when "00111100010000100" => rgb <= "101000";
					when "00111100010000101" => rgb <= "101000";
					when "00111100010000110" => rgb <= "101000";
					when "00111100010000111" => rgb <= "101000";
					when "00111100010001000" => rgb <= "101000";
					when "00111100010001001" => rgb <= "101000";
					when "00111100010001010" => rgb <= "101000";
					when "00111100010001011" => rgb <= "101000";
					when "00111100010001100" => rgb <= "101000";
					when "00111100010001101" => rgb <= "101000";
					when "00111100010001110" => rgb <= "101000";
					when "00111100010001111" => rgb <= "101000";
					when "00111100010010000" => rgb <= "101000";
					when "00111100010010001" => rgb <= "101000";
					when "00111100010010010" => rgb <= "101000";
					when "00111100010010011" => rgb <= "101000";
					when "00111100010010100" => rgb <= "101000";
					when "00111100010010101" => rgb <= "101000";
					when "00111100010010110" => rgb <= "101000";
					when "00111100010010111" => rgb <= "101000";
					when "00111100010011000" => rgb <= "101000";
					when "00111100010011001" => rgb <= "101000";
					when "00111100010011010" => rgb <= "101000";
					when "00111100010011011" => rgb <= "101000";
					when "00111100010011100" => rgb <= "101000";
					when "00111100010011101" => rgb <= "101000";
					when "00111100010011110" => rgb <= "101000";
					when "00111100010011111" => rgb <= "101000";
					when "00111100010100000" => rgb <= "101000";
					when "00111100010100001" => rgb <= "101000";
					when "00111100010100010" => rgb <= "101000";
					when "00111100010100011" => rgb <= "101000";
					when "00111100010100100" => rgb <= "101000";
					when "00111100010100101" => rgb <= "101000";
					when "00111100010100110" => rgb <= "101000";
					when "00111100010100111" => rgb <= "101000";
					when "00111100010101000" => rgb <= "101000";
					when "00111100010101001" => rgb <= "101000";
					when "00111100010101010" => rgb <= "101000";
					when "00111100010101011" => rgb <= "101000";
					when "00111100010101100" => rgb <= "101000";
					when "00111100010101101" => rgb <= "101000";
					when "00111100010101110" => rgb <= "101000";
					when "00111100010101111" => rgb <= "101000";
					when "00111100010110000" => rgb <= "101000";
					when "00111100010110001" => rgb <= "101000";
					when "00111100010110010" => rgb <= "101000";
					when "00111100010110011" => rgb <= "101000";
					when "00111100010110100" => rgb <= "101000";
					when "00111100010110101" => rgb <= "101000";
					when "00111100010110110" => rgb <= "101000";
					when "00111100010110111" => rgb <= "101000";
					when "00111100010111000" => rgb <= "101000";
					when "00111100010111001" => rgb <= "101000";
					when "00111100010111010" => rgb <= "101000";
					when "00111100010111011" => rgb <= "101000";
					when "00111100010111100" => rgb <= "101000";
					when "00111100010111101" => rgb <= "101000";
					when "00111100010111110" => rgb <= "101000";
					when "00111100010111111" => rgb <= "101000";
					when "00111100011000000" => rgb <= "101000";
					when "00111100011000001" => rgb <= "000000";
					when "00111100011000010" => rgb <= "000000";
					when "00111100011000011" => rgb <= "000000";
					when "00111100011000100" => rgb <= "000000";
					when "00111100011000101" => rgb <= "000000";
					when "00111100011000110" => rgb <= "000000";
					when "00111100011000111" => rgb <= "000000";
					when "00111100011001000" => rgb <= "000000";
					when "00111100011001001" => rgb <= "000000";
					when "00111100011001010" => rgb <= "000000";
					when "00111100011001011" => rgb <= "000000";
					when "00111100011001100" => rgb <= "100100";
					when "00111100011001101" => rgb <= "101000";
					when "00111100011001110" => rgb <= "101000";
					when "00111100011001111" => rgb <= "101000";
					when "00111100011010000" => rgb <= "101000";
					when "00111100011010001" => rgb <= "101000";
					when "00111100011010010" => rgb <= "101000";
					when "00111100011010011" => rgb <= "101000";
					when "00111100011010100" => rgb <= "101000";
					when "00111100011010101" => rgb <= "101000";
					when "00111100011010110" => rgb <= "101000";
					when "00111100011010111" => rgb <= "010100";
					when "00111100011011000" => rgb <= "000000";
					when "00111100011011001" => rgb <= "000000";
					when "00111100011011010" => rgb <= "000000";
					when "00111100011011011" => rgb <= "000000";
					when "00111100011011100" => rgb <= "000000";
					when "00111100011011101" => rgb <= "000000";
					when "00111100011011110" => rgb <= "000000";
					when "00111100011011111" => rgb <= "000000";
					when "00111100011100000" => rgb <= "000000";
					when "00111100011100001" => rgb <= "000000";
					when "00111100011100010" => rgb <= "000000";
					when "00111100011100011" => rgb <= "000000";
					when "00111100011100100" => rgb <= "000000";
					when "00111100011100101" => rgb <= "000000";
					when "00111100011100110" => rgb <= "000000";
					when "00111100011100111" => rgb <= "000000";
					when "00111100011101000" => rgb <= "000000";
					when "00111100011101001" => rgb <= "000000";
					when "00111100011101010" => rgb <= "000000";
					when "00111100011101011" => rgb <= "000000";
					when "00111100011101100" => rgb <= "000000";
					when "00111100011101101" => rgb <= "000000";
					when "00111100011101110" => rgb <= "000000";
					when "00111100011101111" => rgb <= "000000";
					when "00111100011110000" => rgb <= "000000";
					when "00111100011110001" => rgb <= "000000";
					when "00111100011110010" => rgb <= "000000";
					when "00111100011110011" => rgb <= "000000";
					when "00111100011110100" => rgb <= "000000";
					when "00111100011110101" => rgb <= "000000";
					when "00111100011110110" => rgb <= "000000";
					when "00111100011110111" => rgb <= "000000";
					when "00111100011111000" => rgb <= "000000";
					when "00111100011111001" => rgb <= "000000";
					when "00111100011111010" => rgb <= "000000";
					when "00111100011111011" => rgb <= "000000";
					when "00111100011111100" => rgb <= "000000";
					when "00111100011111101" => rgb <= "000000";
					when "00111100011111110" => rgb <= "000000";
					when "00111100011111111" => rgb <= "000000";
					when "00111100100000000" => rgb <= "000000";
					when "00111100100000001" => rgb <= "000000";
					when "00111100100000010" => rgb <= "000000";
					when "00111100100000011" => rgb <= "000000";
					when "00111100100000100" => rgb <= "000000";
					when "00111100100000101" => rgb <= "000000";
					when "00111100100000110" => rgb <= "000000";
					when "00111100100000111" => rgb <= "000000";
					when "00111100100001000" => rgb <= "000000";
					when "00111100100001001" => rgb <= "000000";
					when "00111100100001010" => rgb <= "000000";
					when "00111100100001011" => rgb <= "000000";
					when "00111100100001100" => rgb <= "000000";
					when "00111100100001101" => rgb <= "000000";
					when "00111100100001110" => rgb <= "000000";
					when "00111100100001111" => rgb <= "000000";
					when "00111100100010000" => rgb <= "000000";
					when "00111100100010001" => rgb <= "000000";
					when "00111100100010010" => rgb <= "000000";
					when "00111100100010011" => rgb <= "000000";
					when "00111100100010100" => rgb <= "000000";
					when "00111100100010101" => rgb <= "000000";
					when "00111100100010110" => rgb <= "000000";
					when "00111100100010111" => rgb <= "000000";
					when "00111100100011000" => rgb <= "000000";
					when "00111100100011001" => rgb <= "000000";
					when "00111100100011010" => rgb <= "000000";
					when "00111100100011011" => rgb <= "000000";
					when "00111100100011100" => rgb <= "000000";
					when "00111100100011101" => rgb <= "000000";
					when "00111100100011110" => rgb <= "000000";
					when "00111100100011111" => rgb <= "000000";
					when "00111100100100000" => rgb <= "000000";
					when "00111100100100001" => rgb <= "000000";
					when "00111100100100010" => rgb <= "000000";
					when "00111100100100011" => rgb <= "000000";
					when "00111100100100100" => rgb <= "000000";
					when "00111100100100101" => rgb <= "000000";
					when "00111100100100110" => rgb <= "000000";
					when "00111100100100111" => rgb <= "000000";
					when "00111100100101000" => rgb <= "000000";
					when "00111100100101001" => rgb <= "000000";
					when "00111100100101010" => rgb <= "000000";
					when "00111100100101011" => rgb <= "000000";
					when "00111100100101100" => rgb <= "000000";
					when "00111100100101101" => rgb <= "000000";
					when "00111100100101110" => rgb <= "000000";
					when "00111100100101111" => rgb <= "000000";
					when "00111100100110000" => rgb <= "000000";
					when "00111100100110001" => rgb <= "000000";
					when "00111100100110010" => rgb <= "000000";
					when "00111100100110011" => rgb <= "000000";
					when "00111100100110100" => rgb <= "000000";
					when "00111100100110101" => rgb <= "000000";
					when "00111100100110110" => rgb <= "000000";
					when "00111100100110111" => rgb <= "000000";
					when "00111100100111000" => rgb <= "000000";
					when "00111100100111001" => rgb <= "000000";
					when "00111100100111010" => rgb <= "000000";
					when "00111100100111011" => rgb <= "000000";
					when "00111100100111100" => rgb <= "000000";
					when "00111100100111101" => rgb <= "000000";
					when "00111100100111110" => rgb <= "000000";
					when "00111100100111111" => rgb <= "000000";
					when "00111101000000000" => rgb <= "000000";
					when "00111101000000001" => rgb <= "000000";
					when "00111101000000010" => rgb <= "000000";
					when "00111101000000011" => rgb <= "000000";
					when "00111101000000100" => rgb <= "000000";
					when "00111101000000101" => rgb <= "000000";
					when "00111101000000110" => rgb <= "000000";
					when "00111101000000111" => rgb <= "000000";
					when "00111101000001000" => rgb <= "000000";
					when "00111101000001001" => rgb <= "000000";
					when "00111101000001010" => rgb <= "000000";
					when "00111101000001011" => rgb <= "000000";
					when "00111101000001100" => rgb <= "000000";
					when "00111101000001101" => rgb <= "000000";
					when "00111101000001110" => rgb <= "000000";
					when "00111101000001111" => rgb <= "000000";
					when "00111101000010000" => rgb <= "000000";
					when "00111101000010001" => rgb <= "000000";
					when "00111101000010010" => rgb <= "000000";
					when "00111101000010011" => rgb <= "000000";
					when "00111101000010100" => rgb <= "000000";
					when "00111101000010101" => rgb <= "000000";
					when "00111101000010110" => rgb <= "000000";
					when "00111101000010111" => rgb <= "000000";
					when "00111101000011000" => rgb <= "000000";
					when "00111101000011001" => rgb <= "000000";
					when "00111101000011010" => rgb <= "000000";
					when "00111101000011011" => rgb <= "000000";
					when "00111101000011100" => rgb <= "000000";
					when "00111101000011101" => rgb <= "000000";
					when "00111101000011110" => rgb <= "000000";
					when "00111101000011111" => rgb <= "000000";
					when "00111101000100000" => rgb <= "000000";
					when "00111101000100001" => rgb <= "000000";
					when "00111101000100010" => rgb <= "000000";
					when "00111101000100011" => rgb <= "000000";
					when "00111101000100100" => rgb <= "000000";
					when "00111101000100101" => rgb <= "000000";
					when "00111101000100110" => rgb <= "000000";
					when "00111101000100111" => rgb <= "000000";
					when "00111101000101000" => rgb <= "000000";
					when "00111101000101001" => rgb <= "000000";
					when "00111101000101010" => rgb <= "000000";
					when "00111101000101011" => rgb <= "000000";
					when "00111101000101100" => rgb <= "000000";
					when "00111101000101101" => rgb <= "000000";
					when "00111101000101110" => rgb <= "000000";
					when "00111101000101111" => rgb <= "000000";
					when "00111101000110000" => rgb <= "000000";
					when "00111101000110001" => rgb <= "000000";
					when "00111101000110010" => rgb <= "000000";
					when "00111101000110011" => rgb <= "000000";
					when "00111101000110100" => rgb <= "000000";
					when "00111101000110101" => rgb <= "000000";
					when "00111101000110110" => rgb <= "000000";
					when "00111101000110111" => rgb <= "000000";
					when "00111101000111000" => rgb <= "000000";
					when "00111101000111001" => rgb <= "000000";
					when "00111101000111010" => rgb <= "000000";
					when "00111101000111011" => rgb <= "000000";
					when "00111101000111100" => rgb <= "000000";
					when "00111101000111101" => rgb <= "000000";
					when "00111101000111110" => rgb <= "000000";
					when "00111101000111111" => rgb <= "000000";
					when "00111101001000000" => rgb <= "000000";
					when "00111101001000001" => rgb <= "000000";
					when "00111101001000010" => rgb <= "000000";
					when "00111101001000011" => rgb <= "000000";
					when "00111101001000100" => rgb <= "000000";
					when "00111101001000101" => rgb <= "000000";
					when "00111101001000110" => rgb <= "000000";
					when "00111101001000111" => rgb <= "000000";
					when "00111101001001000" => rgb <= "000000";
					when "00111101001001001" => rgb <= "000000";
					when "00111101001001010" => rgb <= "000000";
					when "00111101001001011" => rgb <= "000000";
					when "00111101001001100" => rgb <= "000000";
					when "00111101001001101" => rgb <= "000000";
					when "00111101001001110" => rgb <= "000000";
					when "00111101001001111" => rgb <= "000000";
					when "00111101001010000" => rgb <= "000000";
					when "00111101001010001" => rgb <= "000000";
					when "00111101001010010" => rgb <= "000000";
					when "00111101001010011" => rgb <= "000000";
					when "00111101001010100" => rgb <= "000000";
					when "00111101001010101" => rgb <= "000000";
					when "00111101001010110" => rgb <= "000000";
					when "00111101001010111" => rgb <= "000000";
					when "00111101001011000" => rgb <= "000000";
					when "00111101001011001" => rgb <= "000000";
					when "00111101001011010" => rgb <= "000000";
					when "00111101001011011" => rgb <= "000000";
					when "00111101001011100" => rgb <= "000000";
					when "00111101001011101" => rgb <= "000000";
					when "00111101001011110" => rgb <= "000000";
					when "00111101001011111" => rgb <= "000000";
					when "00111101001100000" => rgb <= "000000";
					when "00111101001100001" => rgb <= "000000";
					when "00111101001100010" => rgb <= "000000";
					when "00111101001100011" => rgb <= "000000";
					when "00111101001100100" => rgb <= "000000";
					when "00111101001100101" => rgb <= "000000";
					when "00111101001100110" => rgb <= "010100";
					when "00111101001100111" => rgb <= "101000";
					when "00111101001101000" => rgb <= "111000";
					when "00111101001101001" => rgb <= "111000";
					when "00111101001101010" => rgb <= "111000";
					when "00111101001101011" => rgb <= "111000";
					when "00111101001101100" => rgb <= "111000";
					when "00111101001101101" => rgb <= "111000";
					when "00111101001101110" => rgb <= "111000";
					when "00111101001101111" => rgb <= "111000";
					when "00111101001110000" => rgb <= "111000";
					when "00111101001110001" => rgb <= "101000";
					when "00111101001110010" => rgb <= "000000";
					when "00111101001110011" => rgb <= "000000";
					when "00111101001110100" => rgb <= "000000";
					when "00111101001110101" => rgb <= "000000";
					when "00111101001110110" => rgb <= "000000";
					when "00111101001110111" => rgb <= "000000";
					when "00111101001111000" => rgb <= "000000";
					when "00111101001111001" => rgb <= "000000";
					when "00111101001111010" => rgb <= "000000";
					when "00111101001111011" => rgb <= "000000";
					when "00111101001111100" => rgb <= "000000";
					when "00111101001111101" => rgb <= "101000";
					when "00111101001111110" => rgb <= "101000";
					when "00111101001111111" => rgb <= "101000";
					when "00111101010000000" => rgb <= "101000";
					when "00111101010000001" => rgb <= "101000";
					when "00111101010000010" => rgb <= "101000";
					when "00111101010000011" => rgb <= "101000";
					when "00111101010000100" => rgb <= "101000";
					when "00111101010000101" => rgb <= "101000";
					when "00111101010000110" => rgb <= "101000";
					when "00111101010000111" => rgb <= "101000";
					when "00111101010001000" => rgb <= "101000";
					when "00111101010001001" => rgb <= "101000";
					when "00111101010001010" => rgb <= "101000";
					when "00111101010001011" => rgb <= "101000";
					when "00111101010001100" => rgb <= "101000";
					when "00111101010001101" => rgb <= "101000";
					when "00111101010001110" => rgb <= "101000";
					when "00111101010001111" => rgb <= "101000";
					when "00111101010010000" => rgb <= "101000";
					when "00111101010010001" => rgb <= "101000";
					when "00111101010010010" => rgb <= "101000";
					when "00111101010010011" => rgb <= "101000";
					when "00111101010010100" => rgb <= "101000";
					when "00111101010010101" => rgb <= "101000";
					when "00111101010010110" => rgb <= "101000";
					when "00111101010010111" => rgb <= "101000";
					when "00111101010011000" => rgb <= "101000";
					when "00111101010011001" => rgb <= "101000";
					when "00111101010011010" => rgb <= "101000";
					when "00111101010011011" => rgb <= "101000";
					when "00111101010011100" => rgb <= "101000";
					when "00111101010011101" => rgb <= "101000";
					when "00111101010011110" => rgb <= "101000";
					when "00111101010011111" => rgb <= "101000";
					when "00111101010100000" => rgb <= "101000";
					when "00111101010100001" => rgb <= "101000";
					when "00111101010100010" => rgb <= "101000";
					when "00111101010100011" => rgb <= "101000";
					when "00111101010100100" => rgb <= "101000";
					when "00111101010100101" => rgb <= "101000";
					when "00111101010100110" => rgb <= "101000";
					when "00111101010100111" => rgb <= "101000";
					when "00111101010101000" => rgb <= "101000";
					when "00111101010101001" => rgb <= "101000";
					when "00111101010101010" => rgb <= "101000";
					when "00111101010101011" => rgb <= "101000";
					when "00111101010101100" => rgb <= "101000";
					when "00111101010101101" => rgb <= "101000";
					when "00111101010101110" => rgb <= "101000";
					when "00111101010101111" => rgb <= "101000";
					when "00111101010110000" => rgb <= "101000";
					when "00111101010110001" => rgb <= "101000";
					when "00111101010110010" => rgb <= "101000";
					when "00111101010110011" => rgb <= "101000";
					when "00111101010110100" => rgb <= "101000";
					when "00111101010110101" => rgb <= "101000";
					when "00111101010110110" => rgb <= "101000";
					when "00111101010110111" => rgb <= "101000";
					when "00111101010111000" => rgb <= "101000";
					when "00111101010111001" => rgb <= "101000";
					when "00111101010111010" => rgb <= "101000";
					when "00111101010111011" => rgb <= "101000";
					when "00111101010111100" => rgb <= "101000";
					when "00111101010111101" => rgb <= "101000";
					when "00111101010111110" => rgb <= "101000";
					when "00111101010111111" => rgb <= "101000";
					when "00111101011000000" => rgb <= "100100";
					when "00111101011000001" => rgb <= "000000";
					when "00111101011000010" => rgb <= "000000";
					when "00111101011000011" => rgb <= "000000";
					when "00111101011000100" => rgb <= "000000";
					when "00111101011000101" => rgb <= "000000";
					when "00111101011000110" => rgb <= "000000";
					when "00111101011000111" => rgb <= "000000";
					when "00111101011001000" => rgb <= "000000";
					when "00111101011001001" => rgb <= "000000";
					when "00111101011001010" => rgb <= "000000";
					when "00111101011001011" => rgb <= "000000";
					when "00111101011001100" => rgb <= "100100";
					when "00111101011001101" => rgb <= "101000";
					when "00111101011001110" => rgb <= "101000";
					when "00111101011001111" => rgb <= "101000";
					when "00111101011010000" => rgb <= "101000";
					when "00111101011010001" => rgb <= "101000";
					when "00111101011010010" => rgb <= "101000";
					when "00111101011010011" => rgb <= "101000";
					when "00111101011010100" => rgb <= "101000";
					when "00111101011010101" => rgb <= "101000";
					when "00111101011010110" => rgb <= "101000";
					when "00111101011010111" => rgb <= "010100";
					when "00111101011011000" => rgb <= "000000";
					when "00111101011011001" => rgb <= "000000";
					when "00111101011011010" => rgb <= "000000";
					when "00111101011011011" => rgb <= "000000";
					when "00111101011011100" => rgb <= "000000";
					when "00111101011011101" => rgb <= "000000";
					when "00111101011011110" => rgb <= "000000";
					when "00111101011011111" => rgb <= "000000";
					when "00111101011100000" => rgb <= "000000";
					when "00111101011100001" => rgb <= "000000";
					when "00111101011100010" => rgb <= "000000";
					when "00111101011100011" => rgb <= "000000";
					when "00111101011100100" => rgb <= "000000";
					when "00111101011100101" => rgb <= "000000";
					when "00111101011100110" => rgb <= "000000";
					when "00111101011100111" => rgb <= "000000";
					when "00111101011101000" => rgb <= "000000";
					when "00111101011101001" => rgb <= "000000";
					when "00111101011101010" => rgb <= "000000";
					when "00111101011101011" => rgb <= "000000";
					when "00111101011101100" => rgb <= "000000";
					when "00111101011101101" => rgb <= "000000";
					when "00111101011101110" => rgb <= "000000";
					when "00111101011101111" => rgb <= "000000";
					when "00111101011110000" => rgb <= "000000";
					when "00111101011110001" => rgb <= "000000";
					when "00111101011110010" => rgb <= "000000";
					when "00111101011110011" => rgb <= "000000";
					when "00111101011110100" => rgb <= "000000";
					when "00111101011110101" => rgb <= "000000";
					when "00111101011110110" => rgb <= "000000";
					when "00111101011110111" => rgb <= "000000";
					when "00111101011111000" => rgb <= "000000";
					when "00111101011111001" => rgb <= "000000";
					when "00111101011111010" => rgb <= "000000";
					when "00111101011111011" => rgb <= "000000";
					when "00111101011111100" => rgb <= "000000";
					when "00111101011111101" => rgb <= "000000";
					when "00111101011111110" => rgb <= "000000";
					when "00111101011111111" => rgb <= "000000";
					when "00111101100000000" => rgb <= "000000";
					when "00111101100000001" => rgb <= "000000";
					when "00111101100000010" => rgb <= "000000";
					when "00111101100000011" => rgb <= "000000";
					when "00111101100000100" => rgb <= "000000";
					when "00111101100000101" => rgb <= "000000";
					when "00111101100000110" => rgb <= "000000";
					when "00111101100000111" => rgb <= "000000";
					when "00111101100001000" => rgb <= "000000";
					when "00111101100001001" => rgb <= "000000";
					when "00111101100001010" => rgb <= "000000";
					when "00111101100001011" => rgb <= "000000";
					when "00111101100001100" => rgb <= "000000";
					when "00111101100001101" => rgb <= "000000";
					when "00111101100001110" => rgb <= "000000";
					when "00111101100001111" => rgb <= "000000";
					when "00111101100010000" => rgb <= "000000";
					when "00111101100010001" => rgb <= "000000";
					when "00111101100010010" => rgb <= "000000";
					when "00111101100010011" => rgb <= "000000";
					when "00111101100010100" => rgb <= "000000";
					when "00111101100010101" => rgb <= "000000";
					when "00111101100010110" => rgb <= "000000";
					when "00111101100010111" => rgb <= "000000";
					when "00111101100011000" => rgb <= "000000";
					when "00111101100011001" => rgb <= "000000";
					when "00111101100011010" => rgb <= "000000";
					when "00111101100011011" => rgb <= "000000";
					when "00111101100011100" => rgb <= "000000";
					when "00111101100011101" => rgb <= "000000";
					when "00111101100011110" => rgb <= "000000";
					when "00111101100011111" => rgb <= "000000";
					when "00111101100100000" => rgb <= "000000";
					when "00111101100100001" => rgb <= "000000";
					when "00111101100100010" => rgb <= "000000";
					when "00111101100100011" => rgb <= "000000";
					when "00111101100100100" => rgb <= "000000";
					when "00111101100100101" => rgb <= "000000";
					when "00111101100100110" => rgb <= "000000";
					when "00111101100100111" => rgb <= "000000";
					when "00111101100101000" => rgb <= "000000";
					when "00111101100101001" => rgb <= "000000";
					when "00111101100101010" => rgb <= "000000";
					when "00111101100101011" => rgb <= "000000";
					when "00111101100101100" => rgb <= "000000";
					when "00111101100101101" => rgb <= "000000";
					when "00111101100101110" => rgb <= "000000";
					when "00111101100101111" => rgb <= "000000";
					when "00111101100110000" => rgb <= "000000";
					when "00111101100110001" => rgb <= "000000";
					when "00111101100110010" => rgb <= "000000";
					when "00111101100110011" => rgb <= "000000";
					when "00111101100110100" => rgb <= "000000";
					when "00111101100110101" => rgb <= "000000";
					when "00111101100110110" => rgb <= "000000";
					when "00111101100110111" => rgb <= "000000";
					when "00111101100111000" => rgb <= "000000";
					when "00111101100111001" => rgb <= "000000";
					when "00111101100111010" => rgb <= "000000";
					when "00111101100111011" => rgb <= "000000";
					when "00111101100111100" => rgb <= "000000";
					when "00111101100111101" => rgb <= "000000";
					when "00111101100111110" => rgb <= "000000";
					when "00111101100111111" => rgb <= "000000";
					when "00111110000000000" => rgb <= "000000";
					when "00111110000000001" => rgb <= "000000";
					when "00111110000000010" => rgb <= "000000";
					when "00111110000000011" => rgb <= "000000";
					when "00111110000000100" => rgb <= "000000";
					when "00111110000000101" => rgb <= "000000";
					when "00111110000000110" => rgb <= "000000";
					when "00111110000000111" => rgb <= "000000";
					when "00111110000001000" => rgb <= "000000";
					when "00111110000001001" => rgb <= "000000";
					when "00111110000001010" => rgb <= "000000";
					when "00111110000001011" => rgb <= "000000";
					when "00111110000001100" => rgb <= "000000";
					when "00111110000001101" => rgb <= "000000";
					when "00111110000001110" => rgb <= "000000";
					when "00111110000001111" => rgb <= "000000";
					when "00111110000010000" => rgb <= "000000";
					when "00111110000010001" => rgb <= "000000";
					when "00111110000010010" => rgb <= "000000";
					when "00111110000010011" => rgb <= "000000";
					when "00111110000010100" => rgb <= "000000";
					when "00111110000010101" => rgb <= "000000";
					when "00111110000010110" => rgb <= "000000";
					when "00111110000010111" => rgb <= "000000";
					when "00111110000011000" => rgb <= "000000";
					when "00111110000011001" => rgb <= "000000";
					when "00111110000011010" => rgb <= "000000";
					when "00111110000011011" => rgb <= "000000";
					when "00111110000011100" => rgb <= "000000";
					when "00111110000011101" => rgb <= "000000";
					when "00111110000011110" => rgb <= "000000";
					when "00111110000011111" => rgb <= "000000";
					when "00111110000100000" => rgb <= "000000";
					when "00111110000100001" => rgb <= "000000";
					when "00111110000100010" => rgb <= "000000";
					when "00111110000100011" => rgb <= "000000";
					when "00111110000100100" => rgb <= "000000";
					when "00111110000100101" => rgb <= "000000";
					when "00111110000100110" => rgb <= "000000";
					when "00111110000100111" => rgb <= "000000";
					when "00111110000101000" => rgb <= "000000";
					when "00111110000101001" => rgb <= "000000";
					when "00111110000101010" => rgb <= "000000";
					when "00111110000101011" => rgb <= "000000";
					when "00111110000101100" => rgb <= "000000";
					when "00111110000101101" => rgb <= "000000";
					when "00111110000101110" => rgb <= "000000";
					when "00111110000101111" => rgb <= "000000";
					when "00111110000110000" => rgb <= "000000";
					when "00111110000110001" => rgb <= "000000";
					when "00111110000110010" => rgb <= "000000";
					when "00111110000110011" => rgb <= "000000";
					when "00111110000110100" => rgb <= "000000";
					when "00111110000110101" => rgb <= "000000";
					when "00111110000110110" => rgb <= "000000";
					when "00111110000110111" => rgb <= "000000";
					when "00111110000111000" => rgb <= "000000";
					when "00111110000111001" => rgb <= "000000";
					when "00111110000111010" => rgb <= "000000";
					when "00111110000111011" => rgb <= "000000";
					when "00111110000111100" => rgb <= "000000";
					when "00111110000111101" => rgb <= "000000";
					when "00111110000111110" => rgb <= "000000";
					when "00111110000111111" => rgb <= "000000";
					when "00111110001000000" => rgb <= "000000";
					when "00111110001000001" => rgb <= "000000";
					when "00111110001000010" => rgb <= "000000";
					when "00111110001000011" => rgb <= "000000";
					when "00111110001000100" => rgb <= "000000";
					when "00111110001000101" => rgb <= "000000";
					when "00111110001000110" => rgb <= "000000";
					when "00111110001000111" => rgb <= "000000";
					when "00111110001001000" => rgb <= "000000";
					when "00111110001001001" => rgb <= "000000";
					when "00111110001001010" => rgb <= "000000";
					when "00111110001001011" => rgb <= "000000";
					when "00111110001001100" => rgb <= "000000";
					when "00111110001001101" => rgb <= "000000";
					when "00111110001001110" => rgb <= "000000";
					when "00111110001001111" => rgb <= "000000";
					when "00111110001010000" => rgb <= "000000";
					when "00111110001010001" => rgb <= "000000";
					when "00111110001010010" => rgb <= "000000";
					when "00111110001010011" => rgb <= "000000";
					when "00111110001010100" => rgb <= "000000";
					when "00111110001010101" => rgb <= "000000";
					when "00111110001010110" => rgb <= "000000";
					when "00111110001010111" => rgb <= "000000";
					when "00111110001011000" => rgb <= "000000";
					when "00111110001011001" => rgb <= "000000";
					when "00111110001011010" => rgb <= "000000";
					when "00111110001011011" => rgb <= "000000";
					when "00111110001011100" => rgb <= "000000";
					when "00111110001011101" => rgb <= "000000";
					when "00111110001011110" => rgb <= "000000";
					when "00111110001011111" => rgb <= "000000";
					when "00111110001100000" => rgb <= "000000";
					when "00111110001100001" => rgb <= "000000";
					when "00111110001100010" => rgb <= "000000";
					when "00111110001100011" => rgb <= "000000";
					when "00111110001100100" => rgb <= "000000";
					when "00111110001100101" => rgb <= "000000";
					when "00111110001100110" => rgb <= "000000";
					when "00111110001100111" => rgb <= "010100";
					when "00111110001101000" => rgb <= "010100";
					when "00111110001101001" => rgb <= "010100";
					when "00111110001101010" => rgb <= "010100";
					when "00111110001101011" => rgb <= "010100";
					when "00111110001101100" => rgb <= "010100";
					when "00111110001101101" => rgb <= "010100";
					when "00111110001101110" => rgb <= "010100";
					when "00111110001101111" => rgb <= "010100";
					when "00111110001110000" => rgb <= "010100";
					when "00111110001110001" => rgb <= "010100";
					when "00111110001110010" => rgb <= "010100";
					when "00111110001110011" => rgb <= "010100";
					when "00111110001110100" => rgb <= "010100";
					when "00111110001110101" => rgb <= "010100";
					when "00111110001110110" => rgb <= "010100";
					when "00111110001110111" => rgb <= "010100";
					when "00111110001111000" => rgb <= "010100";
					when "00111110001111001" => rgb <= "010100";
					when "00111110001111010" => rgb <= "010100";
					when "00111110001111011" => rgb <= "010100";
					when "00111110001111100" => rgb <= "010100";
					when "00111110001111101" => rgb <= "101000";
					when "00111110001111110" => rgb <= "101000";
					when "00111110001111111" => rgb <= "101000";
					when "00111110010000000" => rgb <= "101000";
					when "00111110010000001" => rgb <= "101000";
					when "00111110010000010" => rgb <= "101000";
					when "00111110010000011" => rgb <= "101000";
					when "00111110010000100" => rgb <= "101000";
					when "00111110010000101" => rgb <= "101000";
					when "00111110010000110" => rgb <= "101000";
					when "00111110010000111" => rgb <= "101000";
					when "00111110010001000" => rgb <= "101000";
					when "00111110010001001" => rgb <= "101000";
					when "00111110010001010" => rgb <= "101000";
					when "00111110010001011" => rgb <= "101000";
					when "00111110010001100" => rgb <= "101000";
					when "00111110010001101" => rgb <= "101000";
					when "00111110010001110" => rgb <= "101000";
					when "00111110010001111" => rgb <= "101000";
					when "00111110010010000" => rgb <= "101000";
					when "00111110010010001" => rgb <= "101000";
					when "00111110010010010" => rgb <= "101000";
					when "00111110010010011" => rgb <= "101000";
					when "00111110010010100" => rgb <= "101000";
					when "00111110010010101" => rgb <= "101000";
					when "00111110010010110" => rgb <= "101000";
					when "00111110010010111" => rgb <= "101000";
					when "00111110010011000" => rgb <= "101000";
					when "00111110010011001" => rgb <= "101000";
					when "00111110010011010" => rgb <= "101000";
					when "00111110010011011" => rgb <= "101000";
					when "00111110010011100" => rgb <= "101000";
					when "00111110010011101" => rgb <= "101000";
					when "00111110010011110" => rgb <= "101000";
					when "00111110010011111" => rgb <= "101000";
					when "00111110010100000" => rgb <= "101000";
					when "00111110010100001" => rgb <= "101000";
					when "00111110010100010" => rgb <= "101000";
					when "00111110010100011" => rgb <= "101000";
					when "00111110010100100" => rgb <= "101000";
					when "00111110010100101" => rgb <= "101000";
					when "00111110010100110" => rgb <= "101000";
					when "00111110010100111" => rgb <= "101000";
					when "00111110010101000" => rgb <= "101000";
					when "00111110010101001" => rgb <= "101000";
					when "00111110010101010" => rgb <= "101000";
					when "00111110010101011" => rgb <= "101000";
					when "00111110010101100" => rgb <= "101000";
					when "00111110010101101" => rgb <= "101000";
					when "00111110010101110" => rgb <= "101000";
					when "00111110010101111" => rgb <= "101000";
					when "00111110010110000" => rgb <= "101000";
					when "00111110010110001" => rgb <= "101000";
					when "00111110010110010" => rgb <= "101000";
					when "00111110010110011" => rgb <= "101000";
					when "00111110010110100" => rgb <= "101000";
					when "00111110010110101" => rgb <= "101000";
					when "00111110010110110" => rgb <= "101000";
					when "00111110010110111" => rgb <= "101000";
					when "00111110010111000" => rgb <= "101000";
					when "00111110010111001" => rgb <= "101000";
					when "00111110010111010" => rgb <= "101000";
					when "00111110010111011" => rgb <= "101000";
					when "00111110010111100" => rgb <= "101000";
					when "00111110010111101" => rgb <= "101000";
					when "00111110010111110" => rgb <= "101000";
					when "00111110010111111" => rgb <= "101000";
					when "00111110011000000" => rgb <= "101000";
					when "00111110011000001" => rgb <= "010100";
					when "00111110011000010" => rgb <= "010100";
					when "00111110011000011" => rgb <= "010100";
					when "00111110011000100" => rgb <= "010100";
					when "00111110011000101" => rgb <= "010100";
					when "00111110011000110" => rgb <= "010100";
					when "00111110011000111" => rgb <= "010100";
					when "00111110011001000" => rgb <= "010100";
					when "00111110011001001" => rgb <= "010100";
					when "00111110011001010" => rgb <= "010100";
					when "00111110011001011" => rgb <= "010100";
					when "00111110011001100" => rgb <= "010100";
					when "00111110011001101" => rgb <= "010100";
					when "00111110011001110" => rgb <= "010100";
					when "00111110011001111" => rgb <= "010100";
					when "00111110011010000" => rgb <= "010100";
					when "00111110011010001" => rgb <= "010100";
					when "00111110011010010" => rgb <= "010100";
					when "00111110011010011" => rgb <= "010100";
					when "00111110011010100" => rgb <= "010100";
					when "00111110011010101" => rgb <= "010100";
					when "00111110011010110" => rgb <= "010100";
					when "00111110011010111" => rgb <= "000000";
					when "00111110011011000" => rgb <= "000000";
					when "00111110011011001" => rgb <= "000000";
					when "00111110011011010" => rgb <= "000000";
					when "00111110011011011" => rgb <= "000000";
					when "00111110011011100" => rgb <= "000000";
					when "00111110011011101" => rgb <= "000000";
					when "00111110011011110" => rgb <= "000000";
					when "00111110011011111" => rgb <= "000000";
					when "00111110011100000" => rgb <= "000000";
					when "00111110011100001" => rgb <= "000000";
					when "00111110011100010" => rgb <= "000000";
					when "00111110011100011" => rgb <= "000000";
					when "00111110011100100" => rgb <= "000000";
					when "00111110011100101" => rgb <= "000000";
					when "00111110011100110" => rgb <= "000000";
					when "00111110011100111" => rgb <= "000000";
					when "00111110011101000" => rgb <= "000000";
					when "00111110011101001" => rgb <= "000000";
					when "00111110011101010" => rgb <= "000000";
					when "00111110011101011" => rgb <= "000000";
					when "00111110011101100" => rgb <= "000000";
					when "00111110011101101" => rgb <= "000000";
					when "00111110011101110" => rgb <= "000000";
					when "00111110011101111" => rgb <= "000000";
					when "00111110011110000" => rgb <= "000000";
					when "00111110011110001" => rgb <= "000000";
					when "00111110011110010" => rgb <= "000000";
					when "00111110011110011" => rgb <= "000000";
					when "00111110011110100" => rgb <= "000000";
					when "00111110011110101" => rgb <= "000000";
					when "00111110011110110" => rgb <= "000000";
					when "00111110011110111" => rgb <= "000000";
					when "00111110011111000" => rgb <= "000000";
					when "00111110011111001" => rgb <= "000000";
					when "00111110011111010" => rgb <= "000000";
					when "00111110011111011" => rgb <= "000000";
					when "00111110011111100" => rgb <= "000000";
					when "00111110011111101" => rgb <= "000000";
					when "00111110011111110" => rgb <= "000000";
					when "00111110011111111" => rgb <= "000000";
					when "00111110100000000" => rgb <= "000000";
					when "00111110100000001" => rgb <= "000000";
					when "00111110100000010" => rgb <= "000000";
					when "00111110100000011" => rgb <= "000000";
					when "00111110100000100" => rgb <= "000000";
					when "00111110100000101" => rgb <= "000000";
					when "00111110100000110" => rgb <= "000000";
					when "00111110100000111" => rgb <= "000000";
					when "00111110100001000" => rgb <= "000000";
					when "00111110100001001" => rgb <= "000000";
					when "00111110100001010" => rgb <= "000000";
					when "00111110100001011" => rgb <= "000000";
					when "00111110100001100" => rgb <= "000000";
					when "00111110100001101" => rgb <= "000000";
					when "00111110100001110" => rgb <= "000000";
					when "00111110100001111" => rgb <= "000000";
					when "00111110100010000" => rgb <= "000000";
					when "00111110100010001" => rgb <= "000000";
					when "00111110100010010" => rgb <= "000000";
					when "00111110100010011" => rgb <= "000000";
					when "00111110100010100" => rgb <= "000000";
					when "00111110100010101" => rgb <= "000000";
					when "00111110100010110" => rgb <= "000000";
					when "00111110100010111" => rgb <= "000000";
					when "00111110100011000" => rgb <= "000000";
					when "00111110100011001" => rgb <= "000000";
					when "00111110100011010" => rgb <= "000000";
					when "00111110100011011" => rgb <= "000000";
					when "00111110100011100" => rgb <= "000000";
					when "00111110100011101" => rgb <= "000000";
					when "00111110100011110" => rgb <= "000000";
					when "00111110100011111" => rgb <= "000000";
					when "00111110100100000" => rgb <= "000000";
					when "00111110100100001" => rgb <= "000000";
					when "00111110100100010" => rgb <= "000000";
					when "00111110100100011" => rgb <= "000000";
					when "00111110100100100" => rgb <= "000000";
					when "00111110100100101" => rgb <= "000000";
					when "00111110100100110" => rgb <= "000000";
					when "00111110100100111" => rgb <= "000000";
					when "00111110100101000" => rgb <= "000000";
					when "00111110100101001" => rgb <= "000000";
					when "00111110100101010" => rgb <= "000000";
					when "00111110100101011" => rgb <= "000000";
					when "00111110100101100" => rgb <= "000000";
					when "00111110100101101" => rgb <= "000000";
					when "00111110100101110" => rgb <= "000000";
					when "00111110100101111" => rgb <= "000000";
					when "00111110100110000" => rgb <= "000000";
					when "00111110100110001" => rgb <= "000000";
					when "00111110100110010" => rgb <= "000000";
					when "00111110100110011" => rgb <= "000000";
					when "00111110100110100" => rgb <= "000000";
					when "00111110100110101" => rgb <= "000000";
					when "00111110100110110" => rgb <= "000000";
					when "00111110100110111" => rgb <= "000000";
					when "00111110100111000" => rgb <= "000000";
					when "00111110100111001" => rgb <= "000000";
					when "00111110100111010" => rgb <= "000000";
					when "00111110100111011" => rgb <= "000000";
					when "00111110100111100" => rgb <= "000000";
					when "00111110100111101" => rgb <= "000000";
					when "00111110100111110" => rgb <= "000000";
					when "00111110100111111" => rgb <= "000000";
					when "00111111000000000" => rgb <= "000000";
					when "00111111000000001" => rgb <= "000000";
					when "00111111000000010" => rgb <= "000000";
					when "00111111000000011" => rgb <= "000000";
					when "00111111000000100" => rgb <= "000000";
					when "00111111000000101" => rgb <= "000000";
					when "00111111000000110" => rgb <= "000000";
					when "00111111000000111" => rgb <= "000000";
					when "00111111000001000" => rgb <= "000000";
					when "00111111000001001" => rgb <= "000000";
					when "00111111000001010" => rgb <= "000000";
					when "00111111000001011" => rgb <= "000000";
					when "00111111000001100" => rgb <= "000000";
					when "00111111000001101" => rgb <= "000000";
					when "00111111000001110" => rgb <= "000000";
					when "00111111000001111" => rgb <= "000000";
					when "00111111000010000" => rgb <= "000000";
					when "00111111000010001" => rgb <= "000000";
					when "00111111000010010" => rgb <= "000000";
					when "00111111000010011" => rgb <= "000000";
					when "00111111000010100" => rgb <= "000000";
					when "00111111000010101" => rgb <= "000000";
					when "00111111000010110" => rgb <= "000000";
					when "00111111000010111" => rgb <= "000000";
					when "00111111000011000" => rgb <= "000000";
					when "00111111000011001" => rgb <= "000000";
					when "00111111000011010" => rgb <= "000000";
					when "00111111000011011" => rgb <= "000000";
					when "00111111000011100" => rgb <= "000000";
					when "00111111000011101" => rgb <= "000000";
					when "00111111000011110" => rgb <= "000000";
					when "00111111000011111" => rgb <= "000000";
					when "00111111000100000" => rgb <= "000000";
					when "00111111000100001" => rgb <= "000000";
					when "00111111000100010" => rgb <= "000000";
					when "00111111000100011" => rgb <= "000000";
					when "00111111000100100" => rgb <= "000000";
					when "00111111000100101" => rgb <= "000000";
					when "00111111000100110" => rgb <= "000000";
					when "00111111000100111" => rgb <= "000000";
					when "00111111000101000" => rgb <= "000000";
					when "00111111000101001" => rgb <= "000000";
					when "00111111000101010" => rgb <= "000000";
					when "00111111000101011" => rgb <= "000000";
					when "00111111000101100" => rgb <= "000000";
					when "00111111000101101" => rgb <= "000000";
					when "00111111000101110" => rgb <= "000000";
					when "00111111000101111" => rgb <= "000000";
					when "00111111000110000" => rgb <= "000000";
					when "00111111000110001" => rgb <= "000000";
					when "00111111000110010" => rgb <= "000000";
					when "00111111000110011" => rgb <= "000000";
					when "00111111000110100" => rgb <= "000000";
					when "00111111000110101" => rgb <= "000000";
					when "00111111000110110" => rgb <= "000000";
					when "00111111000110111" => rgb <= "000000";
					when "00111111000111000" => rgb <= "000000";
					when "00111111000111001" => rgb <= "000000";
					when "00111111000111010" => rgb <= "000000";
					when "00111111000111011" => rgb <= "000000";
					when "00111111000111100" => rgb <= "000000";
					when "00111111000111101" => rgb <= "000000";
					when "00111111000111110" => rgb <= "000000";
					when "00111111000111111" => rgb <= "000000";
					when "00111111001000000" => rgb <= "000000";
					when "00111111001000001" => rgb <= "000000";
					when "00111111001000010" => rgb <= "000000";
					when "00111111001000011" => rgb <= "000000";
					when "00111111001000100" => rgb <= "000000";
					when "00111111001000101" => rgb <= "000000";
					when "00111111001000110" => rgb <= "000000";
					when "00111111001000111" => rgb <= "000000";
					when "00111111001001000" => rgb <= "000000";
					when "00111111001001001" => rgb <= "000000";
					when "00111111001001010" => rgb <= "000000";
					when "00111111001001011" => rgb <= "000000";
					when "00111111001001100" => rgb <= "000000";
					when "00111111001001101" => rgb <= "000000";
					when "00111111001001110" => rgb <= "000000";
					when "00111111001001111" => rgb <= "000000";
					when "00111111001010000" => rgb <= "000000";
					when "00111111001010001" => rgb <= "000000";
					when "00111111001010010" => rgb <= "000000";
					when "00111111001010011" => rgb <= "000000";
					when "00111111001010100" => rgb <= "000000";
					when "00111111001010101" => rgb <= "000000";
					when "00111111001010110" => rgb <= "000000";
					when "00111111001010111" => rgb <= "000000";
					when "00111111001011000" => rgb <= "000000";
					when "00111111001011001" => rgb <= "000000";
					when "00111111001011010" => rgb <= "000000";
					when "00111111001011011" => rgb <= "000000";
					when "00111111001011100" => rgb <= "000000";
					when "00111111001011101" => rgb <= "000000";
					when "00111111001011110" => rgb <= "000000";
					when "00111111001011111" => rgb <= "000000";
					when "00111111001100000" => rgb <= "000000";
					when "00111111001100001" => rgb <= "000000";
					when "00111111001100010" => rgb <= "000000";
					when "00111111001100011" => rgb <= "000000";
					when "00111111001100100" => rgb <= "000000";
					when "00111111001100101" => rgb <= "000000";
					when "00111111001100110" => rgb <= "000000";
					when "00111111001100111" => rgb <= "000000";
					when "00111111001101000" => rgb <= "000000";
					when "00111111001101001" => rgb <= "000000";
					when "00111111001101010" => rgb <= "000000";
					when "00111111001101011" => rgb <= "000000";
					when "00111111001101100" => rgb <= "000000";
					when "00111111001101101" => rgb <= "000000";
					when "00111111001101110" => rgb <= "000000";
					when "00111111001101111" => rgb <= "000000";
					when "00111111001110000" => rgb <= "000000";
					when "00111111001110001" => rgb <= "000000";
					when "00111111001110010" => rgb <= "111001";
					when "00111111001110011" => rgb <= "111000";
					when "00111111001110100" => rgb <= "111000";
					when "00111111001110101" => rgb <= "111000";
					when "00111111001110110" => rgb <= "101001";
					when "00111111001110111" => rgb <= "101000";
					when "00111111001111000" => rgb <= "101000";
					when "00111111001111001" => rgb <= "101000";
					when "00111111001111010" => rgb <= "111000";
					when "00111111001111011" => rgb <= "101000";
					when "00111111001111100" => rgb <= "111001";
					when "00111111001111101" => rgb <= "111000";
					when "00111111001111110" => rgb <= "101000";
					when "00111111001111111" => rgb <= "101000";
					when "00111111010000000" => rgb <= "101000";
					when "00111111010000001" => rgb <= "101000";
					when "00111111010000010" => rgb <= "101000";
					when "00111111010000011" => rgb <= "101000";
					when "00111111010000100" => rgb <= "101000";
					when "00111111010000101" => rgb <= "101000";
					when "00111111010000110" => rgb <= "101000";
					when "00111111010000111" => rgb <= "101000";
					when "00111111010001000" => rgb <= "101000";
					when "00111111010001001" => rgb <= "101000";
					when "00111111010001010" => rgb <= "101000";
					when "00111111010001011" => rgb <= "101000";
					when "00111111010001100" => rgb <= "101000";
					when "00111111010001101" => rgb <= "101000";
					when "00111111010001110" => rgb <= "101000";
					when "00111111010001111" => rgb <= "101000";
					when "00111111010010000" => rgb <= "101000";
					when "00111111010010001" => rgb <= "101000";
					when "00111111010010010" => rgb <= "101000";
					when "00111111010010011" => rgb <= "101000";
					when "00111111010010100" => rgb <= "101000";
					when "00111111010010101" => rgb <= "101000";
					when "00111111010010110" => rgb <= "101000";
					when "00111111010010111" => rgb <= "101000";
					when "00111111010011000" => rgb <= "101000";
					when "00111111010011001" => rgb <= "101000";
					when "00111111010011010" => rgb <= "101000";
					when "00111111010011011" => rgb <= "101000";
					when "00111111010011100" => rgb <= "101000";
					when "00111111010011101" => rgb <= "101000";
					when "00111111010011110" => rgb <= "101000";
					when "00111111010011111" => rgb <= "101000";
					when "00111111010100000" => rgb <= "101000";
					when "00111111010100001" => rgb <= "101000";
					when "00111111010100010" => rgb <= "101000";
					when "00111111010100011" => rgb <= "101000";
					when "00111111010100100" => rgb <= "101000";
					when "00111111010100101" => rgb <= "101000";
					when "00111111010100110" => rgb <= "101000";
					when "00111111010100111" => rgb <= "101000";
					when "00111111010101000" => rgb <= "101000";
					when "00111111010101001" => rgb <= "101000";
					when "00111111010101010" => rgb <= "101000";
					when "00111111010101011" => rgb <= "101000";
					when "00111111010101100" => rgb <= "101000";
					when "00111111010101101" => rgb <= "101000";
					when "00111111010101110" => rgb <= "101000";
					when "00111111010101111" => rgb <= "101000";
					when "00111111010110000" => rgb <= "101000";
					when "00111111010110001" => rgb <= "101000";
					when "00111111010110010" => rgb <= "101000";
					when "00111111010110011" => rgb <= "101000";
					when "00111111010110100" => rgb <= "101000";
					when "00111111010110101" => rgb <= "101000";
					when "00111111010110110" => rgb <= "101000";
					when "00111111010110111" => rgb <= "101000";
					when "00111111010111000" => rgb <= "101000";
					when "00111111010111001" => rgb <= "101000";
					when "00111111010111010" => rgb <= "101000";
					when "00111111010111011" => rgb <= "101000";
					when "00111111010111100" => rgb <= "101000";
					when "00111111010111101" => rgb <= "101000";
					when "00111111010111110" => rgb <= "101000";
					when "00111111010111111" => rgb <= "101000";
					when "00111111011000000" => rgb <= "101000";
					when "00111111011000001" => rgb <= "101000";
					when "00111111011000010" => rgb <= "101000";
					when "00111111011000011" => rgb <= "101000";
					when "00111111011000100" => rgb <= "101000";
					when "00111111011000101" => rgb <= "101000";
					when "00111111011000110" => rgb <= "101000";
					when "00111111011000111" => rgb <= "101000";
					when "00111111011001000" => rgb <= "101000";
					when "00111111011001001" => rgb <= "101000";
					when "00111111011001010" => rgb <= "101000";
					when "00111111011001011" => rgb <= "101000";
					when "00111111011001100" => rgb <= "000000";
					when "00111111011001101" => rgb <= "000000";
					when "00111111011001110" => rgb <= "000000";
					when "00111111011001111" => rgb <= "000000";
					when "00111111011010000" => rgb <= "000000";
					when "00111111011010001" => rgb <= "000000";
					when "00111111011010010" => rgb <= "000000";
					when "00111111011010011" => rgb <= "000000";
					when "00111111011010100" => rgb <= "000000";
					when "00111111011010101" => rgb <= "000000";
					when "00111111011010110" => rgb <= "000000";
					when "00111111011010111" => rgb <= "000000";
					when "00111111011011000" => rgb <= "000000";
					when "00111111011011001" => rgb <= "000000";
					when "00111111011011010" => rgb <= "000000";
					when "00111111011011011" => rgb <= "000000";
					when "00111111011011100" => rgb <= "000000";
					when "00111111011011101" => rgb <= "000000";
					when "00111111011011110" => rgb <= "000000";
					when "00111111011011111" => rgb <= "000000";
					when "00111111011100000" => rgb <= "000000";
					when "00111111011100001" => rgb <= "000000";
					when "00111111011100010" => rgb <= "000000";
					when "00111111011100011" => rgb <= "000000";
					when "00111111011100100" => rgb <= "000000";
					when "00111111011100101" => rgb <= "000000";
					when "00111111011100110" => rgb <= "000000";
					when "00111111011100111" => rgb <= "000000";
					when "00111111011101000" => rgb <= "000000";
					when "00111111011101001" => rgb <= "000000";
					when "00111111011101010" => rgb <= "000000";
					when "00111111011101011" => rgb <= "000000";
					when "00111111011101100" => rgb <= "000000";
					when "00111111011101101" => rgb <= "000000";
					when "00111111011101110" => rgb <= "000000";
					when "00111111011101111" => rgb <= "000000";
					when "00111111011110000" => rgb <= "000000";
					when "00111111011110001" => rgb <= "000000";
					when "00111111011110010" => rgb <= "000000";
					when "00111111011110011" => rgb <= "000000";
					when "00111111011110100" => rgb <= "000000";
					when "00111111011110101" => rgb <= "000000";
					when "00111111011110110" => rgb <= "000000";
					when "00111111011110111" => rgb <= "000000";
					when "00111111011111000" => rgb <= "000000";
					when "00111111011111001" => rgb <= "000000";
					when "00111111011111010" => rgb <= "000000";
					when "00111111011111011" => rgb <= "000000";
					when "00111111011111100" => rgb <= "000000";
					when "00111111011111101" => rgb <= "000000";
					when "00111111011111110" => rgb <= "000000";
					when "00111111011111111" => rgb <= "000000";
					when "00111111100000000" => rgb <= "000000";
					when "00111111100000001" => rgb <= "000000";
					when "00111111100000010" => rgb <= "000000";
					when "00111111100000011" => rgb <= "000000";
					when "00111111100000100" => rgb <= "000000";
					when "00111111100000101" => rgb <= "000000";
					when "00111111100000110" => rgb <= "000000";
					when "00111111100000111" => rgb <= "000000";
					when "00111111100001000" => rgb <= "000000";
					when "00111111100001001" => rgb <= "000000";
					when "00111111100001010" => rgb <= "000000";
					when "00111111100001011" => rgb <= "000000";
					when "00111111100001100" => rgb <= "000000";
					when "00111111100001101" => rgb <= "000000";
					when "00111111100001110" => rgb <= "000000";
					when "00111111100001111" => rgb <= "000000";
					when "00111111100010000" => rgb <= "000000";
					when "00111111100010001" => rgb <= "000000";
					when "00111111100010010" => rgb <= "000000";
					when "00111111100010011" => rgb <= "000000";
					when "00111111100010100" => rgb <= "000000";
					when "00111111100010101" => rgb <= "000000";
					when "00111111100010110" => rgb <= "000000";
					when "00111111100010111" => rgb <= "000000";
					when "00111111100011000" => rgb <= "000000";
					when "00111111100011001" => rgb <= "000000";
					when "00111111100011010" => rgb <= "000000";
					when "00111111100011011" => rgb <= "000000";
					when "00111111100011100" => rgb <= "000000";
					when "00111111100011101" => rgb <= "000000";
					when "00111111100011110" => rgb <= "000000";
					when "00111111100011111" => rgb <= "000000";
					when "00111111100100000" => rgb <= "000000";
					when "00111111100100001" => rgb <= "000000";
					when "00111111100100010" => rgb <= "000000";
					when "00111111100100011" => rgb <= "000000";
					when "00111111100100100" => rgb <= "000000";
					when "00111111100100101" => rgb <= "000000";
					when "00111111100100110" => rgb <= "000000";
					when "00111111100100111" => rgb <= "000000";
					when "00111111100101000" => rgb <= "000000";
					when "00111111100101001" => rgb <= "000000";
					when "00111111100101010" => rgb <= "000000";
					when "00111111100101011" => rgb <= "000000";
					when "00111111100101100" => rgb <= "000000";
					when "00111111100101101" => rgb <= "000000";
					when "00111111100101110" => rgb <= "000000";
					when "00111111100101111" => rgb <= "000000";
					when "00111111100110000" => rgb <= "000000";
					when "00111111100110001" => rgb <= "000000";
					when "00111111100110010" => rgb <= "000000";
					when "00111111100110011" => rgb <= "000000";
					when "00111111100110100" => rgb <= "000000";
					when "00111111100110101" => rgb <= "000000";
					when "00111111100110110" => rgb <= "000000";
					when "00111111100110111" => rgb <= "000000";
					when "00111111100111000" => rgb <= "000000";
					when "00111111100111001" => rgb <= "000000";
					when "00111111100111010" => rgb <= "000000";
					when "00111111100111011" => rgb <= "000000";
					when "00111111100111100" => rgb <= "000000";
					when "00111111100111101" => rgb <= "000000";
					when "00111111100111110" => rgb <= "000000";
					when "00111111100111111" => rgb <= "000000";
					when "01000000000000000" => rgb <= "000000";
					when "01000000000000001" => rgb <= "000000";
					when "01000000000000010" => rgb <= "000000";
					when "01000000000000011" => rgb <= "000000";
					when "01000000000000100" => rgb <= "000000";
					when "01000000000000101" => rgb <= "000000";
					when "01000000000000110" => rgb <= "000000";
					when "01000000000000111" => rgb <= "000000";
					when "01000000000001000" => rgb <= "000000";
					when "01000000000001001" => rgb <= "000000";
					when "01000000000001010" => rgb <= "000000";
					when "01000000000001011" => rgb <= "000000";
					when "01000000000001100" => rgb <= "000000";
					when "01000000000001101" => rgb <= "000000";
					when "01000000000001110" => rgb <= "000000";
					when "01000000000001111" => rgb <= "000000";
					when "01000000000010000" => rgb <= "000000";
					when "01000000000010001" => rgb <= "000000";
					when "01000000000010010" => rgb <= "000000";
					when "01000000000010011" => rgb <= "000000";
					when "01000000000010100" => rgb <= "000000";
					when "01000000000010101" => rgb <= "000000";
					when "01000000000010110" => rgb <= "000000";
					when "01000000000010111" => rgb <= "000000";
					when "01000000000011000" => rgb <= "000000";
					when "01000000000011001" => rgb <= "000000";
					when "01000000000011010" => rgb <= "000000";
					when "01000000000011011" => rgb <= "000000";
					when "01000000000011100" => rgb <= "000000";
					when "01000000000011101" => rgb <= "000000";
					when "01000000000011110" => rgb <= "000000";
					when "01000000000011111" => rgb <= "000000";
					when "01000000000100000" => rgb <= "000000";
					when "01000000000100001" => rgb <= "000000";
					when "01000000000100010" => rgb <= "000000";
					when "01000000000100011" => rgb <= "000000";
					when "01000000000100100" => rgb <= "000000";
					when "01000000000100101" => rgb <= "000000";
					when "01000000000100110" => rgb <= "000000";
					when "01000000000100111" => rgb <= "000000";
					when "01000000000101000" => rgb <= "000000";
					when "01000000000101001" => rgb <= "000000";
					when "01000000000101010" => rgb <= "000000";
					when "01000000000101011" => rgb <= "000000";
					when "01000000000101100" => rgb <= "000000";
					when "01000000000101101" => rgb <= "000000";
					when "01000000000101110" => rgb <= "000000";
					when "01000000000101111" => rgb <= "000000";
					when "01000000000110000" => rgb <= "000000";
					when "01000000000110001" => rgb <= "000000";
					when "01000000000110010" => rgb <= "000000";
					when "01000000000110011" => rgb <= "000000";
					when "01000000000110100" => rgb <= "000000";
					when "01000000000110101" => rgb <= "000000";
					when "01000000000110110" => rgb <= "000000";
					when "01000000000110111" => rgb <= "000000";
					when "01000000000111000" => rgb <= "000000";
					when "01000000000111001" => rgb <= "000000";
					when "01000000000111010" => rgb <= "000000";
					when "01000000000111011" => rgb <= "000000";
					when "01000000000111100" => rgb <= "000000";
					when "01000000000111101" => rgb <= "000000";
					when "01000000000111110" => rgb <= "000000";
					when "01000000000111111" => rgb <= "000000";
					when "01000000001000000" => rgb <= "000000";
					when "01000000001000001" => rgb <= "000000";
					when "01000000001000010" => rgb <= "000000";
					when "01000000001000011" => rgb <= "000000";
					when "01000000001000100" => rgb <= "000000";
					when "01000000001000101" => rgb <= "000000";
					when "01000000001000110" => rgb <= "000000";
					when "01000000001000111" => rgb <= "000000";
					when "01000000001001000" => rgb <= "000000";
					when "01000000001001001" => rgb <= "000000";
					when "01000000001001010" => rgb <= "000000";
					when "01000000001001011" => rgb <= "000000";
					when "01000000001001100" => rgb <= "000000";
					when "01000000001001101" => rgb <= "000000";
					when "01000000001001110" => rgb <= "000000";
					when "01000000001001111" => rgb <= "000000";
					when "01000000001010000" => rgb <= "000000";
					when "01000000001010001" => rgb <= "000000";
					when "01000000001010010" => rgb <= "000000";
					when "01000000001010011" => rgb <= "000000";
					when "01000000001010100" => rgb <= "000000";
					when "01000000001010101" => rgb <= "000000";
					when "01000000001010110" => rgb <= "000000";
					when "01000000001010111" => rgb <= "000000";
					when "01000000001011000" => rgb <= "000000";
					when "01000000001011001" => rgb <= "000000";
					when "01000000001011010" => rgb <= "000000";
					when "01000000001011011" => rgb <= "000000";
					when "01000000001011100" => rgb <= "000000";
					when "01000000001011101" => rgb <= "000000";
					when "01000000001011110" => rgb <= "000000";
					when "01000000001011111" => rgb <= "000000";
					when "01000000001100000" => rgb <= "000000";
					when "01000000001100001" => rgb <= "000000";
					when "01000000001100010" => rgb <= "000000";
					when "01000000001100011" => rgb <= "000000";
					when "01000000001100100" => rgb <= "000000";
					when "01000000001100101" => rgb <= "000000";
					when "01000000001100110" => rgb <= "000000";
					when "01000000001100111" => rgb <= "000000";
					when "01000000001101000" => rgb <= "000000";
					when "01000000001101001" => rgb <= "000000";
					when "01000000001101010" => rgb <= "000000";
					when "01000000001101011" => rgb <= "000000";
					when "01000000001101100" => rgb <= "000000";
					when "01000000001101101" => rgb <= "000000";
					when "01000000001101110" => rgb <= "000000";
					when "01000000001101111" => rgb <= "000000";
					when "01000000001110000" => rgb <= "000000";
					when "01000000001110001" => rgb <= "010000";
					when "01000000001110010" => rgb <= "101000";
					when "01000000001110011" => rgb <= "101000";
					when "01000000001110100" => rgb <= "101000";
					when "01000000001110101" => rgb <= "101000";
					when "01000000001110110" => rgb <= "101000";
					when "01000000001110111" => rgb <= "101000";
					when "01000000001111000" => rgb <= "101000";
					when "01000000001111001" => rgb <= "101000";
					when "01000000001111010" => rgb <= "101000";
					when "01000000001111011" => rgb <= "101000";
					when "01000000001111100" => rgb <= "101000";
					when "01000000001111101" => rgb <= "101000";
					when "01000000001111110" => rgb <= "101000";
					when "01000000001111111" => rgb <= "101000";
					when "01000000010000000" => rgb <= "101000";
					when "01000000010000001" => rgb <= "101000";
					when "01000000010000010" => rgb <= "101000";
					when "01000000010000011" => rgb <= "101000";
					when "01000000010000100" => rgb <= "101000";
					when "01000000010000101" => rgb <= "101000";
					when "01000000010000110" => rgb <= "101000";
					when "01000000010000111" => rgb <= "101000";
					when "01000000010001000" => rgb <= "101000";
					when "01000000010001001" => rgb <= "101000";
					when "01000000010001010" => rgb <= "101000";
					when "01000000010001011" => rgb <= "101000";
					when "01000000010001100" => rgb <= "101000";
					when "01000000010001101" => rgb <= "101000";
					when "01000000010001110" => rgb <= "101000";
					when "01000000010001111" => rgb <= "101000";
					when "01000000010010000" => rgb <= "101000";
					when "01000000010010001" => rgb <= "101000";
					when "01000000010010010" => rgb <= "101000";
					when "01000000010010011" => rgb <= "101000";
					when "01000000010010100" => rgb <= "101000";
					when "01000000010010101" => rgb <= "101000";
					when "01000000010010110" => rgb <= "101000";
					when "01000000010010111" => rgb <= "101000";
					when "01000000010011000" => rgb <= "101000";
					when "01000000010011001" => rgb <= "101000";
					when "01000000010011010" => rgb <= "101000";
					when "01000000010011011" => rgb <= "101000";
					when "01000000010011100" => rgb <= "101000";
					when "01000000010011101" => rgb <= "101000";
					when "01000000010011110" => rgb <= "101000";
					when "01000000010011111" => rgb <= "101000";
					when "01000000010100000" => rgb <= "101000";
					when "01000000010100001" => rgb <= "101000";
					when "01000000010100010" => rgb <= "101000";
					when "01000000010100011" => rgb <= "101000";
					when "01000000010100100" => rgb <= "101000";
					when "01000000010100101" => rgb <= "101000";
					when "01000000010100110" => rgb <= "101000";
					when "01000000010100111" => rgb <= "101000";
					when "01000000010101000" => rgb <= "101000";
					when "01000000010101001" => rgb <= "101000";
					when "01000000010101010" => rgb <= "101000";
					when "01000000010101011" => rgb <= "101000";
					when "01000000010101100" => rgb <= "101000";
					when "01000000010101101" => rgb <= "101000";
					when "01000000010101110" => rgb <= "101000";
					when "01000000010101111" => rgb <= "101000";
					when "01000000010110000" => rgb <= "101000";
					when "01000000010110001" => rgb <= "101000";
					when "01000000010110010" => rgb <= "101000";
					when "01000000010110011" => rgb <= "101000";
					when "01000000010110100" => rgb <= "101000";
					when "01000000010110101" => rgb <= "101000";
					when "01000000010110110" => rgb <= "101000";
					when "01000000010110111" => rgb <= "101000";
					when "01000000010111000" => rgb <= "101000";
					when "01000000010111001" => rgb <= "101000";
					when "01000000010111010" => rgb <= "101000";
					when "01000000010111011" => rgb <= "101000";
					when "01000000010111100" => rgb <= "101000";
					when "01000000010111101" => rgb <= "101000";
					when "01000000010111110" => rgb <= "101000";
					when "01000000010111111" => rgb <= "101000";
					when "01000000011000000" => rgb <= "101000";
					when "01000000011000001" => rgb <= "101000";
					when "01000000011000010" => rgb <= "101000";
					when "01000000011000011" => rgb <= "101000";
					when "01000000011000100" => rgb <= "101000";
					when "01000000011000101" => rgb <= "101000";
					when "01000000011000110" => rgb <= "101000";
					when "01000000011000111" => rgb <= "101000";
					when "01000000011001000" => rgb <= "101000";
					when "01000000011001001" => rgb <= "101000";
					when "01000000011001010" => rgb <= "101000";
					when "01000000011001011" => rgb <= "101000";
					when "01000000011001100" => rgb <= "000000";
					when "01000000011001101" => rgb <= "000000";
					when "01000000011001110" => rgb <= "000000";
					when "01000000011001111" => rgb <= "000000";
					when "01000000011010000" => rgb <= "000000";
					when "01000000011010001" => rgb <= "000000";
					when "01000000011010010" => rgb <= "000000";
					when "01000000011010011" => rgb <= "000000";
					when "01000000011010100" => rgb <= "000000";
					when "01000000011010101" => rgb <= "000000";
					when "01000000011010110" => rgb <= "000000";
					when "01000000011010111" => rgb <= "000000";
					when "01000000011011000" => rgb <= "000000";
					when "01000000011011001" => rgb <= "000000";
					when "01000000011011010" => rgb <= "000000";
					when "01000000011011011" => rgb <= "000000";
					when "01000000011011100" => rgb <= "000000";
					when "01000000011011101" => rgb <= "000000";
					when "01000000011011110" => rgb <= "000000";
					when "01000000011011111" => rgb <= "000000";
					when "01000000011100000" => rgb <= "000000";
					when "01000000011100001" => rgb <= "000000";
					when "01000000011100010" => rgb <= "000000";
					when "01000000011100011" => rgb <= "000000";
					when "01000000011100100" => rgb <= "000000";
					when "01000000011100101" => rgb <= "000000";
					when "01000000011100110" => rgb <= "000000";
					when "01000000011100111" => rgb <= "000000";
					when "01000000011101000" => rgb <= "000000";
					when "01000000011101001" => rgb <= "000000";
					when "01000000011101010" => rgb <= "000000";
					when "01000000011101011" => rgb <= "000000";
					when "01000000011101100" => rgb <= "000000";
					when "01000000011101101" => rgb <= "000000";
					when "01000000011101110" => rgb <= "000000";
					when "01000000011101111" => rgb <= "000000";
					when "01000000011110000" => rgb <= "000000";
					when "01000000011110001" => rgb <= "000000";
					when "01000000011110010" => rgb <= "000000";
					when "01000000011110011" => rgb <= "000000";
					when "01000000011110100" => rgb <= "000000";
					when "01000000011110101" => rgb <= "000000";
					when "01000000011110110" => rgb <= "000000";
					when "01000000011110111" => rgb <= "000000";
					when "01000000011111000" => rgb <= "000000";
					when "01000000011111001" => rgb <= "000000";
					when "01000000011111010" => rgb <= "000000";
					when "01000000011111011" => rgb <= "000000";
					when "01000000011111100" => rgb <= "000000";
					when "01000000011111101" => rgb <= "000000";
					when "01000000011111110" => rgb <= "000000";
					when "01000000011111111" => rgb <= "000000";
					when "01000000100000000" => rgb <= "000000";
					when "01000000100000001" => rgb <= "000000";
					when "01000000100000010" => rgb <= "000000";
					when "01000000100000011" => rgb <= "000000";
					when "01000000100000100" => rgb <= "000000";
					when "01000000100000101" => rgb <= "000000";
					when "01000000100000110" => rgb <= "000000";
					when "01000000100000111" => rgb <= "000000";
					when "01000000100001000" => rgb <= "000000";
					when "01000000100001001" => rgb <= "000000";
					when "01000000100001010" => rgb <= "000000";
					when "01000000100001011" => rgb <= "000000";
					when "01000000100001100" => rgb <= "000000";
					when "01000000100001101" => rgb <= "000000";
					when "01000000100001110" => rgb <= "000000";
					when "01000000100001111" => rgb <= "000000";
					when "01000000100010000" => rgb <= "000000";
					when "01000000100010001" => rgb <= "000000";
					when "01000000100010010" => rgb <= "000000";
					when "01000000100010011" => rgb <= "000000";
					when "01000000100010100" => rgb <= "000000";
					when "01000000100010101" => rgb <= "000000";
					when "01000000100010110" => rgb <= "000000";
					when "01000000100010111" => rgb <= "000000";
					when "01000000100011000" => rgb <= "000000";
					when "01000000100011001" => rgb <= "000000";
					when "01000000100011010" => rgb <= "000000";
					when "01000000100011011" => rgb <= "000000";
					when "01000000100011100" => rgb <= "000000";
					when "01000000100011101" => rgb <= "000000";
					when "01000000100011110" => rgb <= "000000";
					when "01000000100011111" => rgb <= "000000";
					when "01000000100100000" => rgb <= "000000";
					when "01000000100100001" => rgb <= "000000";
					when "01000000100100010" => rgb <= "000000";
					when "01000000100100011" => rgb <= "000000";
					when "01000000100100100" => rgb <= "000000";
					when "01000000100100101" => rgb <= "000000";
					when "01000000100100110" => rgb <= "000000";
					when "01000000100100111" => rgb <= "000000";
					when "01000000100101000" => rgb <= "000000";
					when "01000000100101001" => rgb <= "000000";
					when "01000000100101010" => rgb <= "000000";
					when "01000000100101011" => rgb <= "000000";
					when "01000000100101100" => rgb <= "000000";
					when "01000000100101101" => rgb <= "000000";
					when "01000000100101110" => rgb <= "000000";
					when "01000000100101111" => rgb <= "000000";
					when "01000000100110000" => rgb <= "000000";
					when "01000000100110001" => rgb <= "000000";
					when "01000000100110010" => rgb <= "000000";
					when "01000000100110011" => rgb <= "000000";
					when "01000000100110100" => rgb <= "000000";
					when "01000000100110101" => rgb <= "000000";
					when "01000000100110110" => rgb <= "000000";
					when "01000000100110111" => rgb <= "000000";
					when "01000000100111000" => rgb <= "000000";
					when "01000000100111001" => rgb <= "000000";
					when "01000000100111010" => rgb <= "000000";
					when "01000000100111011" => rgb <= "000000";
					when "01000000100111100" => rgb <= "000000";
					when "01000000100111101" => rgb <= "000000";
					when "01000000100111110" => rgb <= "000000";
					when "01000000100111111" => rgb <= "000000";
					when "01000001000000000" => rgb <= "000000";
					when "01000001000000001" => rgb <= "000000";
					when "01000001000000010" => rgb <= "000000";
					when "01000001000000011" => rgb <= "000000";
					when "01000001000000100" => rgb <= "000000";
					when "01000001000000101" => rgb <= "000000";
					when "01000001000000110" => rgb <= "000000";
					when "01000001000000111" => rgb <= "000000";
					when "01000001000001000" => rgb <= "000000";
					when "01000001000001001" => rgb <= "000000";
					when "01000001000001010" => rgb <= "000000";
					when "01000001000001011" => rgb <= "000000";
					when "01000001000001100" => rgb <= "000000";
					when "01000001000001101" => rgb <= "000000";
					when "01000001000001110" => rgb <= "000000";
					when "01000001000001111" => rgb <= "000000";
					when "01000001000010000" => rgb <= "000000";
					when "01000001000010001" => rgb <= "000000";
					when "01000001000010010" => rgb <= "000000";
					when "01000001000010011" => rgb <= "000000";
					when "01000001000010100" => rgb <= "000000";
					when "01000001000010101" => rgb <= "000000";
					when "01000001000010110" => rgb <= "000000";
					when "01000001000010111" => rgb <= "000000";
					when "01000001000011000" => rgb <= "000000";
					when "01000001000011001" => rgb <= "000000";
					when "01000001000011010" => rgb <= "000000";
					when "01000001000011011" => rgb <= "000000";
					when "01000001000011100" => rgb <= "000000";
					when "01000001000011101" => rgb <= "000000";
					when "01000001000011110" => rgb <= "000000";
					when "01000001000011111" => rgb <= "000000";
					when "01000001000100000" => rgb <= "000000";
					when "01000001000100001" => rgb <= "000000";
					when "01000001000100010" => rgb <= "000000";
					when "01000001000100011" => rgb <= "000000";
					when "01000001000100100" => rgb <= "000000";
					when "01000001000100101" => rgb <= "000000";
					when "01000001000100110" => rgb <= "000000";
					when "01000001000100111" => rgb <= "000000";
					when "01000001000101000" => rgb <= "000000";
					when "01000001000101001" => rgb <= "000000";
					when "01000001000101010" => rgb <= "000000";
					when "01000001000101011" => rgb <= "000000";
					when "01000001000101100" => rgb <= "000000";
					when "01000001000101101" => rgb <= "000000";
					when "01000001000101110" => rgb <= "000000";
					when "01000001000101111" => rgb <= "000000";
					when "01000001000110000" => rgb <= "000000";
					when "01000001000110001" => rgb <= "000000";
					when "01000001000110010" => rgb <= "000000";
					when "01000001000110011" => rgb <= "000000";
					when "01000001000110100" => rgb <= "000000";
					when "01000001000110101" => rgb <= "000000";
					when "01000001000110110" => rgb <= "000000";
					when "01000001000110111" => rgb <= "000000";
					when "01000001000111000" => rgb <= "000000";
					when "01000001000111001" => rgb <= "000000";
					when "01000001000111010" => rgb <= "000000";
					when "01000001000111011" => rgb <= "000000";
					when "01000001000111100" => rgb <= "000000";
					when "01000001000111101" => rgb <= "000000";
					when "01000001000111110" => rgb <= "000000";
					when "01000001000111111" => rgb <= "000000";
					when "01000001001000000" => rgb <= "000000";
					when "01000001001000001" => rgb <= "000000";
					when "01000001001000010" => rgb <= "000000";
					when "01000001001000011" => rgb <= "000000";
					when "01000001001000100" => rgb <= "000000";
					when "01000001001000101" => rgb <= "000000";
					when "01000001001000110" => rgb <= "000000";
					when "01000001001000111" => rgb <= "000000";
					when "01000001001001000" => rgb <= "000000";
					when "01000001001001001" => rgb <= "000000";
					when "01000001001001010" => rgb <= "000000";
					when "01000001001001011" => rgb <= "000000";
					when "01000001001001100" => rgb <= "000000";
					when "01000001001001101" => rgb <= "000000";
					when "01000001001001110" => rgb <= "000000";
					when "01000001001001111" => rgb <= "000000";
					when "01000001001010000" => rgb <= "000000";
					when "01000001001010001" => rgb <= "000000";
					when "01000001001010010" => rgb <= "000000";
					when "01000001001010011" => rgb <= "000000";
					when "01000001001010100" => rgb <= "000000";
					when "01000001001010101" => rgb <= "000000";
					when "01000001001010110" => rgb <= "000000";
					when "01000001001010111" => rgb <= "000000";
					when "01000001001011000" => rgb <= "000000";
					when "01000001001011001" => rgb <= "000000";
					when "01000001001011010" => rgb <= "000000";
					when "01000001001011011" => rgb <= "000000";
					when "01000001001011100" => rgb <= "000000";
					when "01000001001011101" => rgb <= "000000";
					when "01000001001011110" => rgb <= "000000";
					when "01000001001011111" => rgb <= "000000";
					when "01000001001100000" => rgb <= "000000";
					when "01000001001100001" => rgb <= "000000";
					when "01000001001100010" => rgb <= "000000";
					when "01000001001100011" => rgb <= "000000";
					when "01000001001100100" => rgb <= "000000";
					when "01000001001100101" => rgb <= "000000";
					when "01000001001100110" => rgb <= "000000";
					when "01000001001100111" => rgb <= "000000";
					when "01000001001101000" => rgb <= "000000";
					when "01000001001101001" => rgb <= "000000";
					when "01000001001101010" => rgb <= "000000";
					when "01000001001101011" => rgb <= "000000";
					when "01000001001101100" => rgb <= "000000";
					when "01000001001101101" => rgb <= "000000";
					when "01000001001101110" => rgb <= "000000";
					when "01000001001101111" => rgb <= "000000";
					when "01000001001110000" => rgb <= "000000";
					when "01000001001110001" => rgb <= "010000";
					when "01000001001110010" => rgb <= "101000";
					when "01000001001110011" => rgb <= "101000";
					when "01000001001110100" => rgb <= "101000";
					when "01000001001110101" => rgb <= "101000";
					when "01000001001110110" => rgb <= "101000";
					when "01000001001110111" => rgb <= "101000";
					when "01000001001111000" => rgb <= "101000";
					when "01000001001111001" => rgb <= "101000";
					when "01000001001111010" => rgb <= "101000";
					when "01000001001111011" => rgb <= "101000";
					when "01000001001111100" => rgb <= "101000";
					when "01000001001111101" => rgb <= "101000";
					when "01000001001111110" => rgb <= "101000";
					when "01000001001111111" => rgb <= "101000";
					when "01000001010000000" => rgb <= "101000";
					when "01000001010000001" => rgb <= "101000";
					when "01000001010000010" => rgb <= "101000";
					when "01000001010000011" => rgb <= "101000";
					when "01000001010000100" => rgb <= "101000";
					when "01000001010000101" => rgb <= "101000";
					when "01000001010000110" => rgb <= "101000";
					when "01000001010000111" => rgb <= "101000";
					when "01000001010001000" => rgb <= "101000";
					when "01000001010001001" => rgb <= "101000";
					when "01000001010001010" => rgb <= "101000";
					when "01000001010001011" => rgb <= "101000";
					when "01000001010001100" => rgb <= "101000";
					when "01000001010001101" => rgb <= "101000";
					when "01000001010001110" => rgb <= "101000";
					when "01000001010001111" => rgb <= "101000";
					when "01000001010010000" => rgb <= "101000";
					when "01000001010010001" => rgb <= "101000";
					when "01000001010010010" => rgb <= "101000";
					when "01000001010010011" => rgb <= "101000";
					when "01000001010010100" => rgb <= "101000";
					when "01000001010010101" => rgb <= "101000";
					when "01000001010010110" => rgb <= "101000";
					when "01000001010010111" => rgb <= "101000";
					when "01000001010011000" => rgb <= "101000";
					when "01000001010011001" => rgb <= "101000";
					when "01000001010011010" => rgb <= "101000";
					when "01000001010011011" => rgb <= "101000";
					when "01000001010011100" => rgb <= "101000";
					when "01000001010011101" => rgb <= "101000";
					when "01000001010011110" => rgb <= "101000";
					when "01000001010011111" => rgb <= "101000";
					when "01000001010100000" => rgb <= "101000";
					when "01000001010100001" => rgb <= "101000";
					when "01000001010100010" => rgb <= "101000";
					when "01000001010100011" => rgb <= "101000";
					when "01000001010100100" => rgb <= "101000";
					when "01000001010100101" => rgb <= "101000";
					when "01000001010100110" => rgb <= "101000";
					when "01000001010100111" => rgb <= "101000";
					when "01000001010101000" => rgb <= "101000";
					when "01000001010101001" => rgb <= "101000";
					when "01000001010101010" => rgb <= "101000";
					when "01000001010101011" => rgb <= "101000";
					when "01000001010101100" => rgb <= "101000";
					when "01000001010101101" => rgb <= "101000";
					when "01000001010101110" => rgb <= "101000";
					when "01000001010101111" => rgb <= "101000";
					when "01000001010110000" => rgb <= "101000";
					when "01000001010110001" => rgb <= "101000";
					when "01000001010110010" => rgb <= "101000";
					when "01000001010110011" => rgb <= "101000";
					when "01000001010110100" => rgb <= "101000";
					when "01000001010110101" => rgb <= "101000";
					when "01000001010110110" => rgb <= "101000";
					when "01000001010110111" => rgb <= "101000";
					when "01000001010111000" => rgb <= "101000";
					when "01000001010111001" => rgb <= "101000";
					when "01000001010111010" => rgb <= "101000";
					when "01000001010111011" => rgb <= "101000";
					when "01000001010111100" => rgb <= "101000";
					when "01000001010111101" => rgb <= "101000";
					when "01000001010111110" => rgb <= "101000";
					when "01000001010111111" => rgb <= "101000";
					when "01000001011000000" => rgb <= "101000";
					when "01000001011000001" => rgb <= "101000";
					when "01000001011000010" => rgb <= "101000";
					when "01000001011000011" => rgb <= "101000";
					when "01000001011000100" => rgb <= "101000";
					when "01000001011000101" => rgb <= "101000";
					when "01000001011000110" => rgb <= "101000";
					when "01000001011000111" => rgb <= "101000";
					when "01000001011001000" => rgb <= "101000";
					when "01000001011001001" => rgb <= "101000";
					when "01000001011001010" => rgb <= "101000";
					when "01000001011001011" => rgb <= "101000";
					when "01000001011001100" => rgb <= "000000";
					when "01000001011001101" => rgb <= "000000";
					when "01000001011001110" => rgb <= "000000";
					when "01000001011001111" => rgb <= "000000";
					when "01000001011010000" => rgb <= "000000";
					when "01000001011010001" => rgb <= "000000";
					when "01000001011010010" => rgb <= "000000";
					when "01000001011010011" => rgb <= "000000";
					when "01000001011010100" => rgb <= "000000";
					when "01000001011010101" => rgb <= "000000";
					when "01000001011010110" => rgb <= "000000";
					when "01000001011010111" => rgb <= "000000";
					when "01000001011011000" => rgb <= "000000";
					when "01000001011011001" => rgb <= "000000";
					when "01000001011011010" => rgb <= "000000";
					when "01000001011011011" => rgb <= "000000";
					when "01000001011011100" => rgb <= "000000";
					when "01000001011011101" => rgb <= "000000";
					when "01000001011011110" => rgb <= "000000";
					when "01000001011011111" => rgb <= "000000";
					when "01000001011100000" => rgb <= "000000";
					when "01000001011100001" => rgb <= "000000";
					when "01000001011100010" => rgb <= "000000";
					when "01000001011100011" => rgb <= "000000";
					when "01000001011100100" => rgb <= "000000";
					when "01000001011100101" => rgb <= "000000";
					when "01000001011100110" => rgb <= "000000";
					when "01000001011100111" => rgb <= "000000";
					when "01000001011101000" => rgb <= "000000";
					when "01000001011101001" => rgb <= "000000";
					when "01000001011101010" => rgb <= "000000";
					when "01000001011101011" => rgb <= "000000";
					when "01000001011101100" => rgb <= "000000";
					when "01000001011101101" => rgb <= "000000";
					when "01000001011101110" => rgb <= "000000";
					when "01000001011101111" => rgb <= "000000";
					when "01000001011110000" => rgb <= "000000";
					when "01000001011110001" => rgb <= "000000";
					when "01000001011110010" => rgb <= "000000";
					when "01000001011110011" => rgb <= "000000";
					when "01000001011110100" => rgb <= "000000";
					when "01000001011110101" => rgb <= "000000";
					when "01000001011110110" => rgb <= "000000";
					when "01000001011110111" => rgb <= "000000";
					when "01000001011111000" => rgb <= "000000";
					when "01000001011111001" => rgb <= "000000";
					when "01000001011111010" => rgb <= "000000";
					when "01000001011111011" => rgb <= "000000";
					when "01000001011111100" => rgb <= "000000";
					when "01000001011111101" => rgb <= "000000";
					when "01000001011111110" => rgb <= "000000";
					when "01000001011111111" => rgb <= "000000";
					when "01000001100000000" => rgb <= "000000";
					when "01000001100000001" => rgb <= "000000";
					when "01000001100000010" => rgb <= "000000";
					when "01000001100000011" => rgb <= "000000";
					when "01000001100000100" => rgb <= "000000";
					when "01000001100000101" => rgb <= "000000";
					when "01000001100000110" => rgb <= "000000";
					when "01000001100000111" => rgb <= "000000";
					when "01000001100001000" => rgb <= "000000";
					when "01000001100001001" => rgb <= "000000";
					when "01000001100001010" => rgb <= "000000";
					when "01000001100001011" => rgb <= "000000";
					when "01000001100001100" => rgb <= "000000";
					when "01000001100001101" => rgb <= "000000";
					when "01000001100001110" => rgb <= "000000";
					when "01000001100001111" => rgb <= "000000";
					when "01000001100010000" => rgb <= "000000";
					when "01000001100010001" => rgb <= "000000";
					when "01000001100010010" => rgb <= "000000";
					when "01000001100010011" => rgb <= "000000";
					when "01000001100010100" => rgb <= "000000";
					when "01000001100010101" => rgb <= "000000";
					when "01000001100010110" => rgb <= "000000";
					when "01000001100010111" => rgb <= "000000";
					when "01000001100011000" => rgb <= "000000";
					when "01000001100011001" => rgb <= "000000";
					when "01000001100011010" => rgb <= "000000";
					when "01000001100011011" => rgb <= "000000";
					when "01000001100011100" => rgb <= "000000";
					when "01000001100011101" => rgb <= "000000";
					when "01000001100011110" => rgb <= "000000";
					when "01000001100011111" => rgb <= "000000";
					when "01000001100100000" => rgb <= "000000";
					when "01000001100100001" => rgb <= "000000";
					when "01000001100100010" => rgb <= "000000";
					when "01000001100100011" => rgb <= "000000";
					when "01000001100100100" => rgb <= "000000";
					when "01000001100100101" => rgb <= "000000";
					when "01000001100100110" => rgb <= "000000";
					when "01000001100100111" => rgb <= "000000";
					when "01000001100101000" => rgb <= "000000";
					when "01000001100101001" => rgb <= "000000";
					when "01000001100101010" => rgb <= "000000";
					when "01000001100101011" => rgb <= "000000";
					when "01000001100101100" => rgb <= "000000";
					when "01000001100101101" => rgb <= "000000";
					when "01000001100101110" => rgb <= "000000";
					when "01000001100101111" => rgb <= "000000";
					when "01000001100110000" => rgb <= "000000";
					when "01000001100110001" => rgb <= "000000";
					when "01000001100110010" => rgb <= "000000";
					when "01000001100110011" => rgb <= "000000";
					when "01000001100110100" => rgb <= "000000";
					when "01000001100110101" => rgb <= "000000";
					when "01000001100110110" => rgb <= "000000";
					when "01000001100110111" => rgb <= "000000";
					when "01000001100111000" => rgb <= "000000";
					when "01000001100111001" => rgb <= "000000";
					when "01000001100111010" => rgb <= "000000";
					when "01000001100111011" => rgb <= "000000";
					when "01000001100111100" => rgb <= "000000";
					when "01000001100111101" => rgb <= "000000";
					when "01000001100111110" => rgb <= "000000";
					when "01000001100111111" => rgb <= "000000";
					when "01000010000000000" => rgb <= "000000";
					when "01000010000000001" => rgb <= "000000";
					when "01000010000000010" => rgb <= "000000";
					when "01000010000000011" => rgb <= "000000";
					when "01000010000000100" => rgb <= "000000";
					when "01000010000000101" => rgb <= "000000";
					when "01000010000000110" => rgb <= "000000";
					when "01000010000000111" => rgb <= "000000";
					when "01000010000001000" => rgb <= "000000";
					when "01000010000001001" => rgb <= "000000";
					when "01000010000001010" => rgb <= "000000";
					when "01000010000001011" => rgb <= "000000";
					when "01000010000001100" => rgb <= "000000";
					when "01000010000001101" => rgb <= "000000";
					when "01000010000001110" => rgb <= "000000";
					when "01000010000001111" => rgb <= "000000";
					when "01000010000010000" => rgb <= "000000";
					when "01000010000010001" => rgb <= "000000";
					when "01000010000010010" => rgb <= "000000";
					when "01000010000010011" => rgb <= "000000";
					when "01000010000010100" => rgb <= "000000";
					when "01000010000010101" => rgb <= "000000";
					when "01000010000010110" => rgb <= "000000";
					when "01000010000010111" => rgb <= "000000";
					when "01000010000011000" => rgb <= "000000";
					when "01000010000011001" => rgb <= "000000";
					when "01000010000011010" => rgb <= "000000";
					when "01000010000011011" => rgb <= "000000";
					when "01000010000011100" => rgb <= "000000";
					when "01000010000011101" => rgb <= "000000";
					when "01000010000011110" => rgb <= "000000";
					when "01000010000011111" => rgb <= "000000";
					when "01000010000100000" => rgb <= "000000";
					when "01000010000100001" => rgb <= "000000";
					when "01000010000100010" => rgb <= "000000";
					when "01000010000100011" => rgb <= "000000";
					when "01000010000100100" => rgb <= "000000";
					when "01000010000100101" => rgb <= "000000";
					when "01000010000100110" => rgb <= "000000";
					when "01000010000100111" => rgb <= "000000";
					when "01000010000101000" => rgb <= "000000";
					when "01000010000101001" => rgb <= "000000";
					when "01000010000101010" => rgb <= "000000";
					when "01000010000101011" => rgb <= "000000";
					when "01000010000101100" => rgb <= "000000";
					when "01000010000101101" => rgb <= "000000";
					when "01000010000101110" => rgb <= "000000";
					when "01000010000101111" => rgb <= "000000";
					when "01000010000110000" => rgb <= "000000";
					when "01000010000110001" => rgb <= "000000";
					when "01000010000110010" => rgb <= "000000";
					when "01000010000110011" => rgb <= "000000";
					when "01000010000110100" => rgb <= "000000";
					when "01000010000110101" => rgb <= "000000";
					when "01000010000110110" => rgb <= "000000";
					when "01000010000110111" => rgb <= "000000";
					when "01000010000111000" => rgb <= "000000";
					when "01000010000111001" => rgb <= "000000";
					when "01000010000111010" => rgb <= "000000";
					when "01000010000111011" => rgb <= "000000";
					when "01000010000111100" => rgb <= "000000";
					when "01000010000111101" => rgb <= "000000";
					when "01000010000111110" => rgb <= "000000";
					when "01000010000111111" => rgb <= "000000";
					when "01000010001000000" => rgb <= "000000";
					when "01000010001000001" => rgb <= "000000";
					when "01000010001000010" => rgb <= "000000";
					when "01000010001000011" => rgb <= "000000";
					when "01000010001000100" => rgb <= "000000";
					when "01000010001000101" => rgb <= "000000";
					when "01000010001000110" => rgb <= "000000";
					when "01000010001000111" => rgb <= "000000";
					when "01000010001001000" => rgb <= "000000";
					when "01000010001001001" => rgb <= "000000";
					when "01000010001001010" => rgb <= "000000";
					when "01000010001001011" => rgb <= "000000";
					when "01000010001001100" => rgb <= "000000";
					when "01000010001001101" => rgb <= "000000";
					when "01000010001001110" => rgb <= "000000";
					when "01000010001001111" => rgb <= "000000";
					when "01000010001010000" => rgb <= "000000";
					when "01000010001010001" => rgb <= "000000";
					when "01000010001010010" => rgb <= "000000";
					when "01000010001010011" => rgb <= "000000";
					when "01000010001010100" => rgb <= "000000";
					when "01000010001010101" => rgb <= "000000";
					when "01000010001010110" => rgb <= "000000";
					when "01000010001010111" => rgb <= "000000";
					when "01000010001011000" => rgb <= "000000";
					when "01000010001011001" => rgb <= "000000";
					when "01000010001011010" => rgb <= "000000";
					when "01000010001011011" => rgb <= "000000";
					when "01000010001011100" => rgb <= "000000";
					when "01000010001011101" => rgb <= "000000";
					when "01000010001011110" => rgb <= "000000";
					when "01000010001011111" => rgb <= "000000";
					when "01000010001100000" => rgb <= "000000";
					when "01000010001100001" => rgb <= "000000";
					when "01000010001100010" => rgb <= "000000";
					when "01000010001100011" => rgb <= "000000";
					when "01000010001100100" => rgb <= "000000";
					when "01000010001100101" => rgb <= "000000";
					when "01000010001100110" => rgb <= "000000";
					when "01000010001100111" => rgb <= "000000";
					when "01000010001101000" => rgb <= "000000";
					when "01000010001101001" => rgb <= "000000";
					when "01000010001101010" => rgb <= "000000";
					when "01000010001101011" => rgb <= "000000";
					when "01000010001101100" => rgb <= "000000";
					when "01000010001101101" => rgb <= "000000";
					when "01000010001101110" => rgb <= "000000";
					when "01000010001101111" => rgb <= "000000";
					when "01000010001110000" => rgb <= "000000";
					when "01000010001110001" => rgb <= "010000";
					when "01000010001110010" => rgb <= "101000";
					when "01000010001110011" => rgb <= "101000";
					when "01000010001110100" => rgb <= "101000";
					when "01000010001110101" => rgb <= "101000";
					when "01000010001110110" => rgb <= "101000";
					when "01000010001110111" => rgb <= "101000";
					when "01000010001111000" => rgb <= "101000";
					when "01000010001111001" => rgb <= "101000";
					when "01000010001111010" => rgb <= "101000";
					when "01000010001111011" => rgb <= "101000";
					when "01000010001111100" => rgb <= "101000";
					when "01000010001111101" => rgb <= "101000";
					when "01000010001111110" => rgb <= "101000";
					when "01000010001111111" => rgb <= "101000";
					when "01000010010000000" => rgb <= "101000";
					when "01000010010000001" => rgb <= "101000";
					when "01000010010000010" => rgb <= "101000";
					when "01000010010000011" => rgb <= "101000";
					when "01000010010000100" => rgb <= "101000";
					when "01000010010000101" => rgb <= "101000";
					when "01000010010000110" => rgb <= "101000";
					when "01000010010000111" => rgb <= "101000";
					when "01000010010001000" => rgb <= "101000";
					when "01000010010001001" => rgb <= "101000";
					when "01000010010001010" => rgb <= "101000";
					when "01000010010001011" => rgb <= "101000";
					when "01000010010001100" => rgb <= "101000";
					when "01000010010001101" => rgb <= "101000";
					when "01000010010001110" => rgb <= "101000";
					when "01000010010001111" => rgb <= "101000";
					when "01000010010010000" => rgb <= "101000";
					when "01000010010010001" => rgb <= "101000";
					when "01000010010010010" => rgb <= "101000";
					when "01000010010010011" => rgb <= "101000";
					when "01000010010010100" => rgb <= "101000";
					when "01000010010010101" => rgb <= "101000";
					when "01000010010010110" => rgb <= "101000";
					when "01000010010010111" => rgb <= "101000";
					when "01000010010011000" => rgb <= "101000";
					when "01000010010011001" => rgb <= "101000";
					when "01000010010011010" => rgb <= "101000";
					when "01000010010011011" => rgb <= "101000";
					when "01000010010011100" => rgb <= "101000";
					when "01000010010011101" => rgb <= "101000";
					when "01000010010011110" => rgb <= "101000";
					when "01000010010011111" => rgb <= "101000";
					when "01000010010100000" => rgb <= "101000";
					when "01000010010100001" => rgb <= "101000";
					when "01000010010100010" => rgb <= "101000";
					when "01000010010100011" => rgb <= "101000";
					when "01000010010100100" => rgb <= "101000";
					when "01000010010100101" => rgb <= "101000";
					when "01000010010100110" => rgb <= "101000";
					when "01000010010100111" => rgb <= "101000";
					when "01000010010101000" => rgb <= "101000";
					when "01000010010101001" => rgb <= "101000";
					when "01000010010101010" => rgb <= "101000";
					when "01000010010101011" => rgb <= "101000";
					when "01000010010101100" => rgb <= "101000";
					when "01000010010101101" => rgb <= "101000";
					when "01000010010101110" => rgb <= "101000";
					when "01000010010101111" => rgb <= "101000";
					when "01000010010110000" => rgb <= "101000";
					when "01000010010110001" => rgb <= "101000";
					when "01000010010110010" => rgb <= "101000";
					when "01000010010110011" => rgb <= "101000";
					when "01000010010110100" => rgb <= "101000";
					when "01000010010110101" => rgb <= "101000";
					when "01000010010110110" => rgb <= "101000";
					when "01000010010110111" => rgb <= "101000";
					when "01000010010111000" => rgb <= "101000";
					when "01000010010111001" => rgb <= "101000";
					when "01000010010111010" => rgb <= "101000";
					when "01000010010111011" => rgb <= "101000";
					when "01000010010111100" => rgb <= "101000";
					when "01000010010111101" => rgb <= "101000";
					when "01000010010111110" => rgb <= "101000";
					when "01000010010111111" => rgb <= "101000";
					when "01000010011000000" => rgb <= "101000";
					when "01000010011000001" => rgb <= "101000";
					when "01000010011000010" => rgb <= "101000";
					when "01000010011000011" => rgb <= "101000";
					when "01000010011000100" => rgb <= "101000";
					when "01000010011000101" => rgb <= "101000";
					when "01000010011000110" => rgb <= "101000";
					when "01000010011000111" => rgb <= "101000";
					when "01000010011001000" => rgb <= "101000";
					when "01000010011001001" => rgb <= "101000";
					when "01000010011001010" => rgb <= "101000";
					when "01000010011001011" => rgb <= "101000";
					when "01000010011001100" => rgb <= "000000";
					when "01000010011001101" => rgb <= "000000";
					when "01000010011001110" => rgb <= "000000";
					when "01000010011001111" => rgb <= "000000";
					when "01000010011010000" => rgb <= "000000";
					when "01000010011010001" => rgb <= "000000";
					when "01000010011010010" => rgb <= "000000";
					when "01000010011010011" => rgb <= "000000";
					when "01000010011010100" => rgb <= "000000";
					when "01000010011010101" => rgb <= "000000";
					when "01000010011010110" => rgb <= "000000";
					when "01000010011010111" => rgb <= "000000";
					when "01000010011011000" => rgb <= "000000";
					when "01000010011011001" => rgb <= "000000";
					when "01000010011011010" => rgb <= "000000";
					when "01000010011011011" => rgb <= "000000";
					when "01000010011011100" => rgb <= "000000";
					when "01000010011011101" => rgb <= "000000";
					when "01000010011011110" => rgb <= "000000";
					when "01000010011011111" => rgb <= "000000";
					when "01000010011100000" => rgb <= "000000";
					when "01000010011100001" => rgb <= "000000";
					when "01000010011100010" => rgb <= "000000";
					when "01000010011100011" => rgb <= "000000";
					when "01000010011100100" => rgb <= "000000";
					when "01000010011100101" => rgb <= "000000";
					when "01000010011100110" => rgb <= "000000";
					when "01000010011100111" => rgb <= "000000";
					when "01000010011101000" => rgb <= "000000";
					when "01000010011101001" => rgb <= "000000";
					when "01000010011101010" => rgb <= "000000";
					when "01000010011101011" => rgb <= "000000";
					when "01000010011101100" => rgb <= "000000";
					when "01000010011101101" => rgb <= "000000";
					when "01000010011101110" => rgb <= "000000";
					when "01000010011101111" => rgb <= "000000";
					when "01000010011110000" => rgb <= "000000";
					when "01000010011110001" => rgb <= "000000";
					when "01000010011110010" => rgb <= "000000";
					when "01000010011110011" => rgb <= "000000";
					when "01000010011110100" => rgb <= "000000";
					when "01000010011110101" => rgb <= "000000";
					when "01000010011110110" => rgb <= "000000";
					when "01000010011110111" => rgb <= "000000";
					when "01000010011111000" => rgb <= "000000";
					when "01000010011111001" => rgb <= "000000";
					when "01000010011111010" => rgb <= "000000";
					when "01000010011111011" => rgb <= "000000";
					when "01000010011111100" => rgb <= "000000";
					when "01000010011111101" => rgb <= "000000";
					when "01000010011111110" => rgb <= "000000";
					when "01000010011111111" => rgb <= "000000";
					when "01000010100000000" => rgb <= "000000";
					when "01000010100000001" => rgb <= "000000";
					when "01000010100000010" => rgb <= "000000";
					when "01000010100000011" => rgb <= "000000";
					when "01000010100000100" => rgb <= "000000";
					when "01000010100000101" => rgb <= "000000";
					when "01000010100000110" => rgb <= "000000";
					when "01000010100000111" => rgb <= "000000";
					when "01000010100001000" => rgb <= "000000";
					when "01000010100001001" => rgb <= "000000";
					when "01000010100001010" => rgb <= "000000";
					when "01000010100001011" => rgb <= "000000";
					when "01000010100001100" => rgb <= "000000";
					when "01000010100001101" => rgb <= "000000";
					when "01000010100001110" => rgb <= "000000";
					when "01000010100001111" => rgb <= "000000";
					when "01000010100010000" => rgb <= "000000";
					when "01000010100010001" => rgb <= "000000";
					when "01000010100010010" => rgb <= "000000";
					when "01000010100010011" => rgb <= "000000";
					when "01000010100010100" => rgb <= "000000";
					when "01000010100010101" => rgb <= "000000";
					when "01000010100010110" => rgb <= "000000";
					when "01000010100010111" => rgb <= "000000";
					when "01000010100011000" => rgb <= "000000";
					when "01000010100011001" => rgb <= "000000";
					when "01000010100011010" => rgb <= "000000";
					when "01000010100011011" => rgb <= "000000";
					when "01000010100011100" => rgb <= "000000";
					when "01000010100011101" => rgb <= "000000";
					when "01000010100011110" => rgb <= "000000";
					when "01000010100011111" => rgb <= "000000";
					when "01000010100100000" => rgb <= "000000";
					when "01000010100100001" => rgb <= "000000";
					when "01000010100100010" => rgb <= "000000";
					when "01000010100100011" => rgb <= "000000";
					when "01000010100100100" => rgb <= "000000";
					when "01000010100100101" => rgb <= "000000";
					when "01000010100100110" => rgb <= "000000";
					when "01000010100100111" => rgb <= "000000";
					when "01000010100101000" => rgb <= "000000";
					when "01000010100101001" => rgb <= "000000";
					when "01000010100101010" => rgb <= "000000";
					when "01000010100101011" => rgb <= "000000";
					when "01000010100101100" => rgb <= "000000";
					when "01000010100101101" => rgb <= "000000";
					when "01000010100101110" => rgb <= "000000";
					when "01000010100101111" => rgb <= "000000";
					when "01000010100110000" => rgb <= "000000";
					when "01000010100110001" => rgb <= "000000";
					when "01000010100110010" => rgb <= "000000";
					when "01000010100110011" => rgb <= "000000";
					when "01000010100110100" => rgb <= "000000";
					when "01000010100110101" => rgb <= "000000";
					when "01000010100110110" => rgb <= "000000";
					when "01000010100110111" => rgb <= "000000";
					when "01000010100111000" => rgb <= "000000";
					when "01000010100111001" => rgb <= "000000";
					when "01000010100111010" => rgb <= "000000";
					when "01000010100111011" => rgb <= "000000";
					when "01000010100111100" => rgb <= "000000";
					when "01000010100111101" => rgb <= "000000";
					when "01000010100111110" => rgb <= "000000";
					when "01000010100111111" => rgb <= "000000";
					when "01000011000000000" => rgb <= "000000";
					when "01000011000000001" => rgb <= "000000";
					when "01000011000000010" => rgb <= "000000";
					when "01000011000000011" => rgb <= "000000";
					when "01000011000000100" => rgb <= "000000";
					when "01000011000000101" => rgb <= "000000";
					when "01000011000000110" => rgb <= "000000";
					when "01000011000000111" => rgb <= "000000";
					when "01000011000001000" => rgb <= "000000";
					when "01000011000001001" => rgb <= "000000";
					when "01000011000001010" => rgb <= "000000";
					when "01000011000001011" => rgb <= "000000";
					when "01000011000001100" => rgb <= "000000";
					when "01000011000001101" => rgb <= "000000";
					when "01000011000001110" => rgb <= "000000";
					when "01000011000001111" => rgb <= "000000";
					when "01000011000010000" => rgb <= "000000";
					when "01000011000010001" => rgb <= "000000";
					when "01000011000010010" => rgb <= "000000";
					when "01000011000010011" => rgb <= "000000";
					when "01000011000010100" => rgb <= "000000";
					when "01000011000010101" => rgb <= "000000";
					when "01000011000010110" => rgb <= "000000";
					when "01000011000010111" => rgb <= "000000";
					when "01000011000011000" => rgb <= "000000";
					when "01000011000011001" => rgb <= "000000";
					when "01000011000011010" => rgb <= "000000";
					when "01000011000011011" => rgb <= "000000";
					when "01000011000011100" => rgb <= "000000";
					when "01000011000011101" => rgb <= "000000";
					when "01000011000011110" => rgb <= "000000";
					when "01000011000011111" => rgb <= "000000";
					when "01000011000100000" => rgb <= "000000";
					when "01000011000100001" => rgb <= "000000";
					when "01000011000100010" => rgb <= "000000";
					when "01000011000100011" => rgb <= "000000";
					when "01000011000100100" => rgb <= "000000";
					when "01000011000100101" => rgb <= "000000";
					when "01000011000100110" => rgb <= "000000";
					when "01000011000100111" => rgb <= "000000";
					when "01000011000101000" => rgb <= "000000";
					when "01000011000101001" => rgb <= "000000";
					when "01000011000101010" => rgb <= "000000";
					when "01000011000101011" => rgb <= "000000";
					when "01000011000101100" => rgb <= "000000";
					when "01000011000101101" => rgb <= "000000";
					when "01000011000101110" => rgb <= "000000";
					when "01000011000101111" => rgb <= "000000";
					when "01000011000110000" => rgb <= "000000";
					when "01000011000110001" => rgb <= "000000";
					when "01000011000110010" => rgb <= "000000";
					when "01000011000110011" => rgb <= "000000";
					when "01000011000110100" => rgb <= "000000";
					when "01000011000110101" => rgb <= "000000";
					when "01000011000110110" => rgb <= "000000";
					when "01000011000110111" => rgb <= "000000";
					when "01000011000111000" => rgb <= "000000";
					when "01000011000111001" => rgb <= "000000";
					when "01000011000111010" => rgb <= "000000";
					when "01000011000111011" => rgb <= "000000";
					when "01000011000111100" => rgb <= "000000";
					when "01000011000111101" => rgb <= "000000";
					when "01000011000111110" => rgb <= "000000";
					when "01000011000111111" => rgb <= "000000";
					when "01000011001000000" => rgb <= "000000";
					when "01000011001000001" => rgb <= "000000";
					when "01000011001000010" => rgb <= "000000";
					when "01000011001000011" => rgb <= "000000";
					when "01000011001000100" => rgb <= "000000";
					when "01000011001000101" => rgb <= "000000";
					when "01000011001000110" => rgb <= "000000";
					when "01000011001000111" => rgb <= "000000";
					when "01000011001001000" => rgb <= "000000";
					when "01000011001001001" => rgb <= "000000";
					when "01000011001001010" => rgb <= "000000";
					when "01000011001001011" => rgb <= "000000";
					when "01000011001001100" => rgb <= "000000";
					when "01000011001001101" => rgb <= "000000";
					when "01000011001001110" => rgb <= "000000";
					when "01000011001001111" => rgb <= "000000";
					when "01000011001010000" => rgb <= "000000";
					when "01000011001010001" => rgb <= "000000";
					when "01000011001010010" => rgb <= "000000";
					when "01000011001010011" => rgb <= "000000";
					when "01000011001010100" => rgb <= "000000";
					when "01000011001010101" => rgb <= "000000";
					when "01000011001010110" => rgb <= "000000";
					when "01000011001010111" => rgb <= "000000";
					when "01000011001011000" => rgb <= "000000";
					when "01000011001011001" => rgb <= "000000";
					when "01000011001011010" => rgb <= "000000";
					when "01000011001011011" => rgb <= "000000";
					when "01000011001011100" => rgb <= "000000";
					when "01000011001011101" => rgb <= "000000";
					when "01000011001011110" => rgb <= "000000";
					when "01000011001011111" => rgb <= "000000";
					when "01000011001100000" => rgb <= "000000";
					when "01000011001100001" => rgb <= "000000";
					when "01000011001100010" => rgb <= "000000";
					when "01000011001100011" => rgb <= "000000";
					when "01000011001100100" => rgb <= "000000";
					when "01000011001100101" => rgb <= "000000";
					when "01000011001100110" => rgb <= "000000";
					when "01000011001100111" => rgb <= "000000";
					when "01000011001101000" => rgb <= "000000";
					when "01000011001101001" => rgb <= "000000";
					when "01000011001101010" => rgb <= "000000";
					when "01000011001101011" => rgb <= "000000";
					when "01000011001101100" => rgb <= "000000";
					when "01000011001101101" => rgb <= "000000";
					when "01000011001101110" => rgb <= "000000";
					when "01000011001101111" => rgb <= "000000";
					when "01000011001110000" => rgb <= "000000";
					when "01000011001110001" => rgb <= "010000";
					when "01000011001110010" => rgb <= "101000";
					when "01000011001110011" => rgb <= "101000";
					when "01000011001110100" => rgb <= "101000";
					when "01000011001110101" => rgb <= "101000";
					when "01000011001110110" => rgb <= "101000";
					when "01000011001110111" => rgb <= "101000";
					when "01000011001111000" => rgb <= "101000";
					when "01000011001111001" => rgb <= "101000";
					when "01000011001111010" => rgb <= "101000";
					when "01000011001111011" => rgb <= "101000";
					when "01000011001111100" => rgb <= "101000";
					when "01000011001111101" => rgb <= "101000";
					when "01000011001111110" => rgb <= "101000";
					when "01000011001111111" => rgb <= "101000";
					when "01000011010000000" => rgb <= "101000";
					when "01000011010000001" => rgb <= "101000";
					when "01000011010000010" => rgb <= "101000";
					when "01000011010000011" => rgb <= "101000";
					when "01000011010000100" => rgb <= "101000";
					when "01000011010000101" => rgb <= "101000";
					when "01000011010000110" => rgb <= "101000";
					when "01000011010000111" => rgb <= "101000";
					when "01000011010001000" => rgb <= "101000";
					when "01000011010001001" => rgb <= "101000";
					when "01000011010001010" => rgb <= "101000";
					when "01000011010001011" => rgb <= "101000";
					when "01000011010001100" => rgb <= "101000";
					when "01000011010001101" => rgb <= "101000";
					when "01000011010001110" => rgb <= "101000";
					when "01000011010001111" => rgb <= "101000";
					when "01000011010010000" => rgb <= "101000";
					when "01000011010010001" => rgb <= "101000";
					when "01000011010010010" => rgb <= "101000";
					when "01000011010010011" => rgb <= "101000";
					when "01000011010010100" => rgb <= "101000";
					when "01000011010010101" => rgb <= "101000";
					when "01000011010010110" => rgb <= "101000";
					when "01000011010010111" => rgb <= "101000";
					when "01000011010011000" => rgb <= "101000";
					when "01000011010011001" => rgb <= "101000";
					when "01000011010011010" => rgb <= "101000";
					when "01000011010011011" => rgb <= "101000";
					when "01000011010011100" => rgb <= "101000";
					when "01000011010011101" => rgb <= "101000";
					when "01000011010011110" => rgb <= "101000";
					when "01000011010011111" => rgb <= "101000";
					when "01000011010100000" => rgb <= "101000";
					when "01000011010100001" => rgb <= "101000";
					when "01000011010100010" => rgb <= "101000";
					when "01000011010100011" => rgb <= "101000";
					when "01000011010100100" => rgb <= "101000";
					when "01000011010100101" => rgb <= "101000";
					when "01000011010100110" => rgb <= "101000";
					when "01000011010100111" => rgb <= "101000";
					when "01000011010101000" => rgb <= "101000";
					when "01000011010101001" => rgb <= "101000";
					when "01000011010101010" => rgb <= "101000";
					when "01000011010101011" => rgb <= "101000";
					when "01000011010101100" => rgb <= "101000";
					when "01000011010101101" => rgb <= "101000";
					when "01000011010101110" => rgb <= "101000";
					when "01000011010101111" => rgb <= "101000";
					when "01000011010110000" => rgb <= "101000";
					when "01000011010110001" => rgb <= "101000";
					when "01000011010110010" => rgb <= "101000";
					when "01000011010110011" => rgb <= "101000";
					when "01000011010110100" => rgb <= "101000";
					when "01000011010110101" => rgb <= "101000";
					when "01000011010110110" => rgb <= "101000";
					when "01000011010110111" => rgb <= "101000";
					when "01000011010111000" => rgb <= "101000";
					when "01000011010111001" => rgb <= "101000";
					when "01000011010111010" => rgb <= "101000";
					when "01000011010111011" => rgb <= "101000";
					when "01000011010111100" => rgb <= "101000";
					when "01000011010111101" => rgb <= "101000";
					when "01000011010111110" => rgb <= "101000";
					when "01000011010111111" => rgb <= "101000";
					when "01000011011000000" => rgb <= "101000";
					when "01000011011000001" => rgb <= "101000";
					when "01000011011000010" => rgb <= "101000";
					when "01000011011000011" => rgb <= "101000";
					when "01000011011000100" => rgb <= "101000";
					when "01000011011000101" => rgb <= "101000";
					when "01000011011000110" => rgb <= "101000";
					when "01000011011000111" => rgb <= "101000";
					when "01000011011001000" => rgb <= "101000";
					when "01000011011001001" => rgb <= "101000";
					when "01000011011001010" => rgb <= "101000";
					when "01000011011001011" => rgb <= "101000";
					when "01000011011001100" => rgb <= "000000";
					when "01000011011001101" => rgb <= "000000";
					when "01000011011001110" => rgb <= "000000";
					when "01000011011001111" => rgb <= "000000";
					when "01000011011010000" => rgb <= "000000";
					when "01000011011010001" => rgb <= "000000";
					when "01000011011010010" => rgb <= "000000";
					when "01000011011010011" => rgb <= "000000";
					when "01000011011010100" => rgb <= "000000";
					when "01000011011010101" => rgb <= "000000";
					when "01000011011010110" => rgb <= "000000";
					when "01000011011010111" => rgb <= "000000";
					when "01000011011011000" => rgb <= "000000";
					when "01000011011011001" => rgb <= "000000";
					when "01000011011011010" => rgb <= "000000";
					when "01000011011011011" => rgb <= "000000";
					when "01000011011011100" => rgb <= "000000";
					when "01000011011011101" => rgb <= "000000";
					when "01000011011011110" => rgb <= "000000";
					when "01000011011011111" => rgb <= "000000";
					when "01000011011100000" => rgb <= "000000";
					when "01000011011100001" => rgb <= "000000";
					when "01000011011100010" => rgb <= "000000";
					when "01000011011100011" => rgb <= "000000";
					when "01000011011100100" => rgb <= "000000";
					when "01000011011100101" => rgb <= "000000";
					when "01000011011100110" => rgb <= "000000";
					when "01000011011100111" => rgb <= "000000";
					when "01000011011101000" => rgb <= "000000";
					when "01000011011101001" => rgb <= "000000";
					when "01000011011101010" => rgb <= "000000";
					when "01000011011101011" => rgb <= "000000";
					when "01000011011101100" => rgb <= "000000";
					when "01000011011101101" => rgb <= "000000";
					when "01000011011101110" => rgb <= "000000";
					when "01000011011101111" => rgb <= "000000";
					when "01000011011110000" => rgb <= "000000";
					when "01000011011110001" => rgb <= "000000";
					when "01000011011110010" => rgb <= "000000";
					when "01000011011110011" => rgb <= "000000";
					when "01000011011110100" => rgb <= "000000";
					when "01000011011110101" => rgb <= "000000";
					when "01000011011110110" => rgb <= "000000";
					when "01000011011110111" => rgb <= "000000";
					when "01000011011111000" => rgb <= "000000";
					when "01000011011111001" => rgb <= "000000";
					when "01000011011111010" => rgb <= "000000";
					when "01000011011111011" => rgb <= "000000";
					when "01000011011111100" => rgb <= "000000";
					when "01000011011111101" => rgb <= "000000";
					when "01000011011111110" => rgb <= "000000";
					when "01000011011111111" => rgb <= "000000";
					when "01000011100000000" => rgb <= "000000";
					when "01000011100000001" => rgb <= "000000";
					when "01000011100000010" => rgb <= "000000";
					when "01000011100000011" => rgb <= "000000";
					when "01000011100000100" => rgb <= "000000";
					when "01000011100000101" => rgb <= "000000";
					when "01000011100000110" => rgb <= "000000";
					when "01000011100000111" => rgb <= "000000";
					when "01000011100001000" => rgb <= "000000";
					when "01000011100001001" => rgb <= "000000";
					when "01000011100001010" => rgb <= "000000";
					when "01000011100001011" => rgb <= "000000";
					when "01000011100001100" => rgb <= "000000";
					when "01000011100001101" => rgb <= "000000";
					when "01000011100001110" => rgb <= "000000";
					when "01000011100001111" => rgb <= "000000";
					when "01000011100010000" => rgb <= "000000";
					when "01000011100010001" => rgb <= "000000";
					when "01000011100010010" => rgb <= "000000";
					when "01000011100010011" => rgb <= "000000";
					when "01000011100010100" => rgb <= "000000";
					when "01000011100010101" => rgb <= "000000";
					when "01000011100010110" => rgb <= "000000";
					when "01000011100010111" => rgb <= "000000";
					when "01000011100011000" => rgb <= "000000";
					when "01000011100011001" => rgb <= "000000";
					when "01000011100011010" => rgb <= "000000";
					when "01000011100011011" => rgb <= "000000";
					when "01000011100011100" => rgb <= "000000";
					when "01000011100011101" => rgb <= "000000";
					when "01000011100011110" => rgb <= "000000";
					when "01000011100011111" => rgb <= "000000";
					when "01000011100100000" => rgb <= "000000";
					when "01000011100100001" => rgb <= "000000";
					when "01000011100100010" => rgb <= "000000";
					when "01000011100100011" => rgb <= "000000";
					when "01000011100100100" => rgb <= "000000";
					when "01000011100100101" => rgb <= "000000";
					when "01000011100100110" => rgb <= "000000";
					when "01000011100100111" => rgb <= "000000";
					when "01000011100101000" => rgb <= "000000";
					when "01000011100101001" => rgb <= "000000";
					when "01000011100101010" => rgb <= "000000";
					when "01000011100101011" => rgb <= "000000";
					when "01000011100101100" => rgb <= "000000";
					when "01000011100101101" => rgb <= "000000";
					when "01000011100101110" => rgb <= "000000";
					when "01000011100101111" => rgb <= "000000";
					when "01000011100110000" => rgb <= "000000";
					when "01000011100110001" => rgb <= "000000";
					when "01000011100110010" => rgb <= "000000";
					when "01000011100110011" => rgb <= "000000";
					when "01000011100110100" => rgb <= "000000";
					when "01000011100110101" => rgb <= "000000";
					when "01000011100110110" => rgb <= "000000";
					when "01000011100110111" => rgb <= "000000";
					when "01000011100111000" => rgb <= "000000";
					when "01000011100111001" => rgb <= "000000";
					when "01000011100111010" => rgb <= "000000";
					when "01000011100111011" => rgb <= "000000";
					when "01000011100111100" => rgb <= "000000";
					when "01000011100111101" => rgb <= "000000";
					when "01000011100111110" => rgb <= "000000";
					when "01000011100111111" => rgb <= "000000";
					when "01000100000000000" => rgb <= "000000";
					when "01000100000000001" => rgb <= "000000";
					when "01000100000000010" => rgb <= "000000";
					when "01000100000000011" => rgb <= "000000";
					when "01000100000000100" => rgb <= "000000";
					when "01000100000000101" => rgb <= "000000";
					when "01000100000000110" => rgb <= "000000";
					when "01000100000000111" => rgb <= "000000";
					when "01000100000001000" => rgb <= "000000";
					when "01000100000001001" => rgb <= "000000";
					when "01000100000001010" => rgb <= "000000";
					when "01000100000001011" => rgb <= "000000";
					when "01000100000001100" => rgb <= "000000";
					when "01000100000001101" => rgb <= "000000";
					when "01000100000001110" => rgb <= "000000";
					when "01000100000001111" => rgb <= "000000";
					when "01000100000010000" => rgb <= "000000";
					when "01000100000010001" => rgb <= "000000";
					when "01000100000010010" => rgb <= "000000";
					when "01000100000010011" => rgb <= "000000";
					when "01000100000010100" => rgb <= "000000";
					when "01000100000010101" => rgb <= "000000";
					when "01000100000010110" => rgb <= "000000";
					when "01000100000010111" => rgb <= "000000";
					when "01000100000011000" => rgb <= "000000";
					when "01000100000011001" => rgb <= "000000";
					when "01000100000011010" => rgb <= "000000";
					when "01000100000011011" => rgb <= "000000";
					when "01000100000011100" => rgb <= "000000";
					when "01000100000011101" => rgb <= "000000";
					when "01000100000011110" => rgb <= "000000";
					when "01000100000011111" => rgb <= "000000";
					when "01000100000100000" => rgb <= "000000";
					when "01000100000100001" => rgb <= "000000";
					when "01000100000100010" => rgb <= "000000";
					when "01000100000100011" => rgb <= "000000";
					when "01000100000100100" => rgb <= "000000";
					when "01000100000100101" => rgb <= "000000";
					when "01000100000100110" => rgb <= "000000";
					when "01000100000100111" => rgb <= "000000";
					when "01000100000101000" => rgb <= "000000";
					when "01000100000101001" => rgb <= "000000";
					when "01000100000101010" => rgb <= "000000";
					when "01000100000101011" => rgb <= "000000";
					when "01000100000101100" => rgb <= "000000";
					when "01000100000101101" => rgb <= "000000";
					when "01000100000101110" => rgb <= "000000";
					when "01000100000101111" => rgb <= "000000";
					when "01000100000110000" => rgb <= "000000";
					when "01000100000110001" => rgb <= "000000";
					when "01000100000110010" => rgb <= "000000";
					when "01000100000110011" => rgb <= "000000";
					when "01000100000110100" => rgb <= "000000";
					when "01000100000110101" => rgb <= "000000";
					when "01000100000110110" => rgb <= "000000";
					when "01000100000110111" => rgb <= "000000";
					when "01000100000111000" => rgb <= "000000";
					when "01000100000111001" => rgb <= "000000";
					when "01000100000111010" => rgb <= "000000";
					when "01000100000111011" => rgb <= "000000";
					when "01000100000111100" => rgb <= "000000";
					when "01000100000111101" => rgb <= "000000";
					when "01000100000111110" => rgb <= "000000";
					when "01000100000111111" => rgb <= "000000";
					when "01000100001000000" => rgb <= "000000";
					when "01000100001000001" => rgb <= "000000";
					when "01000100001000010" => rgb <= "000000";
					when "01000100001000011" => rgb <= "000000";
					when "01000100001000100" => rgb <= "000000";
					when "01000100001000101" => rgb <= "000000";
					when "01000100001000110" => rgb <= "000000";
					when "01000100001000111" => rgb <= "000000";
					when "01000100001001000" => rgb <= "000000";
					when "01000100001001001" => rgb <= "000000";
					when "01000100001001010" => rgb <= "000000";
					when "01000100001001011" => rgb <= "000000";
					when "01000100001001100" => rgb <= "000000";
					when "01000100001001101" => rgb <= "000000";
					when "01000100001001110" => rgb <= "000000";
					when "01000100001001111" => rgb <= "000000";
					when "01000100001010000" => rgb <= "000000";
					when "01000100001010001" => rgb <= "000000";
					when "01000100001010010" => rgb <= "000000";
					when "01000100001010011" => rgb <= "000000";
					when "01000100001010100" => rgb <= "000000";
					when "01000100001010101" => rgb <= "000000";
					when "01000100001010110" => rgb <= "000000";
					when "01000100001010111" => rgb <= "000000";
					when "01000100001011000" => rgb <= "000000";
					when "01000100001011001" => rgb <= "000000";
					when "01000100001011010" => rgb <= "000000";
					when "01000100001011011" => rgb <= "000000";
					when "01000100001011100" => rgb <= "000000";
					when "01000100001011101" => rgb <= "000000";
					when "01000100001011110" => rgb <= "000000";
					when "01000100001011111" => rgb <= "000000";
					when "01000100001100000" => rgb <= "000000";
					when "01000100001100001" => rgb <= "000000";
					when "01000100001100010" => rgb <= "000000";
					when "01000100001100011" => rgb <= "000000";
					when "01000100001100100" => rgb <= "000000";
					when "01000100001100101" => rgb <= "000000";
					when "01000100001100110" => rgb <= "000000";
					when "01000100001100111" => rgb <= "000000";
					when "01000100001101000" => rgb <= "000000";
					when "01000100001101001" => rgb <= "000000";
					when "01000100001101010" => rgb <= "000000";
					when "01000100001101011" => rgb <= "000000";
					when "01000100001101100" => rgb <= "000000";
					when "01000100001101101" => rgb <= "000000";
					when "01000100001101110" => rgb <= "000000";
					when "01000100001101111" => rgb <= "000000";
					when "01000100001110000" => rgb <= "000000";
					when "01000100001110001" => rgb <= "010000";
					when "01000100001110010" => rgb <= "101000";
					when "01000100001110011" => rgb <= "101000";
					when "01000100001110100" => rgb <= "101000";
					when "01000100001110101" => rgb <= "101000";
					when "01000100001110110" => rgb <= "101000";
					when "01000100001110111" => rgb <= "101000";
					when "01000100001111000" => rgb <= "101000";
					when "01000100001111001" => rgb <= "101000";
					when "01000100001111010" => rgb <= "101000";
					when "01000100001111011" => rgb <= "101000";
					when "01000100001111100" => rgb <= "101000";
					when "01000100001111101" => rgb <= "101000";
					when "01000100001111110" => rgb <= "101000";
					when "01000100001111111" => rgb <= "101000";
					when "01000100010000000" => rgb <= "101000";
					when "01000100010000001" => rgb <= "101000";
					when "01000100010000010" => rgb <= "101000";
					when "01000100010000011" => rgb <= "101000";
					when "01000100010000100" => rgb <= "101000";
					when "01000100010000101" => rgb <= "101000";
					when "01000100010000110" => rgb <= "101000";
					when "01000100010000111" => rgb <= "101000";
					when "01000100010001000" => rgb <= "101000";
					when "01000100010001001" => rgb <= "101000";
					when "01000100010001010" => rgb <= "101000";
					when "01000100010001011" => rgb <= "101000";
					when "01000100010001100" => rgb <= "101000";
					when "01000100010001101" => rgb <= "101000";
					when "01000100010001110" => rgb <= "101000";
					when "01000100010001111" => rgb <= "101000";
					when "01000100010010000" => rgb <= "101000";
					when "01000100010010001" => rgb <= "101000";
					when "01000100010010010" => rgb <= "101000";
					when "01000100010010011" => rgb <= "101000";
					when "01000100010010100" => rgb <= "101000";
					when "01000100010010101" => rgb <= "101000";
					when "01000100010010110" => rgb <= "101000";
					when "01000100010010111" => rgb <= "101000";
					when "01000100010011000" => rgb <= "101000";
					when "01000100010011001" => rgb <= "101000";
					when "01000100010011010" => rgb <= "101000";
					when "01000100010011011" => rgb <= "101000";
					when "01000100010011100" => rgb <= "101000";
					when "01000100010011101" => rgb <= "101000";
					when "01000100010011110" => rgb <= "101000";
					when "01000100010011111" => rgb <= "101000";
					when "01000100010100000" => rgb <= "101000";
					when "01000100010100001" => rgb <= "101000";
					when "01000100010100010" => rgb <= "101000";
					when "01000100010100011" => rgb <= "101000";
					when "01000100010100100" => rgb <= "101000";
					when "01000100010100101" => rgb <= "101000";
					when "01000100010100110" => rgb <= "101000";
					when "01000100010100111" => rgb <= "101000";
					when "01000100010101000" => rgb <= "101000";
					when "01000100010101001" => rgb <= "101000";
					when "01000100010101010" => rgb <= "101000";
					when "01000100010101011" => rgb <= "101000";
					when "01000100010101100" => rgb <= "101000";
					when "01000100010101101" => rgb <= "101000";
					when "01000100010101110" => rgb <= "101000";
					when "01000100010101111" => rgb <= "101000";
					when "01000100010110000" => rgb <= "101000";
					when "01000100010110001" => rgb <= "101000";
					when "01000100010110010" => rgb <= "101000";
					when "01000100010110011" => rgb <= "101000";
					when "01000100010110100" => rgb <= "101000";
					when "01000100010110101" => rgb <= "101000";
					when "01000100010110110" => rgb <= "101000";
					when "01000100010110111" => rgb <= "101000";
					when "01000100010111000" => rgb <= "101000";
					when "01000100010111001" => rgb <= "101000";
					when "01000100010111010" => rgb <= "101000";
					when "01000100010111011" => rgb <= "101000";
					when "01000100010111100" => rgb <= "101000";
					when "01000100010111101" => rgb <= "101000";
					when "01000100010111110" => rgb <= "101000";
					when "01000100010111111" => rgb <= "101000";
					when "01000100011000000" => rgb <= "101000";
					when "01000100011000001" => rgb <= "101000";
					when "01000100011000010" => rgb <= "101000";
					when "01000100011000011" => rgb <= "101000";
					when "01000100011000100" => rgb <= "101000";
					when "01000100011000101" => rgb <= "101000";
					when "01000100011000110" => rgb <= "101000";
					when "01000100011000111" => rgb <= "101000";
					when "01000100011001000" => rgb <= "101000";
					when "01000100011001001" => rgb <= "101000";
					when "01000100011001010" => rgb <= "101000";
					when "01000100011001011" => rgb <= "101000";
					when "01000100011001100" => rgb <= "000000";
					when "01000100011001101" => rgb <= "000000";
					when "01000100011001110" => rgb <= "000000";
					when "01000100011001111" => rgb <= "000000";
					when "01000100011010000" => rgb <= "000000";
					when "01000100011010001" => rgb <= "000000";
					when "01000100011010010" => rgb <= "000000";
					when "01000100011010011" => rgb <= "000000";
					when "01000100011010100" => rgb <= "000000";
					when "01000100011010101" => rgb <= "000000";
					when "01000100011010110" => rgb <= "000000";
					when "01000100011010111" => rgb <= "000000";
					when "01000100011011000" => rgb <= "000000";
					when "01000100011011001" => rgb <= "000000";
					when "01000100011011010" => rgb <= "000000";
					when "01000100011011011" => rgb <= "000000";
					when "01000100011011100" => rgb <= "000000";
					when "01000100011011101" => rgb <= "000000";
					when "01000100011011110" => rgb <= "000000";
					when "01000100011011111" => rgb <= "000000";
					when "01000100011100000" => rgb <= "000000";
					when "01000100011100001" => rgb <= "000000";
					when "01000100011100010" => rgb <= "000000";
					when "01000100011100011" => rgb <= "000000";
					when "01000100011100100" => rgb <= "000000";
					when "01000100011100101" => rgb <= "000000";
					when "01000100011100110" => rgb <= "000000";
					when "01000100011100111" => rgb <= "000000";
					when "01000100011101000" => rgb <= "000000";
					when "01000100011101001" => rgb <= "000000";
					when "01000100011101010" => rgb <= "000000";
					when "01000100011101011" => rgb <= "000000";
					when "01000100011101100" => rgb <= "000000";
					when "01000100011101101" => rgb <= "000000";
					when "01000100011101110" => rgb <= "000000";
					when "01000100011101111" => rgb <= "000000";
					when "01000100011110000" => rgb <= "000000";
					when "01000100011110001" => rgb <= "000000";
					when "01000100011110010" => rgb <= "000000";
					when "01000100011110011" => rgb <= "000000";
					when "01000100011110100" => rgb <= "000000";
					when "01000100011110101" => rgb <= "000000";
					when "01000100011110110" => rgb <= "000000";
					when "01000100011110111" => rgb <= "000000";
					when "01000100011111000" => rgb <= "000000";
					when "01000100011111001" => rgb <= "000000";
					when "01000100011111010" => rgb <= "000000";
					when "01000100011111011" => rgb <= "000000";
					when "01000100011111100" => rgb <= "000000";
					when "01000100011111101" => rgb <= "000000";
					when "01000100011111110" => rgb <= "000000";
					when "01000100011111111" => rgb <= "000000";
					when "01000100100000000" => rgb <= "000000";
					when "01000100100000001" => rgb <= "000000";
					when "01000100100000010" => rgb <= "000000";
					when "01000100100000011" => rgb <= "000000";
					when "01000100100000100" => rgb <= "000000";
					when "01000100100000101" => rgb <= "000000";
					when "01000100100000110" => rgb <= "000000";
					when "01000100100000111" => rgb <= "000000";
					when "01000100100001000" => rgb <= "000000";
					when "01000100100001001" => rgb <= "000000";
					when "01000100100001010" => rgb <= "000000";
					when "01000100100001011" => rgb <= "000000";
					when "01000100100001100" => rgb <= "000000";
					when "01000100100001101" => rgb <= "000000";
					when "01000100100001110" => rgb <= "000000";
					when "01000100100001111" => rgb <= "000000";
					when "01000100100010000" => rgb <= "000000";
					when "01000100100010001" => rgb <= "000000";
					when "01000100100010010" => rgb <= "000000";
					when "01000100100010011" => rgb <= "000000";
					when "01000100100010100" => rgb <= "000000";
					when "01000100100010101" => rgb <= "000000";
					when "01000100100010110" => rgb <= "000000";
					when "01000100100010111" => rgb <= "000000";
					when "01000100100011000" => rgb <= "000000";
					when "01000100100011001" => rgb <= "000000";
					when "01000100100011010" => rgb <= "000000";
					when "01000100100011011" => rgb <= "000000";
					when "01000100100011100" => rgb <= "000000";
					when "01000100100011101" => rgb <= "000000";
					when "01000100100011110" => rgb <= "000000";
					when "01000100100011111" => rgb <= "000000";
					when "01000100100100000" => rgb <= "000000";
					when "01000100100100001" => rgb <= "000000";
					when "01000100100100010" => rgb <= "000000";
					when "01000100100100011" => rgb <= "000000";
					when "01000100100100100" => rgb <= "000000";
					when "01000100100100101" => rgb <= "000000";
					when "01000100100100110" => rgb <= "000000";
					when "01000100100100111" => rgb <= "000000";
					when "01000100100101000" => rgb <= "000000";
					when "01000100100101001" => rgb <= "000000";
					when "01000100100101010" => rgb <= "000000";
					when "01000100100101011" => rgb <= "000000";
					when "01000100100101100" => rgb <= "000000";
					when "01000100100101101" => rgb <= "000000";
					when "01000100100101110" => rgb <= "000000";
					when "01000100100101111" => rgb <= "000000";
					when "01000100100110000" => rgb <= "000000";
					when "01000100100110001" => rgb <= "000000";
					when "01000100100110010" => rgb <= "000000";
					when "01000100100110011" => rgb <= "000000";
					when "01000100100110100" => rgb <= "000000";
					when "01000100100110101" => rgb <= "000000";
					when "01000100100110110" => rgb <= "000000";
					when "01000100100110111" => rgb <= "000000";
					when "01000100100111000" => rgb <= "000000";
					when "01000100100111001" => rgb <= "000000";
					when "01000100100111010" => rgb <= "000000";
					when "01000100100111011" => rgb <= "000000";
					when "01000100100111100" => rgb <= "000000";
					when "01000100100111101" => rgb <= "000000";
					when "01000100100111110" => rgb <= "000000";
					when "01000100100111111" => rgb <= "000000";
					when "01000101000000000" => rgb <= "000000";
					when "01000101000000001" => rgb <= "000000";
					when "01000101000000010" => rgb <= "000000";
					when "01000101000000011" => rgb <= "000000";
					when "01000101000000100" => rgb <= "000000";
					when "01000101000000101" => rgb <= "000000";
					when "01000101000000110" => rgb <= "000000";
					when "01000101000000111" => rgb <= "000000";
					when "01000101000001000" => rgb <= "000000";
					when "01000101000001001" => rgb <= "000000";
					when "01000101000001010" => rgb <= "000000";
					when "01000101000001011" => rgb <= "000000";
					when "01000101000001100" => rgb <= "000000";
					when "01000101000001101" => rgb <= "000000";
					when "01000101000001110" => rgb <= "000000";
					when "01000101000001111" => rgb <= "000000";
					when "01000101000010000" => rgb <= "000000";
					when "01000101000010001" => rgb <= "000000";
					when "01000101000010010" => rgb <= "000000";
					when "01000101000010011" => rgb <= "000000";
					when "01000101000010100" => rgb <= "000000";
					when "01000101000010101" => rgb <= "000000";
					when "01000101000010110" => rgb <= "000000";
					when "01000101000010111" => rgb <= "000000";
					when "01000101000011000" => rgb <= "000000";
					when "01000101000011001" => rgb <= "000000";
					when "01000101000011010" => rgb <= "000000";
					when "01000101000011011" => rgb <= "000000";
					when "01000101000011100" => rgb <= "000000";
					when "01000101000011101" => rgb <= "000000";
					when "01000101000011110" => rgb <= "000000";
					when "01000101000011111" => rgb <= "000000";
					when "01000101000100000" => rgb <= "000000";
					when "01000101000100001" => rgb <= "000000";
					when "01000101000100010" => rgb <= "000000";
					when "01000101000100011" => rgb <= "000000";
					when "01000101000100100" => rgb <= "000000";
					when "01000101000100101" => rgb <= "000000";
					when "01000101000100110" => rgb <= "000000";
					when "01000101000100111" => rgb <= "000000";
					when "01000101000101000" => rgb <= "000000";
					when "01000101000101001" => rgb <= "000000";
					when "01000101000101010" => rgb <= "000000";
					when "01000101000101011" => rgb <= "000000";
					when "01000101000101100" => rgb <= "000000";
					when "01000101000101101" => rgb <= "000000";
					when "01000101000101110" => rgb <= "000000";
					when "01000101000101111" => rgb <= "000000";
					when "01000101000110000" => rgb <= "000000";
					when "01000101000110001" => rgb <= "000000";
					when "01000101000110010" => rgb <= "000000";
					when "01000101000110011" => rgb <= "000000";
					when "01000101000110100" => rgb <= "000000";
					when "01000101000110101" => rgb <= "000000";
					when "01000101000110110" => rgb <= "000000";
					when "01000101000110111" => rgb <= "000000";
					when "01000101000111000" => rgb <= "000000";
					when "01000101000111001" => rgb <= "000000";
					when "01000101000111010" => rgb <= "000000";
					when "01000101000111011" => rgb <= "000000";
					when "01000101000111100" => rgb <= "000000";
					when "01000101000111101" => rgb <= "000000";
					when "01000101000111110" => rgb <= "000000";
					when "01000101000111111" => rgb <= "000000";
					when "01000101001000000" => rgb <= "000000";
					when "01000101001000001" => rgb <= "000000";
					when "01000101001000010" => rgb <= "000000";
					when "01000101001000011" => rgb <= "000000";
					when "01000101001000100" => rgb <= "000000";
					when "01000101001000101" => rgb <= "000000";
					when "01000101001000110" => rgb <= "000000";
					when "01000101001000111" => rgb <= "000000";
					when "01000101001001000" => rgb <= "000000";
					when "01000101001001001" => rgb <= "000000";
					when "01000101001001010" => rgb <= "000000";
					when "01000101001001011" => rgb <= "000000";
					when "01000101001001100" => rgb <= "000000";
					when "01000101001001101" => rgb <= "000000";
					when "01000101001001110" => rgb <= "000000";
					when "01000101001001111" => rgb <= "000000";
					when "01000101001010000" => rgb <= "000000";
					when "01000101001010001" => rgb <= "000000";
					when "01000101001010010" => rgb <= "000000";
					when "01000101001010011" => rgb <= "000000";
					when "01000101001010100" => rgb <= "000000";
					when "01000101001010101" => rgb <= "000000";
					when "01000101001010110" => rgb <= "000000";
					when "01000101001010111" => rgb <= "000000";
					when "01000101001011000" => rgb <= "000000";
					when "01000101001011001" => rgb <= "000000";
					when "01000101001011010" => rgb <= "000000";
					when "01000101001011011" => rgb <= "000000";
					when "01000101001011100" => rgb <= "000000";
					when "01000101001011101" => rgb <= "000000";
					when "01000101001011110" => rgb <= "000000";
					when "01000101001011111" => rgb <= "000000";
					when "01000101001100000" => rgb <= "000000";
					when "01000101001100001" => rgb <= "000000";
					when "01000101001100010" => rgb <= "000000";
					when "01000101001100011" => rgb <= "000000";
					when "01000101001100100" => rgb <= "000000";
					when "01000101001100101" => rgb <= "000000";
					when "01000101001100110" => rgb <= "000000";
					when "01000101001100111" => rgb <= "000000";
					when "01000101001101000" => rgb <= "000000";
					when "01000101001101001" => rgb <= "000000";
					when "01000101001101010" => rgb <= "000000";
					when "01000101001101011" => rgb <= "000000";
					when "01000101001101100" => rgb <= "000000";
					when "01000101001101101" => rgb <= "000000";
					when "01000101001101110" => rgb <= "000000";
					when "01000101001101111" => rgb <= "000000";
					when "01000101001110000" => rgb <= "000000";
					when "01000101001110001" => rgb <= "010000";
					when "01000101001110010" => rgb <= "101000";
					when "01000101001110011" => rgb <= "101000";
					when "01000101001110100" => rgb <= "101000";
					when "01000101001110101" => rgb <= "101000";
					when "01000101001110110" => rgb <= "101000";
					when "01000101001110111" => rgb <= "101000";
					when "01000101001111000" => rgb <= "101000";
					when "01000101001111001" => rgb <= "101000";
					when "01000101001111010" => rgb <= "101000";
					when "01000101001111011" => rgb <= "101000";
					when "01000101001111100" => rgb <= "101000";
					when "01000101001111101" => rgb <= "101000";
					when "01000101001111110" => rgb <= "101000";
					when "01000101001111111" => rgb <= "101000";
					when "01000101010000000" => rgb <= "101000";
					when "01000101010000001" => rgb <= "101000";
					when "01000101010000010" => rgb <= "101000";
					when "01000101010000011" => rgb <= "101000";
					when "01000101010000100" => rgb <= "101000";
					when "01000101010000101" => rgb <= "101000";
					when "01000101010000110" => rgb <= "101000";
					when "01000101010000111" => rgb <= "101000";
					when "01000101010001000" => rgb <= "101000";
					when "01000101010001001" => rgb <= "101000";
					when "01000101010001010" => rgb <= "101000";
					when "01000101010001011" => rgb <= "101000";
					when "01000101010001100" => rgb <= "101000";
					when "01000101010001101" => rgb <= "101000";
					when "01000101010001110" => rgb <= "101000";
					when "01000101010001111" => rgb <= "101000";
					when "01000101010010000" => rgb <= "101000";
					when "01000101010010001" => rgb <= "101000";
					when "01000101010010010" => rgb <= "101000";
					when "01000101010010011" => rgb <= "101000";
					when "01000101010010100" => rgb <= "101000";
					when "01000101010010101" => rgb <= "101000";
					when "01000101010010110" => rgb <= "101000";
					when "01000101010010111" => rgb <= "101000";
					when "01000101010011000" => rgb <= "101000";
					when "01000101010011001" => rgb <= "101000";
					when "01000101010011010" => rgb <= "101000";
					when "01000101010011011" => rgb <= "101000";
					when "01000101010011100" => rgb <= "101000";
					when "01000101010011101" => rgb <= "101000";
					when "01000101010011110" => rgb <= "101000";
					when "01000101010011111" => rgb <= "101000";
					when "01000101010100000" => rgb <= "101000";
					when "01000101010100001" => rgb <= "101000";
					when "01000101010100010" => rgb <= "101000";
					when "01000101010100011" => rgb <= "101000";
					when "01000101010100100" => rgb <= "101000";
					when "01000101010100101" => rgb <= "101000";
					when "01000101010100110" => rgb <= "101000";
					when "01000101010100111" => rgb <= "101000";
					when "01000101010101000" => rgb <= "101000";
					when "01000101010101001" => rgb <= "101000";
					when "01000101010101010" => rgb <= "101000";
					when "01000101010101011" => rgb <= "101000";
					when "01000101010101100" => rgb <= "101000";
					when "01000101010101101" => rgb <= "101000";
					when "01000101010101110" => rgb <= "101000";
					when "01000101010101111" => rgb <= "101000";
					when "01000101010110000" => rgb <= "101000";
					when "01000101010110001" => rgb <= "101000";
					when "01000101010110010" => rgb <= "101000";
					when "01000101010110011" => rgb <= "101000";
					when "01000101010110100" => rgb <= "101000";
					when "01000101010110101" => rgb <= "101000";
					when "01000101010110110" => rgb <= "101000";
					when "01000101010110111" => rgb <= "101000";
					when "01000101010111000" => rgb <= "101000";
					when "01000101010111001" => rgb <= "101000";
					when "01000101010111010" => rgb <= "101000";
					when "01000101010111011" => rgb <= "101000";
					when "01000101010111100" => rgb <= "101000";
					when "01000101010111101" => rgb <= "101000";
					when "01000101010111110" => rgb <= "101000";
					when "01000101010111111" => rgb <= "101000";
					when "01000101011000000" => rgb <= "101000";
					when "01000101011000001" => rgb <= "101000";
					when "01000101011000010" => rgb <= "101000";
					when "01000101011000011" => rgb <= "101000";
					when "01000101011000100" => rgb <= "101000";
					when "01000101011000101" => rgb <= "101000";
					when "01000101011000110" => rgb <= "101000";
					when "01000101011000111" => rgb <= "101000";
					when "01000101011001000" => rgb <= "101000";
					when "01000101011001001" => rgb <= "101000";
					when "01000101011001010" => rgb <= "101000";
					when "01000101011001011" => rgb <= "101000";
					when "01000101011001100" => rgb <= "000000";
					when "01000101011001101" => rgb <= "000000";
					when "01000101011001110" => rgb <= "000000";
					when "01000101011001111" => rgb <= "000000";
					when "01000101011010000" => rgb <= "000000";
					when "01000101011010001" => rgb <= "000000";
					when "01000101011010010" => rgb <= "000000";
					when "01000101011010011" => rgb <= "000000";
					when "01000101011010100" => rgb <= "000000";
					when "01000101011010101" => rgb <= "000000";
					when "01000101011010110" => rgb <= "000000";
					when "01000101011010111" => rgb <= "000000";
					when "01000101011011000" => rgb <= "000000";
					when "01000101011011001" => rgb <= "000000";
					when "01000101011011010" => rgb <= "000000";
					when "01000101011011011" => rgb <= "000000";
					when "01000101011011100" => rgb <= "000000";
					when "01000101011011101" => rgb <= "000000";
					when "01000101011011110" => rgb <= "000000";
					when "01000101011011111" => rgb <= "000000";
					when "01000101011100000" => rgb <= "000000";
					when "01000101011100001" => rgb <= "000000";
					when "01000101011100010" => rgb <= "000000";
					when "01000101011100011" => rgb <= "000000";
					when "01000101011100100" => rgb <= "000000";
					when "01000101011100101" => rgb <= "000000";
					when "01000101011100110" => rgb <= "000000";
					when "01000101011100111" => rgb <= "000000";
					when "01000101011101000" => rgb <= "000000";
					when "01000101011101001" => rgb <= "000000";
					when "01000101011101010" => rgb <= "000000";
					when "01000101011101011" => rgb <= "000000";
					when "01000101011101100" => rgb <= "000000";
					when "01000101011101101" => rgb <= "000000";
					when "01000101011101110" => rgb <= "000000";
					when "01000101011101111" => rgb <= "000000";
					when "01000101011110000" => rgb <= "000000";
					when "01000101011110001" => rgb <= "000000";
					when "01000101011110010" => rgb <= "000000";
					when "01000101011110011" => rgb <= "000000";
					when "01000101011110100" => rgb <= "000000";
					when "01000101011110101" => rgb <= "000000";
					when "01000101011110110" => rgb <= "000000";
					when "01000101011110111" => rgb <= "000000";
					when "01000101011111000" => rgb <= "000000";
					when "01000101011111001" => rgb <= "000000";
					when "01000101011111010" => rgb <= "000000";
					when "01000101011111011" => rgb <= "000000";
					when "01000101011111100" => rgb <= "000000";
					when "01000101011111101" => rgb <= "000000";
					when "01000101011111110" => rgb <= "000000";
					when "01000101011111111" => rgb <= "000000";
					when "01000101100000000" => rgb <= "000000";
					when "01000101100000001" => rgb <= "000000";
					when "01000101100000010" => rgb <= "000000";
					when "01000101100000011" => rgb <= "000000";
					when "01000101100000100" => rgb <= "000000";
					when "01000101100000101" => rgb <= "000000";
					when "01000101100000110" => rgb <= "000000";
					when "01000101100000111" => rgb <= "000000";
					when "01000101100001000" => rgb <= "000000";
					when "01000101100001001" => rgb <= "000000";
					when "01000101100001010" => rgb <= "000000";
					when "01000101100001011" => rgb <= "000000";
					when "01000101100001100" => rgb <= "000000";
					when "01000101100001101" => rgb <= "000000";
					when "01000101100001110" => rgb <= "000000";
					when "01000101100001111" => rgb <= "000000";
					when "01000101100010000" => rgb <= "000000";
					when "01000101100010001" => rgb <= "000000";
					when "01000101100010010" => rgb <= "000000";
					when "01000101100010011" => rgb <= "000000";
					when "01000101100010100" => rgb <= "000000";
					when "01000101100010101" => rgb <= "000000";
					when "01000101100010110" => rgb <= "000000";
					when "01000101100010111" => rgb <= "000000";
					when "01000101100011000" => rgb <= "000000";
					when "01000101100011001" => rgb <= "000000";
					when "01000101100011010" => rgb <= "000000";
					when "01000101100011011" => rgb <= "000000";
					when "01000101100011100" => rgb <= "000000";
					when "01000101100011101" => rgb <= "000000";
					when "01000101100011110" => rgb <= "000000";
					when "01000101100011111" => rgb <= "000000";
					when "01000101100100000" => rgb <= "000000";
					when "01000101100100001" => rgb <= "000000";
					when "01000101100100010" => rgb <= "000000";
					when "01000101100100011" => rgb <= "000000";
					when "01000101100100100" => rgb <= "000000";
					when "01000101100100101" => rgb <= "000000";
					when "01000101100100110" => rgb <= "000000";
					when "01000101100100111" => rgb <= "000000";
					when "01000101100101000" => rgb <= "000000";
					when "01000101100101001" => rgb <= "000000";
					when "01000101100101010" => rgb <= "000000";
					when "01000101100101011" => rgb <= "000000";
					when "01000101100101100" => rgb <= "000000";
					when "01000101100101101" => rgb <= "000000";
					when "01000101100101110" => rgb <= "000000";
					when "01000101100101111" => rgb <= "000000";
					when "01000101100110000" => rgb <= "000000";
					when "01000101100110001" => rgb <= "000000";
					when "01000101100110010" => rgb <= "000000";
					when "01000101100110011" => rgb <= "000000";
					when "01000101100110100" => rgb <= "000000";
					when "01000101100110101" => rgb <= "000000";
					when "01000101100110110" => rgb <= "000000";
					when "01000101100110111" => rgb <= "000000";
					when "01000101100111000" => rgb <= "000000";
					when "01000101100111001" => rgb <= "000000";
					when "01000101100111010" => rgb <= "000000";
					when "01000101100111011" => rgb <= "000000";
					when "01000101100111100" => rgb <= "000000";
					when "01000101100111101" => rgb <= "000000";
					when "01000101100111110" => rgb <= "000000";
					when "01000101100111111" => rgb <= "000000";
					when "01000110000000000" => rgb <= "000000";
					when "01000110000000001" => rgb <= "000000";
					when "01000110000000010" => rgb <= "000000";
					when "01000110000000011" => rgb <= "000000";
					when "01000110000000100" => rgb <= "000000";
					when "01000110000000101" => rgb <= "000000";
					when "01000110000000110" => rgb <= "000000";
					when "01000110000000111" => rgb <= "000000";
					when "01000110000001000" => rgb <= "000000";
					when "01000110000001001" => rgb <= "000000";
					when "01000110000001010" => rgb <= "000000";
					when "01000110000001011" => rgb <= "000000";
					when "01000110000001100" => rgb <= "000000";
					when "01000110000001101" => rgb <= "000000";
					when "01000110000001110" => rgb <= "000000";
					when "01000110000001111" => rgb <= "000000";
					when "01000110000010000" => rgb <= "000000";
					when "01000110000010001" => rgb <= "000000";
					when "01000110000010010" => rgb <= "000000";
					when "01000110000010011" => rgb <= "000000";
					when "01000110000010100" => rgb <= "000000";
					when "01000110000010101" => rgb <= "000000";
					when "01000110000010110" => rgb <= "000000";
					when "01000110000010111" => rgb <= "000000";
					when "01000110000011000" => rgb <= "000000";
					when "01000110000011001" => rgb <= "000000";
					when "01000110000011010" => rgb <= "000000";
					when "01000110000011011" => rgb <= "000000";
					when "01000110000011100" => rgb <= "000000";
					when "01000110000011101" => rgb <= "000000";
					when "01000110000011110" => rgb <= "000000";
					when "01000110000011111" => rgb <= "000000";
					when "01000110000100000" => rgb <= "000000";
					when "01000110000100001" => rgb <= "000000";
					when "01000110000100010" => rgb <= "000000";
					when "01000110000100011" => rgb <= "000000";
					when "01000110000100100" => rgb <= "000000";
					when "01000110000100101" => rgb <= "000000";
					when "01000110000100110" => rgb <= "000000";
					when "01000110000100111" => rgb <= "000000";
					when "01000110000101000" => rgb <= "000000";
					when "01000110000101001" => rgb <= "000000";
					when "01000110000101010" => rgb <= "000000";
					when "01000110000101011" => rgb <= "000000";
					when "01000110000101100" => rgb <= "000000";
					when "01000110000101101" => rgb <= "000000";
					when "01000110000101110" => rgb <= "000000";
					when "01000110000101111" => rgb <= "000000";
					when "01000110000110000" => rgb <= "000000";
					when "01000110000110001" => rgb <= "000000";
					when "01000110000110010" => rgb <= "000000";
					when "01000110000110011" => rgb <= "000000";
					when "01000110000110100" => rgb <= "000000";
					when "01000110000110101" => rgb <= "000000";
					when "01000110000110110" => rgb <= "000000";
					when "01000110000110111" => rgb <= "000000";
					when "01000110000111000" => rgb <= "000000";
					when "01000110000111001" => rgb <= "000000";
					when "01000110000111010" => rgb <= "000000";
					when "01000110000111011" => rgb <= "000000";
					when "01000110000111100" => rgb <= "000000";
					when "01000110000111101" => rgb <= "000000";
					when "01000110000111110" => rgb <= "000000";
					when "01000110000111111" => rgb <= "000000";
					when "01000110001000000" => rgb <= "000000";
					when "01000110001000001" => rgb <= "000000";
					when "01000110001000010" => rgb <= "000000";
					when "01000110001000011" => rgb <= "000000";
					when "01000110001000100" => rgb <= "000000";
					when "01000110001000101" => rgb <= "000000";
					when "01000110001000110" => rgb <= "000000";
					when "01000110001000111" => rgb <= "000000";
					when "01000110001001000" => rgb <= "000000";
					when "01000110001001001" => rgb <= "000000";
					when "01000110001001010" => rgb <= "000000";
					when "01000110001001011" => rgb <= "000000";
					when "01000110001001100" => rgb <= "000000";
					when "01000110001001101" => rgb <= "000000";
					when "01000110001001110" => rgb <= "000000";
					when "01000110001001111" => rgb <= "000000";
					when "01000110001010000" => rgb <= "000000";
					when "01000110001010001" => rgb <= "000000";
					when "01000110001010010" => rgb <= "000000";
					when "01000110001010011" => rgb <= "000000";
					when "01000110001010100" => rgb <= "000000";
					when "01000110001010101" => rgb <= "000000";
					when "01000110001010110" => rgb <= "000000";
					when "01000110001010111" => rgb <= "000000";
					when "01000110001011000" => rgb <= "000000";
					when "01000110001011001" => rgb <= "000000";
					when "01000110001011010" => rgb <= "000000";
					when "01000110001011011" => rgb <= "000000";
					when "01000110001011100" => rgb <= "000000";
					when "01000110001011101" => rgb <= "000000";
					when "01000110001011110" => rgb <= "000000";
					when "01000110001011111" => rgb <= "000000";
					when "01000110001100000" => rgb <= "000000";
					when "01000110001100001" => rgb <= "000000";
					when "01000110001100010" => rgb <= "000000";
					when "01000110001100011" => rgb <= "000000";
					when "01000110001100100" => rgb <= "000000";
					when "01000110001100101" => rgb <= "000000";
					when "01000110001100110" => rgb <= "000000";
					when "01000110001100111" => rgb <= "000000";
					when "01000110001101000" => rgb <= "000000";
					when "01000110001101001" => rgb <= "000000";
					when "01000110001101010" => rgb <= "000000";
					when "01000110001101011" => rgb <= "000000";
					when "01000110001101100" => rgb <= "000000";
					when "01000110001101101" => rgb <= "000000";
					when "01000110001101110" => rgb <= "000000";
					when "01000110001101111" => rgb <= "000000";
					when "01000110001110000" => rgb <= "000000";
					when "01000110001110001" => rgb <= "010000";
					when "01000110001110010" => rgb <= "101000";
					when "01000110001110011" => rgb <= "101000";
					when "01000110001110100" => rgb <= "101000";
					when "01000110001110101" => rgb <= "101000";
					when "01000110001110110" => rgb <= "101000";
					when "01000110001110111" => rgb <= "101000";
					when "01000110001111000" => rgb <= "101000";
					when "01000110001111001" => rgb <= "101000";
					when "01000110001111010" => rgb <= "101000";
					when "01000110001111011" => rgb <= "101000";
					when "01000110001111100" => rgb <= "101000";
					when "01000110001111101" => rgb <= "101000";
					when "01000110001111110" => rgb <= "101000";
					when "01000110001111111" => rgb <= "101000";
					when "01000110010000000" => rgb <= "101000";
					when "01000110010000001" => rgb <= "101000";
					when "01000110010000010" => rgb <= "101000";
					when "01000110010000011" => rgb <= "101000";
					when "01000110010000100" => rgb <= "101000";
					when "01000110010000101" => rgb <= "101000";
					when "01000110010000110" => rgb <= "101000";
					when "01000110010000111" => rgb <= "101000";
					when "01000110010001000" => rgb <= "101000";
					when "01000110010001001" => rgb <= "101000";
					when "01000110010001010" => rgb <= "101000";
					when "01000110010001011" => rgb <= "101000";
					when "01000110010001100" => rgb <= "101000";
					when "01000110010001101" => rgb <= "101000";
					when "01000110010001110" => rgb <= "101000";
					when "01000110010001111" => rgb <= "101000";
					when "01000110010010000" => rgb <= "101000";
					when "01000110010010001" => rgb <= "101000";
					when "01000110010010010" => rgb <= "101000";
					when "01000110010010011" => rgb <= "101000";
					when "01000110010010100" => rgb <= "101000";
					when "01000110010010101" => rgb <= "101000";
					when "01000110010010110" => rgb <= "101000";
					when "01000110010010111" => rgb <= "101000";
					when "01000110010011000" => rgb <= "101000";
					when "01000110010011001" => rgb <= "101000";
					when "01000110010011010" => rgb <= "101000";
					when "01000110010011011" => rgb <= "101000";
					when "01000110010011100" => rgb <= "101000";
					when "01000110010011101" => rgb <= "101000";
					when "01000110010011110" => rgb <= "101000";
					when "01000110010011111" => rgb <= "101000";
					when "01000110010100000" => rgb <= "101000";
					when "01000110010100001" => rgb <= "101000";
					when "01000110010100010" => rgb <= "101000";
					when "01000110010100011" => rgb <= "101000";
					when "01000110010100100" => rgb <= "101000";
					when "01000110010100101" => rgb <= "101000";
					when "01000110010100110" => rgb <= "101000";
					when "01000110010100111" => rgb <= "101000";
					when "01000110010101000" => rgb <= "101000";
					when "01000110010101001" => rgb <= "101000";
					when "01000110010101010" => rgb <= "101000";
					when "01000110010101011" => rgb <= "101000";
					when "01000110010101100" => rgb <= "101000";
					when "01000110010101101" => rgb <= "101000";
					when "01000110010101110" => rgb <= "101000";
					when "01000110010101111" => rgb <= "101000";
					when "01000110010110000" => rgb <= "101000";
					when "01000110010110001" => rgb <= "101000";
					when "01000110010110010" => rgb <= "101000";
					when "01000110010110011" => rgb <= "101000";
					when "01000110010110100" => rgb <= "101000";
					when "01000110010110101" => rgb <= "101000";
					when "01000110010110110" => rgb <= "101000";
					when "01000110010110111" => rgb <= "101000";
					when "01000110010111000" => rgb <= "101000";
					when "01000110010111001" => rgb <= "101000";
					when "01000110010111010" => rgb <= "101000";
					when "01000110010111011" => rgb <= "101000";
					when "01000110010111100" => rgb <= "101000";
					when "01000110010111101" => rgb <= "101000";
					when "01000110010111110" => rgb <= "101000";
					when "01000110010111111" => rgb <= "101000";
					when "01000110011000000" => rgb <= "101000";
					when "01000110011000001" => rgb <= "101000";
					when "01000110011000010" => rgb <= "101000";
					when "01000110011000011" => rgb <= "101000";
					when "01000110011000100" => rgb <= "101000";
					when "01000110011000101" => rgb <= "101000";
					when "01000110011000110" => rgb <= "101000";
					when "01000110011000111" => rgb <= "101000";
					when "01000110011001000" => rgb <= "101000";
					when "01000110011001001" => rgb <= "101000";
					when "01000110011001010" => rgb <= "101000";
					when "01000110011001011" => rgb <= "101000";
					when "01000110011001100" => rgb <= "000000";
					when "01000110011001101" => rgb <= "000000";
					when "01000110011001110" => rgb <= "000000";
					when "01000110011001111" => rgb <= "000000";
					when "01000110011010000" => rgb <= "000000";
					when "01000110011010001" => rgb <= "000000";
					when "01000110011010010" => rgb <= "000000";
					when "01000110011010011" => rgb <= "000000";
					when "01000110011010100" => rgb <= "000000";
					when "01000110011010101" => rgb <= "000000";
					when "01000110011010110" => rgb <= "000000";
					when "01000110011010111" => rgb <= "000000";
					when "01000110011011000" => rgb <= "000000";
					when "01000110011011001" => rgb <= "000000";
					when "01000110011011010" => rgb <= "000000";
					when "01000110011011011" => rgb <= "000000";
					when "01000110011011100" => rgb <= "000000";
					when "01000110011011101" => rgb <= "000000";
					when "01000110011011110" => rgb <= "000000";
					when "01000110011011111" => rgb <= "000000";
					when "01000110011100000" => rgb <= "000000";
					when "01000110011100001" => rgb <= "000000";
					when "01000110011100010" => rgb <= "000000";
					when "01000110011100011" => rgb <= "000000";
					when "01000110011100100" => rgb <= "000000";
					when "01000110011100101" => rgb <= "000000";
					when "01000110011100110" => rgb <= "000000";
					when "01000110011100111" => rgb <= "000000";
					when "01000110011101000" => rgb <= "000000";
					when "01000110011101001" => rgb <= "000000";
					when "01000110011101010" => rgb <= "000000";
					when "01000110011101011" => rgb <= "000000";
					when "01000110011101100" => rgb <= "000000";
					when "01000110011101101" => rgb <= "000000";
					when "01000110011101110" => rgb <= "000000";
					when "01000110011101111" => rgb <= "000000";
					when "01000110011110000" => rgb <= "000000";
					when "01000110011110001" => rgb <= "000000";
					when "01000110011110010" => rgb <= "000000";
					when "01000110011110011" => rgb <= "000000";
					when "01000110011110100" => rgb <= "000000";
					when "01000110011110101" => rgb <= "000000";
					when "01000110011110110" => rgb <= "000000";
					when "01000110011110111" => rgb <= "000000";
					when "01000110011111000" => rgb <= "000000";
					when "01000110011111001" => rgb <= "000000";
					when "01000110011111010" => rgb <= "000000";
					when "01000110011111011" => rgb <= "000000";
					when "01000110011111100" => rgb <= "000000";
					when "01000110011111101" => rgb <= "000000";
					when "01000110011111110" => rgb <= "000000";
					when "01000110011111111" => rgb <= "000000";
					when "01000110100000000" => rgb <= "000000";
					when "01000110100000001" => rgb <= "000000";
					when "01000110100000010" => rgb <= "000000";
					when "01000110100000011" => rgb <= "000000";
					when "01000110100000100" => rgb <= "000000";
					when "01000110100000101" => rgb <= "000000";
					when "01000110100000110" => rgb <= "000000";
					when "01000110100000111" => rgb <= "000000";
					when "01000110100001000" => rgb <= "000000";
					when "01000110100001001" => rgb <= "000000";
					when "01000110100001010" => rgb <= "000000";
					when "01000110100001011" => rgb <= "000000";
					when "01000110100001100" => rgb <= "000000";
					when "01000110100001101" => rgb <= "000000";
					when "01000110100001110" => rgb <= "000000";
					when "01000110100001111" => rgb <= "000000";
					when "01000110100010000" => rgb <= "000000";
					when "01000110100010001" => rgb <= "000000";
					when "01000110100010010" => rgb <= "000000";
					when "01000110100010011" => rgb <= "000000";
					when "01000110100010100" => rgb <= "000000";
					when "01000110100010101" => rgb <= "000000";
					when "01000110100010110" => rgb <= "000000";
					when "01000110100010111" => rgb <= "000000";
					when "01000110100011000" => rgb <= "000000";
					when "01000110100011001" => rgb <= "000000";
					when "01000110100011010" => rgb <= "000000";
					when "01000110100011011" => rgb <= "000000";
					when "01000110100011100" => rgb <= "000000";
					when "01000110100011101" => rgb <= "000000";
					when "01000110100011110" => rgb <= "000000";
					when "01000110100011111" => rgb <= "000000";
					when "01000110100100000" => rgb <= "000000";
					when "01000110100100001" => rgb <= "000000";
					when "01000110100100010" => rgb <= "000000";
					when "01000110100100011" => rgb <= "000000";
					when "01000110100100100" => rgb <= "000000";
					when "01000110100100101" => rgb <= "000000";
					when "01000110100100110" => rgb <= "000000";
					when "01000110100100111" => rgb <= "000000";
					when "01000110100101000" => rgb <= "000000";
					when "01000110100101001" => rgb <= "000000";
					when "01000110100101010" => rgb <= "000000";
					when "01000110100101011" => rgb <= "000000";
					when "01000110100101100" => rgb <= "000000";
					when "01000110100101101" => rgb <= "000000";
					when "01000110100101110" => rgb <= "000000";
					when "01000110100101111" => rgb <= "000000";
					when "01000110100110000" => rgb <= "000000";
					when "01000110100110001" => rgb <= "000000";
					when "01000110100110010" => rgb <= "000000";
					when "01000110100110011" => rgb <= "000000";
					when "01000110100110100" => rgb <= "000000";
					when "01000110100110101" => rgb <= "000000";
					when "01000110100110110" => rgb <= "000000";
					when "01000110100110111" => rgb <= "000000";
					when "01000110100111000" => rgb <= "000000";
					when "01000110100111001" => rgb <= "000000";
					when "01000110100111010" => rgb <= "000000";
					when "01000110100111011" => rgb <= "000000";
					when "01000110100111100" => rgb <= "000000";
					when "01000110100111101" => rgb <= "000000";
					when "01000110100111110" => rgb <= "000000";
					when "01000110100111111" => rgb <= "000000";
					when "01000111000000000" => rgb <= "000000";
					when "01000111000000001" => rgb <= "000000";
					when "01000111000000010" => rgb <= "000000";
					when "01000111000000011" => rgb <= "000000";
					when "01000111000000100" => rgb <= "000000";
					when "01000111000000101" => rgb <= "000000";
					when "01000111000000110" => rgb <= "000000";
					when "01000111000000111" => rgb <= "000000";
					when "01000111000001000" => rgb <= "000000";
					when "01000111000001001" => rgb <= "000000";
					when "01000111000001010" => rgb <= "000000";
					when "01000111000001011" => rgb <= "000000";
					when "01000111000001100" => rgb <= "000000";
					when "01000111000001101" => rgb <= "000000";
					when "01000111000001110" => rgb <= "000000";
					when "01000111000001111" => rgb <= "000000";
					when "01000111000010000" => rgb <= "000000";
					when "01000111000010001" => rgb <= "000000";
					when "01000111000010010" => rgb <= "000000";
					when "01000111000010011" => rgb <= "000000";
					when "01000111000010100" => rgb <= "000000";
					when "01000111000010101" => rgb <= "000000";
					when "01000111000010110" => rgb <= "000000";
					when "01000111000010111" => rgb <= "000000";
					when "01000111000011000" => rgb <= "000000";
					when "01000111000011001" => rgb <= "000000";
					when "01000111000011010" => rgb <= "000000";
					when "01000111000011011" => rgb <= "000000";
					when "01000111000011100" => rgb <= "000000";
					when "01000111000011101" => rgb <= "000000";
					when "01000111000011110" => rgb <= "000000";
					when "01000111000011111" => rgb <= "000000";
					when "01000111000100000" => rgb <= "000000";
					when "01000111000100001" => rgb <= "000000";
					when "01000111000100010" => rgb <= "000000";
					when "01000111000100011" => rgb <= "000000";
					when "01000111000100100" => rgb <= "000000";
					when "01000111000100101" => rgb <= "000000";
					when "01000111000100110" => rgb <= "000000";
					when "01000111000100111" => rgb <= "000000";
					when "01000111000101000" => rgb <= "000000";
					when "01000111000101001" => rgb <= "000000";
					when "01000111000101010" => rgb <= "000000";
					when "01000111000101011" => rgb <= "000000";
					when "01000111000101100" => rgb <= "000000";
					when "01000111000101101" => rgb <= "000000";
					when "01000111000101110" => rgb <= "000000";
					when "01000111000101111" => rgb <= "000000";
					when "01000111000110000" => rgb <= "000000";
					when "01000111000110001" => rgb <= "000000";
					when "01000111000110010" => rgb <= "000000";
					when "01000111000110011" => rgb <= "000000";
					when "01000111000110100" => rgb <= "000000";
					when "01000111000110101" => rgb <= "000000";
					when "01000111000110110" => rgb <= "000000";
					when "01000111000110111" => rgb <= "000000";
					when "01000111000111000" => rgb <= "000000";
					when "01000111000111001" => rgb <= "000000";
					when "01000111000111010" => rgb <= "000000";
					when "01000111000111011" => rgb <= "000000";
					when "01000111000111100" => rgb <= "000000";
					when "01000111000111101" => rgb <= "000000";
					when "01000111000111110" => rgb <= "000000";
					when "01000111000111111" => rgb <= "000000";
					when "01000111001000000" => rgb <= "000000";
					when "01000111001000001" => rgb <= "000000";
					when "01000111001000010" => rgb <= "000000";
					when "01000111001000011" => rgb <= "000000";
					when "01000111001000100" => rgb <= "000000";
					when "01000111001000101" => rgb <= "000000";
					when "01000111001000110" => rgb <= "000000";
					when "01000111001000111" => rgb <= "000000";
					when "01000111001001000" => rgb <= "000000";
					when "01000111001001001" => rgb <= "000000";
					when "01000111001001010" => rgb <= "000000";
					when "01000111001001011" => rgb <= "000000";
					when "01000111001001100" => rgb <= "000000";
					when "01000111001001101" => rgb <= "000000";
					when "01000111001001110" => rgb <= "000000";
					when "01000111001001111" => rgb <= "000000";
					when "01000111001010000" => rgb <= "000000";
					when "01000111001010001" => rgb <= "000000";
					when "01000111001010010" => rgb <= "000000";
					when "01000111001010011" => rgb <= "000000";
					when "01000111001010100" => rgb <= "000000";
					when "01000111001010101" => rgb <= "000000";
					when "01000111001010110" => rgb <= "000000";
					when "01000111001010111" => rgb <= "000000";
					when "01000111001011000" => rgb <= "000000";
					when "01000111001011001" => rgb <= "000000";
					when "01000111001011010" => rgb <= "000000";
					when "01000111001011011" => rgb <= "000000";
					when "01000111001011100" => rgb <= "000000";
					when "01000111001011101" => rgb <= "000000";
					when "01000111001011110" => rgb <= "000000";
					when "01000111001011111" => rgb <= "000000";
					when "01000111001100000" => rgb <= "000000";
					when "01000111001100001" => rgb <= "000000";
					when "01000111001100010" => rgb <= "000000";
					when "01000111001100011" => rgb <= "000000";
					when "01000111001100100" => rgb <= "000000";
					when "01000111001100101" => rgb <= "000000";
					when "01000111001100110" => rgb <= "000000";
					when "01000111001100111" => rgb <= "000000";
					when "01000111001101000" => rgb <= "000000";
					when "01000111001101001" => rgb <= "000000";
					when "01000111001101010" => rgb <= "000000";
					when "01000111001101011" => rgb <= "000000";
					when "01000111001101100" => rgb <= "000000";
					when "01000111001101101" => rgb <= "000000";
					when "01000111001101110" => rgb <= "000000";
					when "01000111001101111" => rgb <= "000000";
					when "01000111001110000" => rgb <= "000000";
					when "01000111001110001" => rgb <= "010000";
					when "01000111001110010" => rgb <= "101000";
					when "01000111001110011" => rgb <= "101000";
					when "01000111001110100" => rgb <= "101000";
					when "01000111001110101" => rgb <= "101000";
					when "01000111001110110" => rgb <= "101000";
					when "01000111001110111" => rgb <= "101000";
					when "01000111001111000" => rgb <= "101000";
					when "01000111001111001" => rgb <= "101000";
					when "01000111001111010" => rgb <= "101000";
					when "01000111001111011" => rgb <= "101000";
					when "01000111001111100" => rgb <= "101000";
					when "01000111001111101" => rgb <= "101000";
					when "01000111001111110" => rgb <= "101000";
					when "01000111001111111" => rgb <= "101000";
					when "01000111010000000" => rgb <= "101000";
					when "01000111010000001" => rgb <= "101000";
					when "01000111010000010" => rgb <= "101000";
					when "01000111010000011" => rgb <= "101000";
					when "01000111010000100" => rgb <= "101000";
					when "01000111010000101" => rgb <= "101000";
					when "01000111010000110" => rgb <= "101000";
					when "01000111010000111" => rgb <= "101000";
					when "01000111010001000" => rgb <= "101000";
					when "01000111010001001" => rgb <= "101000";
					when "01000111010001010" => rgb <= "101000";
					when "01000111010001011" => rgb <= "101000";
					when "01000111010001100" => rgb <= "101000";
					when "01000111010001101" => rgb <= "101000";
					when "01000111010001110" => rgb <= "101000";
					when "01000111010001111" => rgb <= "101000";
					when "01000111010010000" => rgb <= "101000";
					when "01000111010010001" => rgb <= "101000";
					when "01000111010010010" => rgb <= "101000";
					when "01000111010010011" => rgb <= "101000";
					when "01000111010010100" => rgb <= "101000";
					when "01000111010010101" => rgb <= "101000";
					when "01000111010010110" => rgb <= "101000";
					when "01000111010010111" => rgb <= "101000";
					when "01000111010011000" => rgb <= "101000";
					when "01000111010011001" => rgb <= "101000";
					when "01000111010011010" => rgb <= "101000";
					when "01000111010011011" => rgb <= "101000";
					when "01000111010011100" => rgb <= "101000";
					when "01000111010011101" => rgb <= "101000";
					when "01000111010011110" => rgb <= "101000";
					when "01000111010011111" => rgb <= "101000";
					when "01000111010100000" => rgb <= "101000";
					when "01000111010100001" => rgb <= "101000";
					when "01000111010100010" => rgb <= "101000";
					when "01000111010100011" => rgb <= "101000";
					when "01000111010100100" => rgb <= "101000";
					when "01000111010100101" => rgb <= "101000";
					when "01000111010100110" => rgb <= "101000";
					when "01000111010100111" => rgb <= "101000";
					when "01000111010101000" => rgb <= "101000";
					when "01000111010101001" => rgb <= "101000";
					when "01000111010101010" => rgb <= "101000";
					when "01000111010101011" => rgb <= "101000";
					when "01000111010101100" => rgb <= "101000";
					when "01000111010101101" => rgb <= "101000";
					when "01000111010101110" => rgb <= "101000";
					when "01000111010101111" => rgb <= "101000";
					when "01000111010110000" => rgb <= "101000";
					when "01000111010110001" => rgb <= "101000";
					when "01000111010110010" => rgb <= "101000";
					when "01000111010110011" => rgb <= "101000";
					when "01000111010110100" => rgb <= "101000";
					when "01000111010110101" => rgb <= "101000";
					when "01000111010110110" => rgb <= "101000";
					when "01000111010110111" => rgb <= "101000";
					when "01000111010111000" => rgb <= "101000";
					when "01000111010111001" => rgb <= "101000";
					when "01000111010111010" => rgb <= "101000";
					when "01000111010111011" => rgb <= "101000";
					when "01000111010111100" => rgb <= "101000";
					when "01000111010111101" => rgb <= "101000";
					when "01000111010111110" => rgb <= "101000";
					when "01000111010111111" => rgb <= "101000";
					when "01000111011000000" => rgb <= "101000";
					when "01000111011000001" => rgb <= "101000";
					when "01000111011000010" => rgb <= "101000";
					when "01000111011000011" => rgb <= "101000";
					when "01000111011000100" => rgb <= "101000";
					when "01000111011000101" => rgb <= "101000";
					when "01000111011000110" => rgb <= "101000";
					when "01000111011000111" => rgb <= "101000";
					when "01000111011001000" => rgb <= "101000";
					when "01000111011001001" => rgb <= "101000";
					when "01000111011001010" => rgb <= "101000";
					when "01000111011001011" => rgb <= "101000";
					when "01000111011001100" => rgb <= "000000";
					when "01000111011001101" => rgb <= "000000";
					when "01000111011001110" => rgb <= "000000";
					when "01000111011001111" => rgb <= "000000";
					when "01000111011010000" => rgb <= "000000";
					when "01000111011010001" => rgb <= "000000";
					when "01000111011010010" => rgb <= "000000";
					when "01000111011010011" => rgb <= "000000";
					when "01000111011010100" => rgb <= "000000";
					when "01000111011010101" => rgb <= "000000";
					when "01000111011010110" => rgb <= "000000";
					when "01000111011010111" => rgb <= "000000";
					when "01000111011011000" => rgb <= "000000";
					when "01000111011011001" => rgb <= "000000";
					when "01000111011011010" => rgb <= "000000";
					when "01000111011011011" => rgb <= "000000";
					when "01000111011011100" => rgb <= "000000";
					when "01000111011011101" => rgb <= "000000";
					when "01000111011011110" => rgb <= "000000";
					when "01000111011011111" => rgb <= "000000";
					when "01000111011100000" => rgb <= "000000";
					when "01000111011100001" => rgb <= "000000";
					when "01000111011100010" => rgb <= "000000";
					when "01000111011100011" => rgb <= "000000";
					when "01000111011100100" => rgb <= "000000";
					when "01000111011100101" => rgb <= "000000";
					when "01000111011100110" => rgb <= "000000";
					when "01000111011100111" => rgb <= "000000";
					when "01000111011101000" => rgb <= "000000";
					when "01000111011101001" => rgb <= "000000";
					when "01000111011101010" => rgb <= "000000";
					when "01000111011101011" => rgb <= "000000";
					when "01000111011101100" => rgb <= "000000";
					when "01000111011101101" => rgb <= "000000";
					when "01000111011101110" => rgb <= "000000";
					when "01000111011101111" => rgb <= "000000";
					when "01000111011110000" => rgb <= "000000";
					when "01000111011110001" => rgb <= "000000";
					when "01000111011110010" => rgb <= "000000";
					when "01000111011110011" => rgb <= "000000";
					when "01000111011110100" => rgb <= "000000";
					when "01000111011110101" => rgb <= "000000";
					when "01000111011110110" => rgb <= "000000";
					when "01000111011110111" => rgb <= "000000";
					when "01000111011111000" => rgb <= "000000";
					when "01000111011111001" => rgb <= "000000";
					when "01000111011111010" => rgb <= "000000";
					when "01000111011111011" => rgb <= "000000";
					when "01000111011111100" => rgb <= "000000";
					when "01000111011111101" => rgb <= "000000";
					when "01000111011111110" => rgb <= "000000";
					when "01000111011111111" => rgb <= "000000";
					when "01000111100000000" => rgb <= "000000";
					when "01000111100000001" => rgb <= "000000";
					when "01000111100000010" => rgb <= "000000";
					when "01000111100000011" => rgb <= "000000";
					when "01000111100000100" => rgb <= "000000";
					when "01000111100000101" => rgb <= "000000";
					when "01000111100000110" => rgb <= "000000";
					when "01000111100000111" => rgb <= "000000";
					when "01000111100001000" => rgb <= "000000";
					when "01000111100001001" => rgb <= "000000";
					when "01000111100001010" => rgb <= "000000";
					when "01000111100001011" => rgb <= "000000";
					when "01000111100001100" => rgb <= "000000";
					when "01000111100001101" => rgb <= "000000";
					when "01000111100001110" => rgb <= "000000";
					when "01000111100001111" => rgb <= "000000";
					when "01000111100010000" => rgb <= "000000";
					when "01000111100010001" => rgb <= "000000";
					when "01000111100010010" => rgb <= "000000";
					when "01000111100010011" => rgb <= "000000";
					when "01000111100010100" => rgb <= "000000";
					when "01000111100010101" => rgb <= "000000";
					when "01000111100010110" => rgb <= "000000";
					when "01000111100010111" => rgb <= "000000";
					when "01000111100011000" => rgb <= "000000";
					when "01000111100011001" => rgb <= "000000";
					when "01000111100011010" => rgb <= "000000";
					when "01000111100011011" => rgb <= "000000";
					when "01000111100011100" => rgb <= "000000";
					when "01000111100011101" => rgb <= "000000";
					when "01000111100011110" => rgb <= "000000";
					when "01000111100011111" => rgb <= "000000";
					when "01000111100100000" => rgb <= "000000";
					when "01000111100100001" => rgb <= "000000";
					when "01000111100100010" => rgb <= "000000";
					when "01000111100100011" => rgb <= "000000";
					when "01000111100100100" => rgb <= "000000";
					when "01000111100100101" => rgb <= "000000";
					when "01000111100100110" => rgb <= "000000";
					when "01000111100100111" => rgb <= "000000";
					when "01000111100101000" => rgb <= "000000";
					when "01000111100101001" => rgb <= "000000";
					when "01000111100101010" => rgb <= "000000";
					when "01000111100101011" => rgb <= "000000";
					when "01000111100101100" => rgb <= "000000";
					when "01000111100101101" => rgb <= "000000";
					when "01000111100101110" => rgb <= "000000";
					when "01000111100101111" => rgb <= "000000";
					when "01000111100110000" => rgb <= "000000";
					when "01000111100110001" => rgb <= "000000";
					when "01000111100110010" => rgb <= "000000";
					when "01000111100110011" => rgb <= "000000";
					when "01000111100110100" => rgb <= "000000";
					when "01000111100110101" => rgb <= "000000";
					when "01000111100110110" => rgb <= "000000";
					when "01000111100110111" => rgb <= "000000";
					when "01000111100111000" => rgb <= "000000";
					when "01000111100111001" => rgb <= "000000";
					when "01000111100111010" => rgb <= "000000";
					when "01000111100111011" => rgb <= "000000";
					when "01000111100111100" => rgb <= "000000";
					when "01000111100111101" => rgb <= "000000";
					when "01000111100111110" => rgb <= "000000";
					when "01000111100111111" => rgb <= "000000";
					when "01001000000000000" => rgb <= "000000";
					when "01001000000000001" => rgb <= "000000";
					when "01001000000000010" => rgb <= "000000";
					when "01001000000000011" => rgb <= "000000";
					when "01001000000000100" => rgb <= "000000";
					when "01001000000000101" => rgb <= "000000";
					when "01001000000000110" => rgb <= "000000";
					when "01001000000000111" => rgb <= "000000";
					when "01001000000001000" => rgb <= "000000";
					when "01001000000001001" => rgb <= "000000";
					when "01001000000001010" => rgb <= "000000";
					when "01001000000001011" => rgb <= "000000";
					when "01001000000001100" => rgb <= "000000";
					when "01001000000001101" => rgb <= "000000";
					when "01001000000001110" => rgb <= "000000";
					when "01001000000001111" => rgb <= "000000";
					when "01001000000010000" => rgb <= "000000";
					when "01001000000010001" => rgb <= "000000";
					when "01001000000010010" => rgb <= "000000";
					when "01001000000010011" => rgb <= "000000";
					when "01001000000010100" => rgb <= "000000";
					when "01001000000010101" => rgb <= "000000";
					when "01001000000010110" => rgb <= "000000";
					when "01001000000010111" => rgb <= "000000";
					when "01001000000011000" => rgb <= "000000";
					when "01001000000011001" => rgb <= "000000";
					when "01001000000011010" => rgb <= "000000";
					when "01001000000011011" => rgb <= "000000";
					when "01001000000011100" => rgb <= "000000";
					when "01001000000011101" => rgb <= "000000";
					when "01001000000011110" => rgb <= "000000";
					when "01001000000011111" => rgb <= "000000";
					when "01001000000100000" => rgb <= "000000";
					when "01001000000100001" => rgb <= "000000";
					when "01001000000100010" => rgb <= "000000";
					when "01001000000100011" => rgb <= "000000";
					when "01001000000100100" => rgb <= "000000";
					when "01001000000100101" => rgb <= "000000";
					when "01001000000100110" => rgb <= "000000";
					when "01001000000100111" => rgb <= "000000";
					when "01001000000101000" => rgb <= "000000";
					when "01001000000101001" => rgb <= "000000";
					when "01001000000101010" => rgb <= "000000";
					when "01001000000101011" => rgb <= "000000";
					when "01001000000101100" => rgb <= "000000";
					when "01001000000101101" => rgb <= "000000";
					when "01001000000101110" => rgb <= "000000";
					when "01001000000101111" => rgb <= "000000";
					when "01001000000110000" => rgb <= "000000";
					when "01001000000110001" => rgb <= "000000";
					when "01001000000110010" => rgb <= "000000";
					when "01001000000110011" => rgb <= "000000";
					when "01001000000110100" => rgb <= "000000";
					when "01001000000110101" => rgb <= "000000";
					when "01001000000110110" => rgb <= "000000";
					when "01001000000110111" => rgb <= "000000";
					when "01001000000111000" => rgb <= "000000";
					when "01001000000111001" => rgb <= "000000";
					when "01001000000111010" => rgb <= "000000";
					when "01001000000111011" => rgb <= "000000";
					when "01001000000111100" => rgb <= "000000";
					when "01001000000111101" => rgb <= "000000";
					when "01001000000111110" => rgb <= "000000";
					when "01001000000111111" => rgb <= "000000";
					when "01001000001000000" => rgb <= "000000";
					when "01001000001000001" => rgb <= "000000";
					when "01001000001000010" => rgb <= "000000";
					when "01001000001000011" => rgb <= "000000";
					when "01001000001000100" => rgb <= "000000";
					when "01001000001000101" => rgb <= "000000";
					when "01001000001000110" => rgb <= "000000";
					when "01001000001000111" => rgb <= "000000";
					when "01001000001001000" => rgb <= "000000";
					when "01001000001001001" => rgb <= "000000";
					when "01001000001001010" => rgb <= "000000";
					when "01001000001001011" => rgb <= "000000";
					when "01001000001001100" => rgb <= "000000";
					when "01001000001001101" => rgb <= "000000";
					when "01001000001001110" => rgb <= "000000";
					when "01001000001001111" => rgb <= "000000";
					when "01001000001010000" => rgb <= "000000";
					when "01001000001010001" => rgb <= "000000";
					when "01001000001010010" => rgb <= "000000";
					when "01001000001010011" => rgb <= "000000";
					when "01001000001010100" => rgb <= "000000";
					when "01001000001010101" => rgb <= "000000";
					when "01001000001010110" => rgb <= "000000";
					when "01001000001010111" => rgb <= "000000";
					when "01001000001011000" => rgb <= "000000";
					when "01001000001011001" => rgb <= "000000";
					when "01001000001011010" => rgb <= "000000";
					when "01001000001011011" => rgb <= "000000";
					when "01001000001011100" => rgb <= "000000";
					when "01001000001011101" => rgb <= "000000";
					when "01001000001011110" => rgb <= "000000";
					when "01001000001011111" => rgb <= "000000";
					when "01001000001100000" => rgb <= "000000";
					when "01001000001100001" => rgb <= "000000";
					when "01001000001100010" => rgb <= "000000";
					when "01001000001100011" => rgb <= "000000";
					when "01001000001100100" => rgb <= "000000";
					when "01001000001100101" => rgb <= "000000";
					when "01001000001100110" => rgb <= "000000";
					when "01001000001100111" => rgb <= "000000";
					when "01001000001101000" => rgb <= "000000";
					when "01001000001101001" => rgb <= "000000";
					when "01001000001101010" => rgb <= "000000";
					when "01001000001101011" => rgb <= "000000";
					when "01001000001101100" => rgb <= "000000";
					when "01001000001101101" => rgb <= "000000";
					when "01001000001101110" => rgb <= "000000";
					when "01001000001101111" => rgb <= "000000";
					when "01001000001110000" => rgb <= "000000";
					when "01001000001110001" => rgb <= "010000";
					when "01001000001110010" => rgb <= "101001";
					when "01001000001110011" => rgb <= "101000";
					when "01001000001110100" => rgb <= "111000";
					when "01001000001110101" => rgb <= "111000";
					when "01001000001110110" => rgb <= "101000";
					when "01001000001110111" => rgb <= "111000";
					when "01001000001111000" => rgb <= "101000";
					when "01001000001111001" => rgb <= "101000";
					when "01001000001111010" => rgb <= "101000";
					when "01001000001111011" => rgb <= "101000";
					when "01001000001111100" => rgb <= "101000";
					when "01001000001111101" => rgb <= "101000";
					when "01001000001111110" => rgb <= "101000";
					when "01001000001111111" => rgb <= "101000";
					when "01001000010000000" => rgb <= "111000";
					when "01001000010000001" => rgb <= "111000";
					when "01001000010000010" => rgb <= "101000";
					when "01001000010000011" => rgb <= "111000";
					when "01001000010000100" => rgb <= "101000";
					when "01001000010000101" => rgb <= "101000";
					when "01001000010000110" => rgb <= "111000";
					when "01001000010000111" => rgb <= "101000";
					when "01001000010001000" => rgb <= "101001";
					when "01001000010001001" => rgb <= "101000";
					when "01001000010001010" => rgb <= "101000";
					when "01001000010001011" => rgb <= "101000";
					when "01001000010001100" => rgb <= "101000";
					when "01001000010001101" => rgb <= "101000";
					when "01001000010001110" => rgb <= "101000";
					when "01001000010001111" => rgb <= "101000";
					when "01001000010010000" => rgb <= "101000";
					when "01001000010010001" => rgb <= "101000";
					when "01001000010010010" => rgb <= "101000";
					when "01001000010010011" => rgb <= "101000";
					when "01001000010010100" => rgb <= "101000";
					when "01001000010010101" => rgb <= "101000";
					when "01001000010010110" => rgb <= "101000";
					when "01001000010010111" => rgb <= "101000";
					when "01001000010011000" => rgb <= "101000";
					when "01001000010011001" => rgb <= "101000";
					when "01001000010011010" => rgb <= "101000";
					when "01001000010011011" => rgb <= "101000";
					when "01001000010011100" => rgb <= "101000";
					when "01001000010011101" => rgb <= "101000";
					when "01001000010011110" => rgb <= "101000";
					when "01001000010011111" => rgb <= "101000";
					when "01001000010100000" => rgb <= "101000";
					when "01001000010100001" => rgb <= "101000";
					when "01001000010100010" => rgb <= "101000";
					when "01001000010100011" => rgb <= "101000";
					when "01001000010100100" => rgb <= "101000";
					when "01001000010100101" => rgb <= "101000";
					when "01001000010100110" => rgb <= "101000";
					when "01001000010100111" => rgb <= "101000";
					when "01001000010101000" => rgb <= "101000";
					when "01001000010101001" => rgb <= "101000";
					when "01001000010101010" => rgb <= "101000";
					when "01001000010101011" => rgb <= "101000";
					when "01001000010101100" => rgb <= "101000";
					when "01001000010101101" => rgb <= "101000";
					when "01001000010101110" => rgb <= "101000";
					when "01001000010101111" => rgb <= "101000";
					when "01001000010110000" => rgb <= "101000";
					when "01001000010110001" => rgb <= "101000";
					when "01001000010110010" => rgb <= "101000";
					when "01001000010110011" => rgb <= "101000";
					when "01001000010110100" => rgb <= "111000";
					when "01001000010110101" => rgb <= "101000";
					when "01001000010110110" => rgb <= "101000";
					when "01001000010110111" => rgb <= "101000";
					when "01001000010111000" => rgb <= "101000";
					when "01001000010111001" => rgb <= "101000";
					when "01001000010111010" => rgb <= "101000";
					when "01001000010111011" => rgb <= "101000";
					when "01001000010111100" => rgb <= "101000";
					when "01001000010111101" => rgb <= "101000";
					when "01001000010111110" => rgb <= "101000";
					when "01001000010111111" => rgb <= "101000";
					when "01001000011000000" => rgb <= "101000";
					when "01001000011000001" => rgb <= "101000";
					when "01001000011000010" => rgb <= "101000";
					when "01001000011000011" => rgb <= "101000";
					when "01001000011000100" => rgb <= "101000";
					when "01001000011000101" => rgb <= "101000";
					when "01001000011000110" => rgb <= "101000";
					when "01001000011000111" => rgb <= "101000";
					when "01001000011001000" => rgb <= "101000";
					when "01001000011001001" => rgb <= "101000";
					when "01001000011001010" => rgb <= "101000";
					when "01001000011001011" => rgb <= "101000";
					when "01001000011001100" => rgb <= "010000";
					when "01001000011001101" => rgb <= "000000";
					when "01001000011001110" => rgb <= "000000";
					when "01001000011001111" => rgb <= "000000";
					when "01001000011010000" => rgb <= "000000";
					when "01001000011010001" => rgb <= "000000";
					when "01001000011010010" => rgb <= "000000";
					when "01001000011010011" => rgb <= "000000";
					when "01001000011010100" => rgb <= "000000";
					when "01001000011010101" => rgb <= "000000";
					when "01001000011010110" => rgb <= "000000";
					when "01001000011010111" => rgb <= "000000";
					when "01001000011011000" => rgb <= "000000";
					when "01001000011011001" => rgb <= "000000";
					when "01001000011011010" => rgb <= "000000";
					when "01001000011011011" => rgb <= "000000";
					when "01001000011011100" => rgb <= "000000";
					when "01001000011011101" => rgb <= "000000";
					when "01001000011011110" => rgb <= "000000";
					when "01001000011011111" => rgb <= "000000";
					when "01001000011100000" => rgb <= "000000";
					when "01001000011100001" => rgb <= "000000";
					when "01001000011100010" => rgb <= "000000";
					when "01001000011100011" => rgb <= "000000";
					when "01001000011100100" => rgb <= "000000";
					when "01001000011100101" => rgb <= "000000";
					when "01001000011100110" => rgb <= "000000";
					when "01001000011100111" => rgb <= "000000";
					when "01001000011101000" => rgb <= "000000";
					when "01001000011101001" => rgb <= "000000";
					when "01001000011101010" => rgb <= "000000";
					when "01001000011101011" => rgb <= "000000";
					when "01001000011101100" => rgb <= "000000";
					when "01001000011101101" => rgb <= "000000";
					when "01001000011101110" => rgb <= "000000";
					when "01001000011101111" => rgb <= "000000";
					when "01001000011110000" => rgb <= "000000";
					when "01001000011110001" => rgb <= "000000";
					when "01001000011110010" => rgb <= "000000";
					when "01001000011110011" => rgb <= "000000";
					when "01001000011110100" => rgb <= "000000";
					when "01001000011110101" => rgb <= "000000";
					when "01001000011110110" => rgb <= "000000";
					when "01001000011110111" => rgb <= "000000";
					when "01001000011111000" => rgb <= "000000";
					when "01001000011111001" => rgb <= "000000";
					when "01001000011111010" => rgb <= "000000";
					when "01001000011111011" => rgb <= "000000";
					when "01001000011111100" => rgb <= "000000";
					when "01001000011111101" => rgb <= "000000";
					when "01001000011111110" => rgb <= "000000";
					when "01001000011111111" => rgb <= "000000";
					when "01001000100000000" => rgb <= "000000";
					when "01001000100000001" => rgb <= "000000";
					when "01001000100000010" => rgb <= "000000";
					when "01001000100000011" => rgb <= "000000";
					when "01001000100000100" => rgb <= "000000";
					when "01001000100000101" => rgb <= "000000";
					when "01001000100000110" => rgb <= "000000";
					when "01001000100000111" => rgb <= "000000";
					when "01001000100001000" => rgb <= "000000";
					when "01001000100001001" => rgb <= "000000";
					when "01001000100001010" => rgb <= "000000";
					when "01001000100001011" => rgb <= "000000";
					when "01001000100001100" => rgb <= "000000";
					when "01001000100001101" => rgb <= "000000";
					when "01001000100001110" => rgb <= "000000";
					when "01001000100001111" => rgb <= "000000";
					when "01001000100010000" => rgb <= "000000";
					when "01001000100010001" => rgb <= "000000";
					when "01001000100010010" => rgb <= "000000";
					when "01001000100010011" => rgb <= "000000";
					when "01001000100010100" => rgb <= "000000";
					when "01001000100010101" => rgb <= "000000";
					when "01001000100010110" => rgb <= "000000";
					when "01001000100010111" => rgb <= "000000";
					when "01001000100011000" => rgb <= "000000";
					when "01001000100011001" => rgb <= "000000";
					when "01001000100011010" => rgb <= "000000";
					when "01001000100011011" => rgb <= "000000";
					when "01001000100011100" => rgb <= "000000";
					when "01001000100011101" => rgb <= "000000";
					when "01001000100011110" => rgb <= "000000";
					when "01001000100011111" => rgb <= "000000";
					when "01001000100100000" => rgb <= "000000";
					when "01001000100100001" => rgb <= "000000";
					when "01001000100100010" => rgb <= "000000";
					when "01001000100100011" => rgb <= "000000";
					when "01001000100100100" => rgb <= "000000";
					when "01001000100100101" => rgb <= "000000";
					when "01001000100100110" => rgb <= "000000";
					when "01001000100100111" => rgb <= "000000";
					when "01001000100101000" => rgb <= "000000";
					when "01001000100101001" => rgb <= "000000";
					when "01001000100101010" => rgb <= "000000";
					when "01001000100101011" => rgb <= "000000";
					when "01001000100101100" => rgb <= "000000";
					when "01001000100101101" => rgb <= "000000";
					when "01001000100101110" => rgb <= "000000";
					when "01001000100101111" => rgb <= "000000";
					when "01001000100110000" => rgb <= "000000";
					when "01001000100110001" => rgb <= "000000";
					when "01001000100110010" => rgb <= "000000";
					when "01001000100110011" => rgb <= "000000";
					when "01001000100110100" => rgb <= "000000";
					when "01001000100110101" => rgb <= "000000";
					when "01001000100110110" => rgb <= "000000";
					when "01001000100110111" => rgb <= "000000";
					when "01001000100111000" => rgb <= "000000";
					when "01001000100111001" => rgb <= "000000";
					when "01001000100111010" => rgb <= "000000";
					when "01001000100111011" => rgb <= "000000";
					when "01001000100111100" => rgb <= "000000";
					when "01001000100111101" => rgb <= "000000";
					when "01001000100111110" => rgb <= "000000";
					when "01001000100111111" => rgb <= "000000";
					when "01001001000000000" => rgb <= "000000";
					when "01001001000000001" => rgb <= "000000";
					when "01001001000000010" => rgb <= "000000";
					when "01001001000000011" => rgb <= "000000";
					when "01001001000000100" => rgb <= "000000";
					when "01001001000000101" => rgb <= "000000";
					when "01001001000000110" => rgb <= "000000";
					when "01001001000000111" => rgb <= "000000";
					when "01001001000001000" => rgb <= "000000";
					when "01001001000001001" => rgb <= "000000";
					when "01001001000001010" => rgb <= "000000";
					when "01001001000001011" => rgb <= "000000";
					when "01001001000001100" => rgb <= "000000";
					when "01001001000001101" => rgb <= "000000";
					when "01001001000001110" => rgb <= "000000";
					when "01001001000001111" => rgb <= "000000";
					when "01001001000010000" => rgb <= "000000";
					when "01001001000010001" => rgb <= "000000";
					when "01001001000010010" => rgb <= "000000";
					when "01001001000010011" => rgb <= "000000";
					when "01001001000010100" => rgb <= "000000";
					when "01001001000010101" => rgb <= "000000";
					when "01001001000010110" => rgb <= "000000";
					when "01001001000010111" => rgb <= "000000";
					when "01001001000011000" => rgb <= "000000";
					when "01001001000011001" => rgb <= "000000";
					when "01001001000011010" => rgb <= "000000";
					when "01001001000011011" => rgb <= "000000";
					when "01001001000011100" => rgb <= "000000";
					when "01001001000011101" => rgb <= "000000";
					when "01001001000011110" => rgb <= "000000";
					when "01001001000011111" => rgb <= "000000";
					when "01001001000100000" => rgb <= "000000";
					when "01001001000100001" => rgb <= "000000";
					when "01001001000100010" => rgb <= "000000";
					when "01001001000100011" => rgb <= "000000";
					when "01001001000100100" => rgb <= "000000";
					when "01001001000100101" => rgb <= "000000";
					when "01001001000100110" => rgb <= "000000";
					when "01001001000100111" => rgb <= "000000";
					when "01001001000101000" => rgb <= "000000";
					when "01001001000101001" => rgb <= "000000";
					when "01001001000101010" => rgb <= "000000";
					when "01001001000101011" => rgb <= "000000";
					when "01001001000101100" => rgb <= "000000";
					when "01001001000101101" => rgb <= "000000";
					when "01001001000101110" => rgb <= "000000";
					when "01001001000101111" => rgb <= "000000";
					when "01001001000110000" => rgb <= "000000";
					when "01001001000110001" => rgb <= "000000";
					when "01001001000110010" => rgb <= "000000";
					when "01001001000110011" => rgb <= "000000";
					when "01001001000110100" => rgb <= "000000";
					when "01001001000110101" => rgb <= "000000";
					when "01001001000110110" => rgb <= "000000";
					when "01001001000110111" => rgb <= "000000";
					when "01001001000111000" => rgb <= "000000";
					when "01001001000111001" => rgb <= "000000";
					when "01001001000111010" => rgb <= "000000";
					when "01001001000111011" => rgb <= "000000";
					when "01001001000111100" => rgb <= "000000";
					when "01001001000111101" => rgb <= "000000";
					when "01001001000111110" => rgb <= "000000";
					when "01001001000111111" => rgb <= "000000";
					when "01001001001000000" => rgb <= "000000";
					when "01001001001000001" => rgb <= "000000";
					when "01001001001000010" => rgb <= "000000";
					when "01001001001000011" => rgb <= "000000";
					when "01001001001000100" => rgb <= "000000";
					when "01001001001000101" => rgb <= "000000";
					when "01001001001000110" => rgb <= "000000";
					when "01001001001000111" => rgb <= "000000";
					when "01001001001001000" => rgb <= "000000";
					when "01001001001001001" => rgb <= "000000";
					when "01001001001001010" => rgb <= "000000";
					when "01001001001001011" => rgb <= "000000";
					when "01001001001001100" => rgb <= "000000";
					when "01001001001001101" => rgb <= "000000";
					when "01001001001001110" => rgb <= "000000";
					when "01001001001001111" => rgb <= "000000";
					when "01001001001010000" => rgb <= "000000";
					when "01001001001010001" => rgb <= "000000";
					when "01001001001010010" => rgb <= "000000";
					when "01001001001010011" => rgb <= "000000";
					when "01001001001010100" => rgb <= "000000";
					when "01001001001010101" => rgb <= "000000";
					when "01001001001010110" => rgb <= "000000";
					when "01001001001010111" => rgb <= "000000";
					when "01001001001011000" => rgb <= "000000";
					when "01001001001011001" => rgb <= "000000";
					when "01001001001011010" => rgb <= "000000";
					when "01001001001011011" => rgb <= "000000";
					when "01001001001011100" => rgb <= "000000";
					when "01001001001011101" => rgb <= "000000";
					when "01001001001011110" => rgb <= "000000";
					when "01001001001011111" => rgb <= "000000";
					when "01001001001100000" => rgb <= "000000";
					when "01001001001100001" => rgb <= "000000";
					when "01001001001100010" => rgb <= "000000";
					when "01001001001100011" => rgb <= "000000";
					when "01001001001100100" => rgb <= "000000";
					when "01001001001100101" => rgb <= "000000";
					when "01001001001100110" => rgb <= "000000";
					when "01001001001100111" => rgb <= "000000";
					when "01001001001101000" => rgb <= "000000";
					when "01001001001101001" => rgb <= "000000";
					when "01001001001101010" => rgb <= "000000";
					when "01001001001101011" => rgb <= "000000";
					when "01001001001101100" => rgb <= "000000";
					when "01001001001101101" => rgb <= "000000";
					when "01001001001101110" => rgb <= "000000";
					when "01001001001101111" => rgb <= "000000";
					when "01001001001110000" => rgb <= "000000";
					when "01001001001110001" => rgb <= "000000";
					when "01001001001110010" => rgb <= "101000";
					when "01001001001110011" => rgb <= "101000";
					when "01001001001110100" => rgb <= "101000";
					when "01001001001110101" => rgb <= "101000";
					when "01001001001110110" => rgb <= "101000";
					when "01001001001110111" => rgb <= "101000";
					when "01001001001111000" => rgb <= "101000";
					when "01001001001111001" => rgb <= "101000";
					when "01001001001111010" => rgb <= "101000";
					when "01001001001111011" => rgb <= "101000";
					when "01001001001111100" => rgb <= "101000";
					when "01001001001111101" => rgb <= "101000";
					when "01001001001111110" => rgb <= "101000";
					when "01001001001111111" => rgb <= "101000";
					when "01001001010000000" => rgb <= "101000";
					when "01001001010000001" => rgb <= "101000";
					when "01001001010000010" => rgb <= "101000";
					when "01001001010000011" => rgb <= "101000";
					when "01001001010000100" => rgb <= "101000";
					when "01001001010000101" => rgb <= "101000";
					when "01001001010000110" => rgb <= "101000";
					when "01001001010000111" => rgb <= "101000";
					when "01001001010001000" => rgb <= "101000";
					when "01001001010001001" => rgb <= "101000";
					when "01001001010001010" => rgb <= "101000";
					when "01001001010001011" => rgb <= "101000";
					when "01001001010001100" => rgb <= "101000";
					when "01001001010001101" => rgb <= "101000";
					when "01001001010001110" => rgb <= "101000";
					when "01001001010001111" => rgb <= "101000";
					when "01001001010010000" => rgb <= "101000";
					when "01001001010010001" => rgb <= "101000";
					when "01001001010010010" => rgb <= "101000";
					when "01001001010010011" => rgb <= "101000";
					when "01001001010010100" => rgb <= "101000";
					when "01001001010010101" => rgb <= "101000";
					when "01001001010010110" => rgb <= "101000";
					when "01001001010010111" => rgb <= "101000";
					when "01001001010011000" => rgb <= "101000";
					when "01001001010011001" => rgb <= "101000";
					when "01001001010011010" => rgb <= "101000";
					when "01001001010011011" => rgb <= "101000";
					when "01001001010011100" => rgb <= "101000";
					when "01001001010011101" => rgb <= "101000";
					when "01001001010011110" => rgb <= "101000";
					when "01001001010011111" => rgb <= "101000";
					when "01001001010100000" => rgb <= "101000";
					when "01001001010100001" => rgb <= "101000";
					when "01001001010100010" => rgb <= "101000";
					when "01001001010100011" => rgb <= "101000";
					when "01001001010100100" => rgb <= "101000";
					when "01001001010100101" => rgb <= "101000";
					when "01001001010100110" => rgb <= "101000";
					when "01001001010100111" => rgb <= "101000";
					when "01001001010101000" => rgb <= "101000";
					when "01001001010101001" => rgb <= "101000";
					when "01001001010101010" => rgb <= "101000";
					when "01001001010101011" => rgb <= "101000";
					when "01001001010101100" => rgb <= "101000";
					when "01001001010101101" => rgb <= "101000";
					when "01001001010101110" => rgb <= "101000";
					when "01001001010101111" => rgb <= "101000";
					when "01001001010110000" => rgb <= "101000";
					when "01001001010110001" => rgb <= "101000";
					when "01001001010110010" => rgb <= "101000";
					when "01001001010110011" => rgb <= "101000";
					when "01001001010110100" => rgb <= "111000";
					when "01001001010110101" => rgb <= "101000";
					when "01001001010110110" => rgb <= "010100";
					when "01001001010110111" => rgb <= "100100";
					when "01001001010111000" => rgb <= "100100";
					when "01001001010111001" => rgb <= "100100";
					when "01001001010111010" => rgb <= "100100";
					when "01001001010111011" => rgb <= "100100";
					when "01001001010111100" => rgb <= "100100";
					when "01001001010111101" => rgb <= "100100";
					when "01001001010111110" => rgb <= "100100";
					when "01001001010111111" => rgb <= "100100";
					when "01001001011000000" => rgb <= "100100";
					when "01001001011000001" => rgb <= "100100";
					when "01001001011000010" => rgb <= "100100";
					when "01001001011000011" => rgb <= "100100";
					when "01001001011000100" => rgb <= "100100";
					when "01001001011000101" => rgb <= "100100";
					when "01001001011000110" => rgb <= "100100";
					when "01001001011000111" => rgb <= "100100";
					when "01001001011001000" => rgb <= "100100";
					when "01001001011001001" => rgb <= "100100";
					when "01001001011001010" => rgb <= "100100";
					when "01001001011001011" => rgb <= "100100";
					when "01001001011001100" => rgb <= "000000";
					when "01001001011001101" => rgb <= "000000";
					when "01001001011001110" => rgb <= "000000";
					when "01001001011001111" => rgb <= "000000";
					when "01001001011010000" => rgb <= "000000";
					when "01001001011010001" => rgb <= "000000";
					when "01001001011010010" => rgb <= "000000";
					when "01001001011010011" => rgb <= "000000";
					when "01001001011010100" => rgb <= "000000";
					when "01001001011010101" => rgb <= "000000";
					when "01001001011010110" => rgb <= "000000";
					when "01001001011010111" => rgb <= "000000";
					when "01001001011011000" => rgb <= "000000";
					when "01001001011011001" => rgb <= "000000";
					when "01001001011011010" => rgb <= "000000";
					when "01001001011011011" => rgb <= "000000";
					when "01001001011011100" => rgb <= "000000";
					when "01001001011011101" => rgb <= "000000";
					when "01001001011011110" => rgb <= "000000";
					when "01001001011011111" => rgb <= "000000";
					when "01001001011100000" => rgb <= "000000";
					when "01001001011100001" => rgb <= "000000";
					when "01001001011100010" => rgb <= "000000";
					when "01001001011100011" => rgb <= "000000";
					when "01001001011100100" => rgb <= "000000";
					when "01001001011100101" => rgb <= "000000";
					when "01001001011100110" => rgb <= "000000";
					when "01001001011100111" => rgb <= "000000";
					when "01001001011101000" => rgb <= "000000";
					when "01001001011101001" => rgb <= "000000";
					when "01001001011101010" => rgb <= "000000";
					when "01001001011101011" => rgb <= "000000";
					when "01001001011101100" => rgb <= "000000";
					when "01001001011101101" => rgb <= "000000";
					when "01001001011101110" => rgb <= "000000";
					when "01001001011101111" => rgb <= "000000";
					when "01001001011110000" => rgb <= "000000";
					when "01001001011110001" => rgb <= "000000";
					when "01001001011110010" => rgb <= "000000";
					when "01001001011110011" => rgb <= "000000";
					when "01001001011110100" => rgb <= "000000";
					when "01001001011110101" => rgb <= "000000";
					when "01001001011110110" => rgb <= "000000";
					when "01001001011110111" => rgb <= "000000";
					when "01001001011111000" => rgb <= "000000";
					when "01001001011111001" => rgb <= "000000";
					when "01001001011111010" => rgb <= "000000";
					when "01001001011111011" => rgb <= "000000";
					when "01001001011111100" => rgb <= "000000";
					when "01001001011111101" => rgb <= "000000";
					when "01001001011111110" => rgb <= "000000";
					when "01001001011111111" => rgb <= "000000";
					when "01001001100000000" => rgb <= "000000";
					when "01001001100000001" => rgb <= "000000";
					when "01001001100000010" => rgb <= "000000";
					when "01001001100000011" => rgb <= "000000";
					when "01001001100000100" => rgb <= "000000";
					when "01001001100000101" => rgb <= "000000";
					when "01001001100000110" => rgb <= "000000";
					when "01001001100000111" => rgb <= "000000";
					when "01001001100001000" => rgb <= "000000";
					when "01001001100001001" => rgb <= "000000";
					when "01001001100001010" => rgb <= "000000";
					when "01001001100001011" => rgb <= "000000";
					when "01001001100001100" => rgb <= "000000";
					when "01001001100001101" => rgb <= "000000";
					when "01001001100001110" => rgb <= "000000";
					when "01001001100001111" => rgb <= "000000";
					when "01001001100010000" => rgb <= "000000";
					when "01001001100010001" => rgb <= "000000";
					when "01001001100010010" => rgb <= "000000";
					when "01001001100010011" => rgb <= "000000";
					when "01001001100010100" => rgb <= "000000";
					when "01001001100010101" => rgb <= "000000";
					when "01001001100010110" => rgb <= "000000";
					when "01001001100010111" => rgb <= "000000";
					when "01001001100011000" => rgb <= "000000";
					when "01001001100011001" => rgb <= "000000";
					when "01001001100011010" => rgb <= "000000";
					when "01001001100011011" => rgb <= "000000";
					when "01001001100011100" => rgb <= "000000";
					when "01001001100011101" => rgb <= "000000";
					when "01001001100011110" => rgb <= "000000";
					when "01001001100011111" => rgb <= "000000";
					when "01001001100100000" => rgb <= "000000";
					when "01001001100100001" => rgb <= "000000";
					when "01001001100100010" => rgb <= "000000";
					when "01001001100100011" => rgb <= "000000";
					when "01001001100100100" => rgb <= "000000";
					when "01001001100100101" => rgb <= "000000";
					when "01001001100100110" => rgb <= "000000";
					when "01001001100100111" => rgb <= "000000";
					when "01001001100101000" => rgb <= "000000";
					when "01001001100101001" => rgb <= "000000";
					when "01001001100101010" => rgb <= "000000";
					when "01001001100101011" => rgb <= "000000";
					when "01001001100101100" => rgb <= "000000";
					when "01001001100101101" => rgb <= "000000";
					when "01001001100101110" => rgb <= "000000";
					when "01001001100101111" => rgb <= "000000";
					when "01001001100110000" => rgb <= "000000";
					when "01001001100110001" => rgb <= "000000";
					when "01001001100110010" => rgb <= "000000";
					when "01001001100110011" => rgb <= "000000";
					when "01001001100110100" => rgb <= "000000";
					when "01001001100110101" => rgb <= "000000";
					when "01001001100110110" => rgb <= "000000";
					when "01001001100110111" => rgb <= "000000";
					when "01001001100111000" => rgb <= "000000";
					when "01001001100111001" => rgb <= "000000";
					when "01001001100111010" => rgb <= "000000";
					when "01001001100111011" => rgb <= "000000";
					when "01001001100111100" => rgb <= "000000";
					when "01001001100111101" => rgb <= "000000";
					when "01001001100111110" => rgb <= "000000";
					when "01001001100111111" => rgb <= "000000";
					when "01001010000000000" => rgb <= "000000";
					when "01001010000000001" => rgb <= "000000";
					when "01001010000000010" => rgb <= "000000";
					when "01001010000000011" => rgb <= "000000";
					when "01001010000000100" => rgb <= "000000";
					when "01001010000000101" => rgb <= "000000";
					when "01001010000000110" => rgb <= "000000";
					when "01001010000000111" => rgb <= "000000";
					when "01001010000001000" => rgb <= "000000";
					when "01001010000001001" => rgb <= "000000";
					when "01001010000001010" => rgb <= "000000";
					when "01001010000001011" => rgb <= "000000";
					when "01001010000001100" => rgb <= "000000";
					when "01001010000001101" => rgb <= "000000";
					when "01001010000001110" => rgb <= "000000";
					when "01001010000001111" => rgb <= "000000";
					when "01001010000010000" => rgb <= "000000";
					when "01001010000010001" => rgb <= "000000";
					when "01001010000010010" => rgb <= "000000";
					when "01001010000010011" => rgb <= "000000";
					when "01001010000010100" => rgb <= "000000";
					when "01001010000010101" => rgb <= "000000";
					when "01001010000010110" => rgb <= "000000";
					when "01001010000010111" => rgb <= "000000";
					when "01001010000011000" => rgb <= "000000";
					when "01001010000011001" => rgb <= "000000";
					when "01001010000011010" => rgb <= "000000";
					when "01001010000011011" => rgb <= "000000";
					when "01001010000011100" => rgb <= "000000";
					when "01001010000011101" => rgb <= "000000";
					when "01001010000011110" => rgb <= "000000";
					when "01001010000011111" => rgb <= "000000";
					when "01001010000100000" => rgb <= "000000";
					when "01001010000100001" => rgb <= "000000";
					when "01001010000100010" => rgb <= "000000";
					when "01001010000100011" => rgb <= "000000";
					when "01001010000100100" => rgb <= "000000";
					when "01001010000100101" => rgb <= "000000";
					when "01001010000100110" => rgb <= "000000";
					when "01001010000100111" => rgb <= "000000";
					when "01001010000101000" => rgb <= "000000";
					when "01001010000101001" => rgb <= "000000";
					when "01001010000101010" => rgb <= "000000";
					when "01001010000101011" => rgb <= "000000";
					when "01001010000101100" => rgb <= "000000";
					when "01001010000101101" => rgb <= "000000";
					when "01001010000101110" => rgb <= "000000";
					when "01001010000101111" => rgb <= "000000";
					when "01001010000110000" => rgb <= "000000";
					when "01001010000110001" => rgb <= "000000";
					when "01001010000110010" => rgb <= "000000";
					when "01001010000110011" => rgb <= "000000";
					when "01001010000110100" => rgb <= "000000";
					when "01001010000110101" => rgb <= "000000";
					when "01001010000110110" => rgb <= "000000";
					when "01001010000110111" => rgb <= "000000";
					when "01001010000111000" => rgb <= "000000";
					when "01001010000111001" => rgb <= "000000";
					when "01001010000111010" => rgb <= "000000";
					when "01001010000111011" => rgb <= "000000";
					when "01001010000111100" => rgb <= "000000";
					when "01001010000111101" => rgb <= "000000";
					when "01001010000111110" => rgb <= "000000";
					when "01001010000111111" => rgb <= "000000";
					when "01001010001000000" => rgb <= "000000";
					when "01001010001000001" => rgb <= "000000";
					when "01001010001000010" => rgb <= "000000";
					when "01001010001000011" => rgb <= "000000";
					when "01001010001000100" => rgb <= "000000";
					when "01001010001000101" => rgb <= "000000";
					when "01001010001000110" => rgb <= "000000";
					when "01001010001000111" => rgb <= "000000";
					when "01001010001001000" => rgb <= "000000";
					when "01001010001001001" => rgb <= "000000";
					when "01001010001001010" => rgb <= "000000";
					when "01001010001001011" => rgb <= "000000";
					when "01001010001001100" => rgb <= "000000";
					when "01001010001001101" => rgb <= "000000";
					when "01001010001001110" => rgb <= "000000";
					when "01001010001001111" => rgb <= "000000";
					when "01001010001010000" => rgb <= "000000";
					when "01001010001010001" => rgb <= "000000";
					when "01001010001010010" => rgb <= "000000";
					when "01001010001010011" => rgb <= "000000";
					when "01001010001010100" => rgb <= "000000";
					when "01001010001010101" => rgb <= "000000";
					when "01001010001010110" => rgb <= "000000";
					when "01001010001010111" => rgb <= "000000";
					when "01001010001011000" => rgb <= "000000";
					when "01001010001011001" => rgb <= "000000";
					when "01001010001011010" => rgb <= "000000";
					when "01001010001011011" => rgb <= "000000";
					when "01001010001011100" => rgb <= "000000";
					when "01001010001011101" => rgb <= "000000";
					when "01001010001011110" => rgb <= "000000";
					when "01001010001011111" => rgb <= "000000";
					when "01001010001100000" => rgb <= "000000";
					when "01001010001100001" => rgb <= "000000";
					when "01001010001100010" => rgb <= "000000";
					when "01001010001100011" => rgb <= "000000";
					when "01001010001100100" => rgb <= "000000";
					when "01001010001100101" => rgb <= "000000";
					when "01001010001100110" => rgb <= "000000";
					when "01001010001100111" => rgb <= "000000";
					when "01001010001101000" => rgb <= "000000";
					when "01001010001101001" => rgb <= "000000";
					when "01001010001101010" => rgb <= "000000";
					when "01001010001101011" => rgb <= "000000";
					when "01001010001101100" => rgb <= "000000";
					when "01001010001101101" => rgb <= "000000";
					when "01001010001101110" => rgb <= "000000";
					when "01001010001101111" => rgb <= "000000";
					when "01001010001110000" => rgb <= "000000";
					when "01001010001110001" => rgb <= "000000";
					when "01001010001110010" => rgb <= "000000";
					when "01001010001110011" => rgb <= "000000";
					when "01001010001110100" => rgb <= "000000";
					when "01001010001110101" => rgb <= "000000";
					when "01001010001110110" => rgb <= "000000";
					when "01001010001110111" => rgb <= "000000";
					when "01001010001111000" => rgb <= "000000";
					when "01001010001111001" => rgb <= "000000";
					when "01001010001111010" => rgb <= "000000";
					when "01001010001111011" => rgb <= "000000";
					when "01001010001111100" => rgb <= "000000";
					when "01001010001111101" => rgb <= "000000";
					when "01001010001111110" => rgb <= "000000";
					when "01001010001111111" => rgb <= "000000";
					when "01001010010000000" => rgb <= "000000";
					when "01001010010000001" => rgb <= "000000";
					when "01001010010000010" => rgb <= "000000";
					when "01001010010000011" => rgb <= "000000";
					when "01001010010000100" => rgb <= "000000";
					when "01001010010000101" => rgb <= "000000";
					when "01001010010000110" => rgb <= "000000";
					when "01001010010000111" => rgb <= "000000";
					when "01001010010001000" => rgb <= "100100";
					when "01001010010001001" => rgb <= "101000";
					when "01001010010001010" => rgb <= "101000";
					when "01001010010001011" => rgb <= "101000";
					when "01001010010001100" => rgb <= "101000";
					when "01001010010001101" => rgb <= "101000";
					when "01001010010001110" => rgb <= "101000";
					when "01001010010001111" => rgb <= "101000";
					when "01001010010010000" => rgb <= "101000";
					when "01001010010010001" => rgb <= "101000";
					when "01001010010010010" => rgb <= "101000";
					when "01001010010010011" => rgb <= "101000";
					when "01001010010010100" => rgb <= "101000";
					when "01001010010010101" => rgb <= "101000";
					when "01001010010010110" => rgb <= "101000";
					when "01001010010010111" => rgb <= "101000";
					when "01001010010011000" => rgb <= "101000";
					when "01001010010011001" => rgb <= "101000";
					when "01001010010011010" => rgb <= "101000";
					when "01001010010011011" => rgb <= "101000";
					when "01001010010011100" => rgb <= "101000";
					when "01001010010011101" => rgb <= "101000";
					when "01001010010011110" => rgb <= "101000";
					when "01001010010011111" => rgb <= "101000";
					when "01001010010100000" => rgb <= "101000";
					when "01001010010100001" => rgb <= "101000";
					when "01001010010100010" => rgb <= "101000";
					when "01001010010100011" => rgb <= "101000";
					when "01001010010100100" => rgb <= "101000";
					when "01001010010100101" => rgb <= "101000";
					when "01001010010100110" => rgb <= "101000";
					when "01001010010100111" => rgb <= "101000";
					when "01001010010101000" => rgb <= "101000";
					when "01001010010101001" => rgb <= "101000";
					when "01001010010101010" => rgb <= "101000";
					when "01001010010101011" => rgb <= "101000";
					when "01001010010101100" => rgb <= "101000";
					when "01001010010101101" => rgb <= "101000";
					when "01001010010101110" => rgb <= "101000";
					when "01001010010101111" => rgb <= "101000";
					when "01001010010110000" => rgb <= "101000";
					when "01001010010110001" => rgb <= "101000";
					when "01001010010110010" => rgb <= "101000";
					when "01001010010110011" => rgb <= "101000";
					when "01001010010110100" => rgb <= "101000";
					when "01001010010110101" => rgb <= "010100";
					when "01001010010110110" => rgb <= "000000";
					when "01001010010110111" => rgb <= "000000";
					when "01001010010111000" => rgb <= "000000";
					when "01001010010111001" => rgb <= "000000";
					when "01001010010111010" => rgb <= "000000";
					when "01001010010111011" => rgb <= "000000";
					when "01001010010111100" => rgb <= "000000";
					when "01001010010111101" => rgb <= "000000";
					when "01001010010111110" => rgb <= "000000";
					when "01001010010111111" => rgb <= "000000";
					when "01001010011000000" => rgb <= "000000";
					when "01001010011000001" => rgb <= "000000";
					when "01001010011000010" => rgb <= "000000";
					when "01001010011000011" => rgb <= "000000";
					when "01001010011000100" => rgb <= "000000";
					when "01001010011000101" => rgb <= "000000";
					when "01001010011000110" => rgb <= "000000";
					when "01001010011000111" => rgb <= "000000";
					when "01001010011001000" => rgb <= "000000";
					when "01001010011001001" => rgb <= "000000";
					when "01001010011001010" => rgb <= "000000";
					when "01001010011001011" => rgb <= "000000";
					when "01001010011001100" => rgb <= "000000";
					when "01001010011001101" => rgb <= "000000";
					when "01001010011001110" => rgb <= "000000";
					when "01001010011001111" => rgb <= "000000";
					when "01001010011010000" => rgb <= "000000";
					when "01001010011010001" => rgb <= "000000";
					when "01001010011010010" => rgb <= "000000";
					when "01001010011010011" => rgb <= "000000";
					when "01001010011010100" => rgb <= "000000";
					when "01001010011010101" => rgb <= "000000";
					when "01001010011010110" => rgb <= "000000";
					when "01001010011010111" => rgb <= "000000";
					when "01001010011011000" => rgb <= "000000";
					when "01001010011011001" => rgb <= "000000";
					when "01001010011011010" => rgb <= "000000";
					when "01001010011011011" => rgb <= "000000";
					when "01001010011011100" => rgb <= "000000";
					when "01001010011011101" => rgb <= "000000";
					when "01001010011011110" => rgb <= "000000";
					when "01001010011011111" => rgb <= "000000";
					when "01001010011100000" => rgb <= "000000";
					when "01001010011100001" => rgb <= "000000";
					when "01001010011100010" => rgb <= "000000";
					when "01001010011100011" => rgb <= "000000";
					when "01001010011100100" => rgb <= "000000";
					when "01001010011100101" => rgb <= "000000";
					when "01001010011100110" => rgb <= "000000";
					when "01001010011100111" => rgb <= "000000";
					when "01001010011101000" => rgb <= "000000";
					when "01001010011101001" => rgb <= "000000";
					when "01001010011101010" => rgb <= "000000";
					when "01001010011101011" => rgb <= "000000";
					when "01001010011101100" => rgb <= "000000";
					when "01001010011101101" => rgb <= "000000";
					when "01001010011101110" => rgb <= "000000";
					when "01001010011101111" => rgb <= "000000";
					when "01001010011110000" => rgb <= "000000";
					when "01001010011110001" => rgb <= "000000";
					when "01001010011110010" => rgb <= "000000";
					when "01001010011110011" => rgb <= "000000";
					when "01001010011110100" => rgb <= "000000";
					when "01001010011110101" => rgb <= "000000";
					when "01001010011110110" => rgb <= "000000";
					when "01001010011110111" => rgb <= "000000";
					when "01001010011111000" => rgb <= "000000";
					when "01001010011111001" => rgb <= "000000";
					when "01001010011111010" => rgb <= "000000";
					when "01001010011111011" => rgb <= "000000";
					when "01001010011111100" => rgb <= "000000";
					when "01001010011111101" => rgb <= "000000";
					when "01001010011111110" => rgb <= "000000";
					when "01001010011111111" => rgb <= "000000";
					when "01001010100000000" => rgb <= "000000";
					when "01001010100000001" => rgb <= "000000";
					when "01001010100000010" => rgb <= "000000";
					when "01001010100000011" => rgb <= "000000";
					when "01001010100000100" => rgb <= "000000";
					when "01001010100000101" => rgb <= "000000";
					when "01001010100000110" => rgb <= "000000";
					when "01001010100000111" => rgb <= "000000";
					when "01001010100001000" => rgb <= "000000";
					when "01001010100001001" => rgb <= "000000";
					when "01001010100001010" => rgb <= "000000";
					when "01001010100001011" => rgb <= "000000";
					when "01001010100001100" => rgb <= "000000";
					when "01001010100001101" => rgb <= "000000";
					when "01001010100001110" => rgb <= "000000";
					when "01001010100001111" => rgb <= "000000";
					when "01001010100010000" => rgb <= "000000";
					when "01001010100010001" => rgb <= "000000";
					when "01001010100010010" => rgb <= "000000";
					when "01001010100010011" => rgb <= "000000";
					when "01001010100010100" => rgb <= "000000";
					when "01001010100010101" => rgb <= "000000";
					when "01001010100010110" => rgb <= "000000";
					when "01001010100010111" => rgb <= "000000";
					when "01001010100011000" => rgb <= "000000";
					when "01001010100011001" => rgb <= "000000";
					when "01001010100011010" => rgb <= "000000";
					when "01001010100011011" => rgb <= "000000";
					when "01001010100011100" => rgb <= "000000";
					when "01001010100011101" => rgb <= "000000";
					when "01001010100011110" => rgb <= "000000";
					when "01001010100011111" => rgb <= "000000";
					when "01001010100100000" => rgb <= "000000";
					when "01001010100100001" => rgb <= "000000";
					when "01001010100100010" => rgb <= "000000";
					when "01001010100100011" => rgb <= "000000";
					when "01001010100100100" => rgb <= "000000";
					when "01001010100100101" => rgb <= "000000";
					when "01001010100100110" => rgb <= "000000";
					when "01001010100100111" => rgb <= "000000";
					when "01001010100101000" => rgb <= "000000";
					when "01001010100101001" => rgb <= "000000";
					when "01001010100101010" => rgb <= "000000";
					when "01001010100101011" => rgb <= "000000";
					when "01001010100101100" => rgb <= "000000";
					when "01001010100101101" => rgb <= "000000";
					when "01001010100101110" => rgb <= "000000";
					when "01001010100101111" => rgb <= "000000";
					when "01001010100110000" => rgb <= "000000";
					when "01001010100110001" => rgb <= "000000";
					when "01001010100110010" => rgb <= "000000";
					when "01001010100110011" => rgb <= "000000";
					when "01001010100110100" => rgb <= "000000";
					when "01001010100110101" => rgb <= "000000";
					when "01001010100110110" => rgb <= "000000";
					when "01001010100110111" => rgb <= "000000";
					when "01001010100111000" => rgb <= "000000";
					when "01001010100111001" => rgb <= "000000";
					when "01001010100111010" => rgb <= "000000";
					when "01001010100111011" => rgb <= "000000";
					when "01001010100111100" => rgb <= "000000";
					when "01001010100111101" => rgb <= "000000";
					when "01001010100111110" => rgb <= "000000";
					when "01001010100111111" => rgb <= "000000";
					when "01001011000000000" => rgb <= "000000";
					when "01001011000000001" => rgb <= "000000";
					when "01001011000000010" => rgb <= "000000";
					when "01001011000000011" => rgb <= "000000";
					when "01001011000000100" => rgb <= "000000";
					when "01001011000000101" => rgb <= "000000";
					when "01001011000000110" => rgb <= "000000";
					when "01001011000000111" => rgb <= "000000";
					when "01001011000001000" => rgb <= "000000";
					when "01001011000001001" => rgb <= "000000";
					when "01001011000001010" => rgb <= "000000";
					when "01001011000001011" => rgb <= "000000";
					when "01001011000001100" => rgb <= "000000";
					when "01001011000001101" => rgb <= "000000";
					when "01001011000001110" => rgb <= "000000";
					when "01001011000001111" => rgb <= "000000";
					when "01001011000010000" => rgb <= "000000";
					when "01001011000010001" => rgb <= "000000";
					when "01001011000010010" => rgb <= "000000";
					when "01001011000010011" => rgb <= "000000";
					when "01001011000010100" => rgb <= "000000";
					when "01001011000010101" => rgb <= "000000";
					when "01001011000010110" => rgb <= "000000";
					when "01001011000010111" => rgb <= "000000";
					when "01001011000011000" => rgb <= "000000";
					when "01001011000011001" => rgb <= "000000";
					when "01001011000011010" => rgb <= "000000";
					when "01001011000011011" => rgb <= "000000";
					when "01001011000011100" => rgb <= "000000";
					when "01001011000011101" => rgb <= "000000";
					when "01001011000011110" => rgb <= "000000";
					when "01001011000011111" => rgb <= "000000";
					when "01001011000100000" => rgb <= "000000";
					when "01001011000100001" => rgb <= "000000";
					when "01001011000100010" => rgb <= "000000";
					when "01001011000100011" => rgb <= "000000";
					when "01001011000100100" => rgb <= "000000";
					when "01001011000100101" => rgb <= "000000";
					when "01001011000100110" => rgb <= "000000";
					when "01001011000100111" => rgb <= "000000";
					when "01001011000101000" => rgb <= "000000";
					when "01001011000101001" => rgb <= "000000";
					when "01001011000101010" => rgb <= "000000";
					when "01001011000101011" => rgb <= "000000";
					when "01001011000101100" => rgb <= "000000";
					when "01001011000101101" => rgb <= "000000";
					when "01001011000101110" => rgb <= "000000";
					when "01001011000101111" => rgb <= "000000";
					when "01001011000110000" => rgb <= "000000";
					when "01001011000110001" => rgb <= "000000";
					when "01001011000110010" => rgb <= "000000";
					when "01001011000110011" => rgb <= "000000";
					when "01001011000110100" => rgb <= "000000";
					when "01001011000110101" => rgb <= "000000";
					when "01001011000110110" => rgb <= "000000";
					when "01001011000110111" => rgb <= "000000";
					when "01001011000111000" => rgb <= "000000";
					when "01001011000111001" => rgb <= "000000";
					when "01001011000111010" => rgb <= "000000";
					when "01001011000111011" => rgb <= "000000";
					when "01001011000111100" => rgb <= "000000";
					when "01001011000111101" => rgb <= "000000";
					when "01001011000111110" => rgb <= "000000";
					when "01001011000111111" => rgb <= "000000";
					when "01001011001000000" => rgb <= "000000";
					when "01001011001000001" => rgb <= "000000";
					when "01001011001000010" => rgb <= "000000";
					when "01001011001000011" => rgb <= "000000";
					when "01001011001000100" => rgb <= "000000";
					when "01001011001000101" => rgb <= "000000";
					when "01001011001000110" => rgb <= "000000";
					when "01001011001000111" => rgb <= "000000";
					when "01001011001001000" => rgb <= "000000";
					when "01001011001001001" => rgb <= "000000";
					when "01001011001001010" => rgb <= "000000";
					when "01001011001001011" => rgb <= "000000";
					when "01001011001001100" => rgb <= "000000";
					when "01001011001001101" => rgb <= "000000";
					when "01001011001001110" => rgb <= "000000";
					when "01001011001001111" => rgb <= "000000";
					when "01001011001010000" => rgb <= "000000";
					when "01001011001010001" => rgb <= "000000";
					when "01001011001010010" => rgb <= "000000";
					when "01001011001010011" => rgb <= "000000";
					when "01001011001010100" => rgb <= "000000";
					when "01001011001010101" => rgb <= "000000";
					when "01001011001010110" => rgb <= "000000";
					when "01001011001010111" => rgb <= "000000";
					when "01001011001011000" => rgb <= "000000";
					when "01001011001011001" => rgb <= "000000";
					when "01001011001011010" => rgb <= "000000";
					when "01001011001011011" => rgb <= "000000";
					when "01001011001011100" => rgb <= "000000";
					when "01001011001011101" => rgb <= "000000";
					when "01001011001011110" => rgb <= "000000";
					when "01001011001011111" => rgb <= "000000";
					when "01001011001100000" => rgb <= "000000";
					when "01001011001100001" => rgb <= "000000";
					when "01001011001100010" => rgb <= "000000";
					when "01001011001100011" => rgb <= "000000";
					when "01001011001100100" => rgb <= "000000";
					when "01001011001100101" => rgb <= "000000";
					when "01001011001100110" => rgb <= "000000";
					when "01001011001100111" => rgb <= "000000";
					when "01001011001101000" => rgb <= "000000";
					when "01001011001101001" => rgb <= "000000";
					when "01001011001101010" => rgb <= "000000";
					when "01001011001101011" => rgb <= "000000";
					when "01001011001101100" => rgb <= "000000";
					when "01001011001101101" => rgb <= "000000";
					when "01001011001101110" => rgb <= "000000";
					when "01001011001101111" => rgb <= "000000";
					when "01001011001110000" => rgb <= "000000";
					when "01001011001110001" => rgb <= "000000";
					when "01001011001110010" => rgb <= "000000";
					when "01001011001110011" => rgb <= "000000";
					when "01001011001110100" => rgb <= "000000";
					when "01001011001110101" => rgb <= "000000";
					when "01001011001110110" => rgb <= "000000";
					when "01001011001110111" => rgb <= "000000";
					when "01001011001111000" => rgb <= "000000";
					when "01001011001111001" => rgb <= "000000";
					when "01001011001111010" => rgb <= "000000";
					when "01001011001111011" => rgb <= "000000";
					when "01001011001111100" => rgb <= "000000";
					when "01001011001111101" => rgb <= "000000";
					when "01001011001111110" => rgb <= "000000";
					when "01001011001111111" => rgb <= "000000";
					when "01001011010000000" => rgb <= "000000";
					when "01001011010000001" => rgb <= "000000";
					when "01001011010000010" => rgb <= "000000";
					when "01001011010000011" => rgb <= "000000";
					when "01001011010000100" => rgb <= "000000";
					when "01001011010000101" => rgb <= "000000";
					when "01001011010000110" => rgb <= "000000";
					when "01001011010000111" => rgb <= "000000";
					when "01001011010001000" => rgb <= "100100";
					when "01001011010001001" => rgb <= "101000";
					when "01001011010001010" => rgb <= "101000";
					when "01001011010001011" => rgb <= "101000";
					when "01001011010001100" => rgb <= "101000";
					when "01001011010001101" => rgb <= "101000";
					when "01001011010001110" => rgb <= "101000";
					when "01001011010001111" => rgb <= "101000";
					when "01001011010010000" => rgb <= "101000";
					when "01001011010010001" => rgb <= "101000";
					when "01001011010010010" => rgb <= "101000";
					when "01001011010010011" => rgb <= "101000";
					when "01001011010010100" => rgb <= "101000";
					when "01001011010010101" => rgb <= "101000";
					when "01001011010010110" => rgb <= "101000";
					when "01001011010010111" => rgb <= "101000";
					when "01001011010011000" => rgb <= "101000";
					when "01001011010011001" => rgb <= "101000";
					when "01001011010011010" => rgb <= "101000";
					when "01001011010011011" => rgb <= "101000";
					when "01001011010011100" => rgb <= "101000";
					when "01001011010011101" => rgb <= "101000";
					when "01001011010011110" => rgb <= "101000";
					when "01001011010011111" => rgb <= "101000";
					when "01001011010100000" => rgb <= "101000";
					when "01001011010100001" => rgb <= "101000";
					when "01001011010100010" => rgb <= "101000";
					when "01001011010100011" => rgb <= "101000";
					when "01001011010100100" => rgb <= "101000";
					when "01001011010100101" => rgb <= "101000";
					when "01001011010100110" => rgb <= "101000";
					when "01001011010100111" => rgb <= "101000";
					when "01001011010101000" => rgb <= "101000";
					when "01001011010101001" => rgb <= "101000";
					when "01001011010101010" => rgb <= "101000";
					when "01001011010101011" => rgb <= "101000";
					when "01001011010101100" => rgb <= "101000";
					when "01001011010101101" => rgb <= "101000";
					when "01001011010101110" => rgb <= "101000";
					when "01001011010101111" => rgb <= "101000";
					when "01001011010110000" => rgb <= "101000";
					when "01001011010110001" => rgb <= "101000";
					when "01001011010110010" => rgb <= "101000";
					when "01001011010110011" => rgb <= "101000";
					when "01001011010110100" => rgb <= "101000";
					when "01001011010110101" => rgb <= "010100";
					when "01001011010110110" => rgb <= "000000";
					when "01001011010110111" => rgb <= "000000";
					when "01001011010111000" => rgb <= "000000";
					when "01001011010111001" => rgb <= "000000";
					when "01001011010111010" => rgb <= "000000";
					when "01001011010111011" => rgb <= "000000";
					when "01001011010111100" => rgb <= "000000";
					when "01001011010111101" => rgb <= "000000";
					when "01001011010111110" => rgb <= "000000";
					when "01001011010111111" => rgb <= "000000";
					when "01001011011000000" => rgb <= "000000";
					when "01001011011000001" => rgb <= "000000";
					when "01001011011000010" => rgb <= "000000";
					when "01001011011000011" => rgb <= "000000";
					when "01001011011000100" => rgb <= "000000";
					when "01001011011000101" => rgb <= "000000";
					when "01001011011000110" => rgb <= "000000";
					when "01001011011000111" => rgb <= "000000";
					when "01001011011001000" => rgb <= "000000";
					when "01001011011001001" => rgb <= "000000";
					when "01001011011001010" => rgb <= "000000";
					when "01001011011001011" => rgb <= "000000";
					when "01001011011001100" => rgb <= "000000";
					when "01001011011001101" => rgb <= "000000";
					when "01001011011001110" => rgb <= "000000";
					when "01001011011001111" => rgb <= "000000";
					when "01001011011010000" => rgb <= "000000";
					when "01001011011010001" => rgb <= "000000";
					when "01001011011010010" => rgb <= "000000";
					when "01001011011010011" => rgb <= "000000";
					when "01001011011010100" => rgb <= "000000";
					when "01001011011010101" => rgb <= "000000";
					when "01001011011010110" => rgb <= "000000";
					when "01001011011010111" => rgb <= "000000";
					when "01001011011011000" => rgb <= "000000";
					when "01001011011011001" => rgb <= "000000";
					when "01001011011011010" => rgb <= "000000";
					when "01001011011011011" => rgb <= "000000";
					when "01001011011011100" => rgb <= "000000";
					when "01001011011011101" => rgb <= "000000";
					when "01001011011011110" => rgb <= "000000";
					when "01001011011011111" => rgb <= "000000";
					when "01001011011100000" => rgb <= "000000";
					when "01001011011100001" => rgb <= "000000";
					when "01001011011100010" => rgb <= "000000";
					when "01001011011100011" => rgb <= "000000";
					when "01001011011100100" => rgb <= "000000";
					when "01001011011100101" => rgb <= "000000";
					when "01001011011100110" => rgb <= "000000";
					when "01001011011100111" => rgb <= "000000";
					when "01001011011101000" => rgb <= "000000";
					when "01001011011101001" => rgb <= "000000";
					when "01001011011101010" => rgb <= "000000";
					when "01001011011101011" => rgb <= "000000";
					when "01001011011101100" => rgb <= "000000";
					when "01001011011101101" => rgb <= "000000";
					when "01001011011101110" => rgb <= "000000";
					when "01001011011101111" => rgb <= "000000";
					when "01001011011110000" => rgb <= "000000";
					when "01001011011110001" => rgb <= "000000";
					when "01001011011110010" => rgb <= "000000";
					when "01001011011110011" => rgb <= "000000";
					when "01001011011110100" => rgb <= "000000";
					when "01001011011110101" => rgb <= "000000";
					when "01001011011110110" => rgb <= "000000";
					when "01001011011110111" => rgb <= "000000";
					when "01001011011111000" => rgb <= "000000";
					when "01001011011111001" => rgb <= "000000";
					when "01001011011111010" => rgb <= "000000";
					when "01001011011111011" => rgb <= "000000";
					when "01001011011111100" => rgb <= "000000";
					when "01001011011111101" => rgb <= "000000";
					when "01001011011111110" => rgb <= "000000";
					when "01001011011111111" => rgb <= "000000";
					when "01001011100000000" => rgb <= "000000";
					when "01001011100000001" => rgb <= "000000";
					when "01001011100000010" => rgb <= "000000";
					when "01001011100000011" => rgb <= "000000";
					when "01001011100000100" => rgb <= "000000";
					when "01001011100000101" => rgb <= "000000";
					when "01001011100000110" => rgb <= "000000";
					when "01001011100000111" => rgb <= "000000";
					when "01001011100001000" => rgb <= "000000";
					when "01001011100001001" => rgb <= "000000";
					when "01001011100001010" => rgb <= "000000";
					when "01001011100001011" => rgb <= "000000";
					when "01001011100001100" => rgb <= "000000";
					when "01001011100001101" => rgb <= "000000";
					when "01001011100001110" => rgb <= "000000";
					when "01001011100001111" => rgb <= "000000";
					when "01001011100010000" => rgb <= "000000";
					when "01001011100010001" => rgb <= "000000";
					when "01001011100010010" => rgb <= "000000";
					when "01001011100010011" => rgb <= "000000";
					when "01001011100010100" => rgb <= "000000";
					when "01001011100010101" => rgb <= "000000";
					when "01001011100010110" => rgb <= "000000";
					when "01001011100010111" => rgb <= "000000";
					when "01001011100011000" => rgb <= "000000";
					when "01001011100011001" => rgb <= "000000";
					when "01001011100011010" => rgb <= "000000";
					when "01001011100011011" => rgb <= "000000";
					when "01001011100011100" => rgb <= "000000";
					when "01001011100011101" => rgb <= "000000";
					when "01001011100011110" => rgb <= "000000";
					when "01001011100011111" => rgb <= "000000";
					when "01001011100100000" => rgb <= "000000";
					when "01001011100100001" => rgb <= "000000";
					when "01001011100100010" => rgb <= "000000";
					when "01001011100100011" => rgb <= "000000";
					when "01001011100100100" => rgb <= "000000";
					when "01001011100100101" => rgb <= "000000";
					when "01001011100100110" => rgb <= "000000";
					when "01001011100100111" => rgb <= "000000";
					when "01001011100101000" => rgb <= "000000";
					when "01001011100101001" => rgb <= "000000";
					when "01001011100101010" => rgb <= "000000";
					when "01001011100101011" => rgb <= "000000";
					when "01001011100101100" => rgb <= "000000";
					when "01001011100101101" => rgb <= "000000";
					when "01001011100101110" => rgb <= "000000";
					when "01001011100101111" => rgb <= "000000";
					when "01001011100110000" => rgb <= "000000";
					when "01001011100110001" => rgb <= "000000";
					when "01001011100110010" => rgb <= "000000";
					when "01001011100110011" => rgb <= "000000";
					when "01001011100110100" => rgb <= "000000";
					when "01001011100110101" => rgb <= "000000";
					when "01001011100110110" => rgb <= "000000";
					when "01001011100110111" => rgb <= "000000";
					when "01001011100111000" => rgb <= "000000";
					when "01001011100111001" => rgb <= "000000";
					when "01001011100111010" => rgb <= "000000";
					when "01001011100111011" => rgb <= "000000";
					when "01001011100111100" => rgb <= "000000";
					when "01001011100111101" => rgb <= "000000";
					when "01001011100111110" => rgb <= "000000";
					when "01001011100111111" => rgb <= "000000";
					when "01001100000000000" => rgb <= "000000";
					when "01001100000000001" => rgb <= "000000";
					when "01001100000000010" => rgb <= "000000";
					when "01001100000000011" => rgb <= "000000";
					when "01001100000000100" => rgb <= "000000";
					when "01001100000000101" => rgb <= "000000";
					when "01001100000000110" => rgb <= "000000";
					when "01001100000000111" => rgb <= "000000";
					when "01001100000001000" => rgb <= "000000";
					when "01001100000001001" => rgb <= "000000";
					when "01001100000001010" => rgb <= "000000";
					when "01001100000001011" => rgb <= "000000";
					when "01001100000001100" => rgb <= "000000";
					when "01001100000001101" => rgb <= "000000";
					when "01001100000001110" => rgb <= "000000";
					when "01001100000001111" => rgb <= "000000";
					when "01001100000010000" => rgb <= "000000";
					when "01001100000010001" => rgb <= "000000";
					when "01001100000010010" => rgb <= "000000";
					when "01001100000010011" => rgb <= "000000";
					when "01001100000010100" => rgb <= "000000";
					when "01001100000010101" => rgb <= "000000";
					when "01001100000010110" => rgb <= "000000";
					when "01001100000010111" => rgb <= "000000";
					when "01001100000011000" => rgb <= "000000";
					when "01001100000011001" => rgb <= "000000";
					when "01001100000011010" => rgb <= "000000";
					when "01001100000011011" => rgb <= "000000";
					when "01001100000011100" => rgb <= "000000";
					when "01001100000011101" => rgb <= "000000";
					when "01001100000011110" => rgb <= "000000";
					when "01001100000011111" => rgb <= "000000";
					when "01001100000100000" => rgb <= "000000";
					when "01001100000100001" => rgb <= "000000";
					when "01001100000100010" => rgb <= "000000";
					when "01001100000100011" => rgb <= "000000";
					when "01001100000100100" => rgb <= "000000";
					when "01001100000100101" => rgb <= "000000";
					when "01001100000100110" => rgb <= "000000";
					when "01001100000100111" => rgb <= "000000";
					when "01001100000101000" => rgb <= "000000";
					when "01001100000101001" => rgb <= "000000";
					when "01001100000101010" => rgb <= "000000";
					when "01001100000101011" => rgb <= "000000";
					when "01001100000101100" => rgb <= "000000";
					when "01001100000101101" => rgb <= "000000";
					when "01001100000101110" => rgb <= "000000";
					when "01001100000101111" => rgb <= "000000";
					when "01001100000110000" => rgb <= "000000";
					when "01001100000110001" => rgb <= "000000";
					when "01001100000110010" => rgb <= "000000";
					when "01001100000110011" => rgb <= "000000";
					when "01001100000110100" => rgb <= "000000";
					when "01001100000110101" => rgb <= "000000";
					when "01001100000110110" => rgb <= "000000";
					when "01001100000110111" => rgb <= "000000";
					when "01001100000111000" => rgb <= "000000";
					when "01001100000111001" => rgb <= "000000";
					when "01001100000111010" => rgb <= "000000";
					when "01001100000111011" => rgb <= "000000";
					when "01001100000111100" => rgb <= "000000";
					when "01001100000111101" => rgb <= "000000";
					when "01001100000111110" => rgb <= "000000";
					when "01001100000111111" => rgb <= "000000";
					when "01001100001000000" => rgb <= "000000";
					when "01001100001000001" => rgb <= "000000";
					when "01001100001000010" => rgb <= "000000";
					when "01001100001000011" => rgb <= "000000";
					when "01001100001000100" => rgb <= "000000";
					when "01001100001000101" => rgb <= "000000";
					when "01001100001000110" => rgb <= "000000";
					when "01001100001000111" => rgb <= "000000";
					when "01001100001001000" => rgb <= "000000";
					when "01001100001001001" => rgb <= "000000";
					when "01001100001001010" => rgb <= "000000";
					when "01001100001001011" => rgb <= "000000";
					when "01001100001001100" => rgb <= "000000";
					when "01001100001001101" => rgb <= "000000";
					when "01001100001001110" => rgb <= "000000";
					when "01001100001001111" => rgb <= "000000";
					when "01001100001010000" => rgb <= "000000";
					when "01001100001010001" => rgb <= "000000";
					when "01001100001010010" => rgb <= "000000";
					when "01001100001010011" => rgb <= "000000";
					when "01001100001010100" => rgb <= "000000";
					when "01001100001010101" => rgb <= "000000";
					when "01001100001010110" => rgb <= "000000";
					when "01001100001010111" => rgb <= "000000";
					when "01001100001011000" => rgb <= "000000";
					when "01001100001011001" => rgb <= "000000";
					when "01001100001011010" => rgb <= "000000";
					when "01001100001011011" => rgb <= "000000";
					when "01001100001011100" => rgb <= "000000";
					when "01001100001011101" => rgb <= "000000";
					when "01001100001011110" => rgb <= "000000";
					when "01001100001011111" => rgb <= "000000";
					when "01001100001100000" => rgb <= "000000";
					when "01001100001100001" => rgb <= "000000";
					when "01001100001100010" => rgb <= "000000";
					when "01001100001100011" => rgb <= "000000";
					when "01001100001100100" => rgb <= "000000";
					when "01001100001100101" => rgb <= "000000";
					when "01001100001100110" => rgb <= "000000";
					when "01001100001100111" => rgb <= "000000";
					when "01001100001101000" => rgb <= "000000";
					when "01001100001101001" => rgb <= "000000";
					when "01001100001101010" => rgb <= "000000";
					when "01001100001101011" => rgb <= "000000";
					when "01001100001101100" => rgb <= "000000";
					when "01001100001101101" => rgb <= "000000";
					when "01001100001101110" => rgb <= "000000";
					when "01001100001101111" => rgb <= "000000";
					when "01001100001110000" => rgb <= "000000";
					when "01001100001110001" => rgb <= "000000";
					when "01001100001110010" => rgb <= "000000";
					when "01001100001110011" => rgb <= "000000";
					when "01001100001110100" => rgb <= "000000";
					when "01001100001110101" => rgb <= "000000";
					when "01001100001110110" => rgb <= "000000";
					when "01001100001110111" => rgb <= "000000";
					when "01001100001111000" => rgb <= "000000";
					when "01001100001111001" => rgb <= "000000";
					when "01001100001111010" => rgb <= "000000";
					when "01001100001111011" => rgb <= "000000";
					when "01001100001111100" => rgb <= "000000";
					when "01001100001111101" => rgb <= "000000";
					when "01001100001111110" => rgb <= "000000";
					when "01001100001111111" => rgb <= "000000";
					when "01001100010000000" => rgb <= "000000";
					when "01001100010000001" => rgb <= "000000";
					when "01001100010000010" => rgb <= "000000";
					when "01001100010000011" => rgb <= "000000";
					when "01001100010000100" => rgb <= "000000";
					when "01001100010000101" => rgb <= "000000";
					when "01001100010000110" => rgb <= "000000";
					when "01001100010000111" => rgb <= "000000";
					when "01001100010001000" => rgb <= "100100";
					when "01001100010001001" => rgb <= "101000";
					when "01001100010001010" => rgb <= "101000";
					when "01001100010001011" => rgb <= "101000";
					when "01001100010001100" => rgb <= "101000";
					when "01001100010001101" => rgb <= "101000";
					when "01001100010001110" => rgb <= "101000";
					when "01001100010001111" => rgb <= "101000";
					when "01001100010010000" => rgb <= "101000";
					when "01001100010010001" => rgb <= "101000";
					when "01001100010010010" => rgb <= "101000";
					when "01001100010010011" => rgb <= "101000";
					when "01001100010010100" => rgb <= "101000";
					when "01001100010010101" => rgb <= "101000";
					when "01001100010010110" => rgb <= "101000";
					when "01001100010010111" => rgb <= "101000";
					when "01001100010011000" => rgb <= "101000";
					when "01001100010011001" => rgb <= "101000";
					when "01001100010011010" => rgb <= "101000";
					when "01001100010011011" => rgb <= "101000";
					when "01001100010011100" => rgb <= "101000";
					when "01001100010011101" => rgb <= "101000";
					when "01001100010011110" => rgb <= "101000";
					when "01001100010011111" => rgb <= "101000";
					when "01001100010100000" => rgb <= "101000";
					when "01001100010100001" => rgb <= "101000";
					when "01001100010100010" => rgb <= "101000";
					when "01001100010100011" => rgb <= "101000";
					when "01001100010100100" => rgb <= "101000";
					when "01001100010100101" => rgb <= "101000";
					when "01001100010100110" => rgb <= "101000";
					when "01001100010100111" => rgb <= "101000";
					when "01001100010101000" => rgb <= "101000";
					when "01001100010101001" => rgb <= "101000";
					when "01001100010101010" => rgb <= "101000";
					when "01001100010101011" => rgb <= "101000";
					when "01001100010101100" => rgb <= "101000";
					when "01001100010101101" => rgb <= "101000";
					when "01001100010101110" => rgb <= "101000";
					when "01001100010101111" => rgb <= "101000";
					when "01001100010110000" => rgb <= "101000";
					when "01001100010110001" => rgb <= "101000";
					when "01001100010110010" => rgb <= "101000";
					when "01001100010110011" => rgb <= "101000";
					when "01001100010110100" => rgb <= "101000";
					when "01001100010110101" => rgb <= "010100";
					when "01001100010110110" => rgb <= "000000";
					when "01001100010110111" => rgb <= "000000";
					when "01001100010111000" => rgb <= "000000";
					when "01001100010111001" => rgb <= "000000";
					when "01001100010111010" => rgb <= "000000";
					when "01001100010111011" => rgb <= "000000";
					when "01001100010111100" => rgb <= "000000";
					when "01001100010111101" => rgb <= "000000";
					when "01001100010111110" => rgb <= "000000";
					when "01001100010111111" => rgb <= "000000";
					when "01001100011000000" => rgb <= "000000";
					when "01001100011000001" => rgb <= "000000";
					when "01001100011000010" => rgb <= "000000";
					when "01001100011000011" => rgb <= "000000";
					when "01001100011000100" => rgb <= "000000";
					when "01001100011000101" => rgb <= "000000";
					when "01001100011000110" => rgb <= "000000";
					when "01001100011000111" => rgb <= "000000";
					when "01001100011001000" => rgb <= "000000";
					when "01001100011001001" => rgb <= "000000";
					when "01001100011001010" => rgb <= "000000";
					when "01001100011001011" => rgb <= "000000";
					when "01001100011001100" => rgb <= "000000";
					when "01001100011001101" => rgb <= "000000";
					when "01001100011001110" => rgb <= "000000";
					when "01001100011001111" => rgb <= "000000";
					when "01001100011010000" => rgb <= "000000";
					when "01001100011010001" => rgb <= "000000";
					when "01001100011010010" => rgb <= "000000";
					when "01001100011010011" => rgb <= "000000";
					when "01001100011010100" => rgb <= "000000";
					when "01001100011010101" => rgb <= "000000";
					when "01001100011010110" => rgb <= "000000";
					when "01001100011010111" => rgb <= "000000";
					when "01001100011011000" => rgb <= "000000";
					when "01001100011011001" => rgb <= "000000";
					when "01001100011011010" => rgb <= "000000";
					when "01001100011011011" => rgb <= "000000";
					when "01001100011011100" => rgb <= "000000";
					when "01001100011011101" => rgb <= "000000";
					when "01001100011011110" => rgb <= "000000";
					when "01001100011011111" => rgb <= "000000";
					when "01001100011100000" => rgb <= "000000";
					when "01001100011100001" => rgb <= "000000";
					when "01001100011100010" => rgb <= "000000";
					when "01001100011100011" => rgb <= "000000";
					when "01001100011100100" => rgb <= "000000";
					when "01001100011100101" => rgb <= "000000";
					when "01001100011100110" => rgb <= "000000";
					when "01001100011100111" => rgb <= "000000";
					when "01001100011101000" => rgb <= "000000";
					when "01001100011101001" => rgb <= "000000";
					when "01001100011101010" => rgb <= "000000";
					when "01001100011101011" => rgb <= "000000";
					when "01001100011101100" => rgb <= "000000";
					when "01001100011101101" => rgb <= "000000";
					when "01001100011101110" => rgb <= "000000";
					when "01001100011101111" => rgb <= "000000";
					when "01001100011110000" => rgb <= "000000";
					when "01001100011110001" => rgb <= "000000";
					when "01001100011110010" => rgb <= "000000";
					when "01001100011110011" => rgb <= "000000";
					when "01001100011110100" => rgb <= "000000";
					when "01001100011110101" => rgb <= "000000";
					when "01001100011110110" => rgb <= "000000";
					when "01001100011110111" => rgb <= "000000";
					when "01001100011111000" => rgb <= "000000";
					when "01001100011111001" => rgb <= "000000";
					when "01001100011111010" => rgb <= "000000";
					when "01001100011111011" => rgb <= "000000";
					when "01001100011111100" => rgb <= "000000";
					when "01001100011111101" => rgb <= "000000";
					when "01001100011111110" => rgb <= "000000";
					when "01001100011111111" => rgb <= "000000";
					when "01001100100000000" => rgb <= "000000";
					when "01001100100000001" => rgb <= "000000";
					when "01001100100000010" => rgb <= "000000";
					when "01001100100000011" => rgb <= "000000";
					when "01001100100000100" => rgb <= "000000";
					when "01001100100000101" => rgb <= "000000";
					when "01001100100000110" => rgb <= "000000";
					when "01001100100000111" => rgb <= "000000";
					when "01001100100001000" => rgb <= "000000";
					when "01001100100001001" => rgb <= "000000";
					when "01001100100001010" => rgb <= "000000";
					when "01001100100001011" => rgb <= "000000";
					when "01001100100001100" => rgb <= "000000";
					when "01001100100001101" => rgb <= "000000";
					when "01001100100001110" => rgb <= "000000";
					when "01001100100001111" => rgb <= "000000";
					when "01001100100010000" => rgb <= "000000";
					when "01001100100010001" => rgb <= "000000";
					when "01001100100010010" => rgb <= "000000";
					when "01001100100010011" => rgb <= "000000";
					when "01001100100010100" => rgb <= "000000";
					when "01001100100010101" => rgb <= "000000";
					when "01001100100010110" => rgb <= "000000";
					when "01001100100010111" => rgb <= "000000";
					when "01001100100011000" => rgb <= "000000";
					when "01001100100011001" => rgb <= "000000";
					when "01001100100011010" => rgb <= "000000";
					when "01001100100011011" => rgb <= "000000";
					when "01001100100011100" => rgb <= "000000";
					when "01001100100011101" => rgb <= "000000";
					when "01001100100011110" => rgb <= "000000";
					when "01001100100011111" => rgb <= "000000";
					when "01001100100100000" => rgb <= "000000";
					when "01001100100100001" => rgb <= "000000";
					when "01001100100100010" => rgb <= "000000";
					when "01001100100100011" => rgb <= "000000";
					when "01001100100100100" => rgb <= "000000";
					when "01001100100100101" => rgb <= "000000";
					when "01001100100100110" => rgb <= "000000";
					when "01001100100100111" => rgb <= "000000";
					when "01001100100101000" => rgb <= "000000";
					when "01001100100101001" => rgb <= "000000";
					when "01001100100101010" => rgb <= "000000";
					when "01001100100101011" => rgb <= "000000";
					when "01001100100101100" => rgb <= "000000";
					when "01001100100101101" => rgb <= "000000";
					when "01001100100101110" => rgb <= "000000";
					when "01001100100101111" => rgb <= "000000";
					when "01001100100110000" => rgb <= "000000";
					when "01001100100110001" => rgb <= "000000";
					when "01001100100110010" => rgb <= "000000";
					when "01001100100110011" => rgb <= "000000";
					when "01001100100110100" => rgb <= "000000";
					when "01001100100110101" => rgb <= "000000";
					when "01001100100110110" => rgb <= "000000";
					when "01001100100110111" => rgb <= "000000";
					when "01001100100111000" => rgb <= "000000";
					when "01001100100111001" => rgb <= "000000";
					when "01001100100111010" => rgb <= "000000";
					when "01001100100111011" => rgb <= "000000";
					when "01001100100111100" => rgb <= "000000";
					when "01001100100111101" => rgb <= "000000";
					when "01001100100111110" => rgb <= "000000";
					when "01001100100111111" => rgb <= "000000";
					when "01001101000000000" => rgb <= "000000";
					when "01001101000000001" => rgb <= "000000";
					when "01001101000000010" => rgb <= "000000";
					when "01001101000000011" => rgb <= "000000";
					when "01001101000000100" => rgb <= "000000";
					when "01001101000000101" => rgb <= "000000";
					when "01001101000000110" => rgb <= "000000";
					when "01001101000000111" => rgb <= "000000";
					when "01001101000001000" => rgb <= "000000";
					when "01001101000001001" => rgb <= "000000";
					when "01001101000001010" => rgb <= "000000";
					when "01001101000001011" => rgb <= "000000";
					when "01001101000001100" => rgb <= "000000";
					when "01001101000001101" => rgb <= "000000";
					when "01001101000001110" => rgb <= "000000";
					when "01001101000001111" => rgb <= "000000";
					when "01001101000010000" => rgb <= "000000";
					when "01001101000010001" => rgb <= "000000";
					when "01001101000010010" => rgb <= "000000";
					when "01001101000010011" => rgb <= "000000";
					when "01001101000010100" => rgb <= "000000";
					when "01001101000010101" => rgb <= "000000";
					when "01001101000010110" => rgb <= "000000";
					when "01001101000010111" => rgb <= "000000";
					when "01001101000011000" => rgb <= "000000";
					when "01001101000011001" => rgb <= "000000";
					when "01001101000011010" => rgb <= "000000";
					when "01001101000011011" => rgb <= "000000";
					when "01001101000011100" => rgb <= "000000";
					when "01001101000011101" => rgb <= "000000";
					when "01001101000011110" => rgb <= "000000";
					when "01001101000011111" => rgb <= "000000";
					when "01001101000100000" => rgb <= "000000";
					when "01001101000100001" => rgb <= "000000";
					when "01001101000100010" => rgb <= "000000";
					when "01001101000100011" => rgb <= "000000";
					when "01001101000100100" => rgb <= "000000";
					when "01001101000100101" => rgb <= "000000";
					when "01001101000100110" => rgb <= "000000";
					when "01001101000100111" => rgb <= "000000";
					when "01001101000101000" => rgb <= "000000";
					when "01001101000101001" => rgb <= "000000";
					when "01001101000101010" => rgb <= "000000";
					when "01001101000101011" => rgb <= "000000";
					when "01001101000101100" => rgb <= "000000";
					when "01001101000101101" => rgb <= "000000";
					when "01001101000101110" => rgb <= "000000";
					when "01001101000101111" => rgb <= "000000";
					when "01001101000110000" => rgb <= "000000";
					when "01001101000110001" => rgb <= "000000";
					when "01001101000110010" => rgb <= "000000";
					when "01001101000110011" => rgb <= "000000";
					when "01001101000110100" => rgb <= "000000";
					when "01001101000110101" => rgb <= "000000";
					when "01001101000110110" => rgb <= "000000";
					when "01001101000110111" => rgb <= "000000";
					when "01001101000111000" => rgb <= "000000";
					when "01001101000111001" => rgb <= "000000";
					when "01001101000111010" => rgb <= "000000";
					when "01001101000111011" => rgb <= "000000";
					when "01001101000111100" => rgb <= "000000";
					when "01001101000111101" => rgb <= "000000";
					when "01001101000111110" => rgb <= "000000";
					when "01001101000111111" => rgb <= "000000";
					when "01001101001000000" => rgb <= "000000";
					when "01001101001000001" => rgb <= "000000";
					when "01001101001000010" => rgb <= "000000";
					when "01001101001000011" => rgb <= "000000";
					when "01001101001000100" => rgb <= "000000";
					when "01001101001000101" => rgb <= "000000";
					when "01001101001000110" => rgb <= "000000";
					when "01001101001000111" => rgb <= "000000";
					when "01001101001001000" => rgb <= "000000";
					when "01001101001001001" => rgb <= "000000";
					when "01001101001001010" => rgb <= "000000";
					when "01001101001001011" => rgb <= "000000";
					when "01001101001001100" => rgb <= "000000";
					when "01001101001001101" => rgb <= "000000";
					when "01001101001001110" => rgb <= "000000";
					when "01001101001001111" => rgb <= "000000";
					when "01001101001010000" => rgb <= "000000";
					when "01001101001010001" => rgb <= "000000";
					when "01001101001010010" => rgb <= "000000";
					when "01001101001010011" => rgb <= "000000";
					when "01001101001010100" => rgb <= "000000";
					when "01001101001010101" => rgb <= "000000";
					when "01001101001010110" => rgb <= "000000";
					when "01001101001010111" => rgb <= "000000";
					when "01001101001011000" => rgb <= "000000";
					when "01001101001011001" => rgb <= "000000";
					when "01001101001011010" => rgb <= "000000";
					when "01001101001011011" => rgb <= "000000";
					when "01001101001011100" => rgb <= "000000";
					when "01001101001011101" => rgb <= "000000";
					when "01001101001011110" => rgb <= "000000";
					when "01001101001011111" => rgb <= "000000";
					when "01001101001100000" => rgb <= "000000";
					when "01001101001100001" => rgb <= "000000";
					when "01001101001100010" => rgb <= "000000";
					when "01001101001100011" => rgb <= "000000";
					when "01001101001100100" => rgb <= "000000";
					when "01001101001100101" => rgb <= "000000";
					when "01001101001100110" => rgb <= "000000";
					when "01001101001100111" => rgb <= "000000";
					when "01001101001101000" => rgb <= "000000";
					when "01001101001101001" => rgb <= "000000";
					when "01001101001101010" => rgb <= "000000";
					when "01001101001101011" => rgb <= "000000";
					when "01001101001101100" => rgb <= "000000";
					when "01001101001101101" => rgb <= "000000";
					when "01001101001101110" => rgb <= "000000";
					when "01001101001101111" => rgb <= "000000";
					when "01001101001110000" => rgb <= "000000";
					when "01001101001110001" => rgb <= "000000";
					when "01001101001110010" => rgb <= "000000";
					when "01001101001110011" => rgb <= "000000";
					when "01001101001110100" => rgb <= "000000";
					when "01001101001110101" => rgb <= "000000";
					when "01001101001110110" => rgb <= "000000";
					when "01001101001110111" => rgb <= "000000";
					when "01001101001111000" => rgb <= "000000";
					when "01001101001111001" => rgb <= "000000";
					when "01001101001111010" => rgb <= "000000";
					when "01001101001111011" => rgb <= "000000";
					when "01001101001111100" => rgb <= "000000";
					when "01001101001111101" => rgb <= "000000";
					when "01001101001111110" => rgb <= "000000";
					when "01001101001111111" => rgb <= "000000";
					when "01001101010000000" => rgb <= "000000";
					when "01001101010000001" => rgb <= "000000";
					when "01001101010000010" => rgb <= "000000";
					when "01001101010000011" => rgb <= "000000";
					when "01001101010000100" => rgb <= "000000";
					when "01001101010000101" => rgb <= "000000";
					when "01001101010000110" => rgb <= "000000";
					when "01001101010000111" => rgb <= "000000";
					when "01001101010001000" => rgb <= "100100";
					when "01001101010001001" => rgb <= "101000";
					when "01001101010001010" => rgb <= "101000";
					when "01001101010001011" => rgb <= "101000";
					when "01001101010001100" => rgb <= "101000";
					when "01001101010001101" => rgb <= "101000";
					when "01001101010001110" => rgb <= "101000";
					when "01001101010001111" => rgb <= "101000";
					when "01001101010010000" => rgb <= "101000";
					when "01001101010010001" => rgb <= "101000";
					when "01001101010010010" => rgb <= "101000";
					when "01001101010010011" => rgb <= "101000";
					when "01001101010010100" => rgb <= "101000";
					when "01001101010010101" => rgb <= "101000";
					when "01001101010010110" => rgb <= "101000";
					when "01001101010010111" => rgb <= "101000";
					when "01001101010011000" => rgb <= "101000";
					when "01001101010011001" => rgb <= "101000";
					when "01001101010011010" => rgb <= "101000";
					when "01001101010011011" => rgb <= "101000";
					when "01001101010011100" => rgb <= "101000";
					when "01001101010011101" => rgb <= "101000";
					when "01001101010011110" => rgb <= "101000";
					when "01001101010011111" => rgb <= "101000";
					when "01001101010100000" => rgb <= "101000";
					when "01001101010100001" => rgb <= "101000";
					when "01001101010100010" => rgb <= "101000";
					when "01001101010100011" => rgb <= "101000";
					when "01001101010100100" => rgb <= "101000";
					when "01001101010100101" => rgb <= "101000";
					when "01001101010100110" => rgb <= "101000";
					when "01001101010100111" => rgb <= "101000";
					when "01001101010101000" => rgb <= "101000";
					when "01001101010101001" => rgb <= "101000";
					when "01001101010101010" => rgb <= "101000";
					when "01001101010101011" => rgb <= "101000";
					when "01001101010101100" => rgb <= "101000";
					when "01001101010101101" => rgb <= "101000";
					when "01001101010101110" => rgb <= "101000";
					when "01001101010101111" => rgb <= "101000";
					when "01001101010110000" => rgb <= "101000";
					when "01001101010110001" => rgb <= "101000";
					when "01001101010110010" => rgb <= "101000";
					when "01001101010110011" => rgb <= "101000";
					when "01001101010110100" => rgb <= "101000";
					when "01001101010110101" => rgb <= "010100";
					when "01001101010110110" => rgb <= "000000";
					when "01001101010110111" => rgb <= "000000";
					when "01001101010111000" => rgb <= "000000";
					when "01001101010111001" => rgb <= "000000";
					when "01001101010111010" => rgb <= "000000";
					when "01001101010111011" => rgb <= "000000";
					when "01001101010111100" => rgb <= "000000";
					when "01001101010111101" => rgb <= "000000";
					when "01001101010111110" => rgb <= "000000";
					when "01001101010111111" => rgb <= "000000";
					when "01001101011000000" => rgb <= "000000";
					when "01001101011000001" => rgb <= "000000";
					when "01001101011000010" => rgb <= "000000";
					when "01001101011000011" => rgb <= "000000";
					when "01001101011000100" => rgb <= "000000";
					when "01001101011000101" => rgb <= "000000";
					when "01001101011000110" => rgb <= "000000";
					when "01001101011000111" => rgb <= "000000";
					when "01001101011001000" => rgb <= "000000";
					when "01001101011001001" => rgb <= "000000";
					when "01001101011001010" => rgb <= "000000";
					when "01001101011001011" => rgb <= "000000";
					when "01001101011001100" => rgb <= "000000";
					when "01001101011001101" => rgb <= "000000";
					when "01001101011001110" => rgb <= "000000";
					when "01001101011001111" => rgb <= "000000";
					when "01001101011010000" => rgb <= "000000";
					when "01001101011010001" => rgb <= "000000";
					when "01001101011010010" => rgb <= "000000";
					when "01001101011010011" => rgb <= "000000";
					when "01001101011010100" => rgb <= "000000";
					when "01001101011010101" => rgb <= "000000";
					when "01001101011010110" => rgb <= "000000";
					when "01001101011010111" => rgb <= "000000";
					when "01001101011011000" => rgb <= "000000";
					when "01001101011011001" => rgb <= "000000";
					when "01001101011011010" => rgb <= "000000";
					when "01001101011011011" => rgb <= "000000";
					when "01001101011011100" => rgb <= "000000";
					when "01001101011011101" => rgb <= "000000";
					when "01001101011011110" => rgb <= "000000";
					when "01001101011011111" => rgb <= "000000";
					when "01001101011100000" => rgb <= "000000";
					when "01001101011100001" => rgb <= "000000";
					when "01001101011100010" => rgb <= "000000";
					when "01001101011100011" => rgb <= "000000";
					when "01001101011100100" => rgb <= "000000";
					when "01001101011100101" => rgb <= "000000";
					when "01001101011100110" => rgb <= "000000";
					when "01001101011100111" => rgb <= "000000";
					when "01001101011101000" => rgb <= "000000";
					when "01001101011101001" => rgb <= "000000";
					when "01001101011101010" => rgb <= "000000";
					when "01001101011101011" => rgb <= "000000";
					when "01001101011101100" => rgb <= "000000";
					when "01001101011101101" => rgb <= "000000";
					when "01001101011101110" => rgb <= "000000";
					when "01001101011101111" => rgb <= "000000";
					when "01001101011110000" => rgb <= "000000";
					when "01001101011110001" => rgb <= "000000";
					when "01001101011110010" => rgb <= "000000";
					when "01001101011110011" => rgb <= "000000";
					when "01001101011110100" => rgb <= "000000";
					when "01001101011110101" => rgb <= "000000";
					when "01001101011110110" => rgb <= "000000";
					when "01001101011110111" => rgb <= "000000";
					when "01001101011111000" => rgb <= "000000";
					when "01001101011111001" => rgb <= "000000";
					when "01001101011111010" => rgb <= "000000";
					when "01001101011111011" => rgb <= "000000";
					when "01001101011111100" => rgb <= "000000";
					when "01001101011111101" => rgb <= "000000";
					when "01001101011111110" => rgb <= "000000";
					when "01001101011111111" => rgb <= "000000";
					when "01001101100000000" => rgb <= "000000";
					when "01001101100000001" => rgb <= "000000";
					when "01001101100000010" => rgb <= "000000";
					when "01001101100000011" => rgb <= "000000";
					when "01001101100000100" => rgb <= "000000";
					when "01001101100000101" => rgb <= "000000";
					when "01001101100000110" => rgb <= "000000";
					when "01001101100000111" => rgb <= "000000";
					when "01001101100001000" => rgb <= "000000";
					when "01001101100001001" => rgb <= "000000";
					when "01001101100001010" => rgb <= "000000";
					when "01001101100001011" => rgb <= "000000";
					when "01001101100001100" => rgb <= "000000";
					when "01001101100001101" => rgb <= "000000";
					when "01001101100001110" => rgb <= "000000";
					when "01001101100001111" => rgb <= "000000";
					when "01001101100010000" => rgb <= "000000";
					when "01001101100010001" => rgb <= "000000";
					when "01001101100010010" => rgb <= "000000";
					when "01001101100010011" => rgb <= "000000";
					when "01001101100010100" => rgb <= "000000";
					when "01001101100010101" => rgb <= "000000";
					when "01001101100010110" => rgb <= "000000";
					when "01001101100010111" => rgb <= "000000";
					when "01001101100011000" => rgb <= "000000";
					when "01001101100011001" => rgb <= "000000";
					when "01001101100011010" => rgb <= "000000";
					when "01001101100011011" => rgb <= "000000";
					when "01001101100011100" => rgb <= "000000";
					when "01001101100011101" => rgb <= "000000";
					when "01001101100011110" => rgb <= "000000";
					when "01001101100011111" => rgb <= "000000";
					when "01001101100100000" => rgb <= "000000";
					when "01001101100100001" => rgb <= "000000";
					when "01001101100100010" => rgb <= "000000";
					when "01001101100100011" => rgb <= "000000";
					when "01001101100100100" => rgb <= "000000";
					when "01001101100100101" => rgb <= "000000";
					when "01001101100100110" => rgb <= "000000";
					when "01001101100100111" => rgb <= "000000";
					when "01001101100101000" => rgb <= "000000";
					when "01001101100101001" => rgb <= "000000";
					when "01001101100101010" => rgb <= "000000";
					when "01001101100101011" => rgb <= "000000";
					when "01001101100101100" => rgb <= "000000";
					when "01001101100101101" => rgb <= "000000";
					when "01001101100101110" => rgb <= "000000";
					when "01001101100101111" => rgb <= "000000";
					when "01001101100110000" => rgb <= "000000";
					when "01001101100110001" => rgb <= "000000";
					when "01001101100110010" => rgb <= "000000";
					when "01001101100110011" => rgb <= "000000";
					when "01001101100110100" => rgb <= "000000";
					when "01001101100110101" => rgb <= "000000";
					when "01001101100110110" => rgb <= "000000";
					when "01001101100110111" => rgb <= "000000";
					when "01001101100111000" => rgb <= "000000";
					when "01001101100111001" => rgb <= "000000";
					when "01001101100111010" => rgb <= "000000";
					when "01001101100111011" => rgb <= "000000";
					when "01001101100111100" => rgb <= "000000";
					when "01001101100111101" => rgb <= "000000";
					when "01001101100111110" => rgb <= "000000";
					when "01001101100111111" => rgb <= "000000";
					when "01001110000000000" => rgb <= "000000";
					when "01001110000000001" => rgb <= "000000";
					when "01001110000000010" => rgb <= "000000";
					when "01001110000000011" => rgb <= "000000";
					when "01001110000000100" => rgb <= "000000";
					when "01001110000000101" => rgb <= "000000";
					when "01001110000000110" => rgb <= "000000";
					when "01001110000000111" => rgb <= "000000";
					when "01001110000001000" => rgb <= "000000";
					when "01001110000001001" => rgb <= "000000";
					when "01001110000001010" => rgb <= "000000";
					when "01001110000001011" => rgb <= "000000";
					when "01001110000001100" => rgb <= "000000";
					when "01001110000001101" => rgb <= "000000";
					when "01001110000001110" => rgb <= "000000";
					when "01001110000001111" => rgb <= "000000";
					when "01001110000010000" => rgb <= "000000";
					when "01001110000010001" => rgb <= "000000";
					when "01001110000010010" => rgb <= "000000";
					when "01001110000010011" => rgb <= "000000";
					when "01001110000010100" => rgb <= "000000";
					when "01001110000010101" => rgb <= "000000";
					when "01001110000010110" => rgb <= "000000";
					when "01001110000010111" => rgb <= "000000";
					when "01001110000011000" => rgb <= "000000";
					when "01001110000011001" => rgb <= "000000";
					when "01001110000011010" => rgb <= "000000";
					when "01001110000011011" => rgb <= "000000";
					when "01001110000011100" => rgb <= "000000";
					when "01001110000011101" => rgb <= "000000";
					when "01001110000011110" => rgb <= "000000";
					when "01001110000011111" => rgb <= "000000";
					when "01001110000100000" => rgb <= "000000";
					when "01001110000100001" => rgb <= "000000";
					when "01001110000100010" => rgb <= "000000";
					when "01001110000100011" => rgb <= "000000";
					when "01001110000100100" => rgb <= "000000";
					when "01001110000100101" => rgb <= "000000";
					when "01001110000100110" => rgb <= "000000";
					when "01001110000100111" => rgb <= "000000";
					when "01001110000101000" => rgb <= "000000";
					when "01001110000101001" => rgb <= "000000";
					when "01001110000101010" => rgb <= "000000";
					when "01001110000101011" => rgb <= "000000";
					when "01001110000101100" => rgb <= "000000";
					when "01001110000101101" => rgb <= "000000";
					when "01001110000101110" => rgb <= "000000";
					when "01001110000101111" => rgb <= "000000";
					when "01001110000110000" => rgb <= "000000";
					when "01001110000110001" => rgb <= "000000";
					when "01001110000110010" => rgb <= "000000";
					when "01001110000110011" => rgb <= "000000";
					when "01001110000110100" => rgb <= "000000";
					when "01001110000110101" => rgb <= "000000";
					when "01001110000110110" => rgb <= "000000";
					when "01001110000110111" => rgb <= "000000";
					when "01001110000111000" => rgb <= "000000";
					when "01001110000111001" => rgb <= "000000";
					when "01001110000111010" => rgb <= "000000";
					when "01001110000111011" => rgb <= "000000";
					when "01001110000111100" => rgb <= "000000";
					when "01001110000111101" => rgb <= "000000";
					when "01001110000111110" => rgb <= "000000";
					when "01001110000111111" => rgb <= "000000";
					when "01001110001000000" => rgb <= "000000";
					when "01001110001000001" => rgb <= "000000";
					when "01001110001000010" => rgb <= "000000";
					when "01001110001000011" => rgb <= "000000";
					when "01001110001000100" => rgb <= "000000";
					when "01001110001000101" => rgb <= "000000";
					when "01001110001000110" => rgb <= "000000";
					when "01001110001000111" => rgb <= "000000";
					when "01001110001001000" => rgb <= "000000";
					when "01001110001001001" => rgb <= "000000";
					when "01001110001001010" => rgb <= "000000";
					when "01001110001001011" => rgb <= "000000";
					when "01001110001001100" => rgb <= "000000";
					when "01001110001001101" => rgb <= "000000";
					when "01001110001001110" => rgb <= "000000";
					when "01001110001001111" => rgb <= "000000";
					when "01001110001010000" => rgb <= "000000";
					when "01001110001010001" => rgb <= "000000";
					when "01001110001010010" => rgb <= "000000";
					when "01001110001010011" => rgb <= "000000";
					when "01001110001010100" => rgb <= "000000";
					when "01001110001010101" => rgb <= "000000";
					when "01001110001010110" => rgb <= "000000";
					when "01001110001010111" => rgb <= "000000";
					when "01001110001011000" => rgb <= "000000";
					when "01001110001011001" => rgb <= "000000";
					when "01001110001011010" => rgb <= "000000";
					when "01001110001011011" => rgb <= "000000";
					when "01001110001011100" => rgb <= "000000";
					when "01001110001011101" => rgb <= "000000";
					when "01001110001011110" => rgb <= "000000";
					when "01001110001011111" => rgb <= "000000";
					when "01001110001100000" => rgb <= "000000";
					when "01001110001100001" => rgb <= "000000";
					when "01001110001100010" => rgb <= "000000";
					when "01001110001100011" => rgb <= "000000";
					when "01001110001100100" => rgb <= "000000";
					when "01001110001100101" => rgb <= "000000";
					when "01001110001100110" => rgb <= "000000";
					when "01001110001100111" => rgb <= "000000";
					when "01001110001101000" => rgb <= "000000";
					when "01001110001101001" => rgb <= "000000";
					when "01001110001101010" => rgb <= "000000";
					when "01001110001101011" => rgb <= "000000";
					when "01001110001101100" => rgb <= "000000";
					when "01001110001101101" => rgb <= "000000";
					when "01001110001101110" => rgb <= "000000";
					when "01001110001101111" => rgb <= "000000";
					when "01001110001110000" => rgb <= "000000";
					when "01001110001110001" => rgb <= "000000";
					when "01001110001110010" => rgb <= "000000";
					when "01001110001110011" => rgb <= "000000";
					when "01001110001110100" => rgb <= "000000";
					when "01001110001110101" => rgb <= "000000";
					when "01001110001110110" => rgb <= "000000";
					when "01001110001110111" => rgb <= "000000";
					when "01001110001111000" => rgb <= "000000";
					when "01001110001111001" => rgb <= "000000";
					when "01001110001111010" => rgb <= "000000";
					when "01001110001111011" => rgb <= "000000";
					when "01001110001111100" => rgb <= "000000";
					when "01001110001111101" => rgb <= "000000";
					when "01001110001111110" => rgb <= "000000";
					when "01001110001111111" => rgb <= "000000";
					when "01001110010000000" => rgb <= "000000";
					when "01001110010000001" => rgb <= "000000";
					when "01001110010000010" => rgb <= "000000";
					when "01001110010000011" => rgb <= "000000";
					when "01001110010000100" => rgb <= "000000";
					when "01001110010000101" => rgb <= "000000";
					when "01001110010000110" => rgb <= "000000";
					when "01001110010000111" => rgb <= "000000";
					when "01001110010001000" => rgb <= "100100";
					when "01001110010001001" => rgb <= "101000";
					when "01001110010001010" => rgb <= "101000";
					when "01001110010001011" => rgb <= "101000";
					when "01001110010001100" => rgb <= "101000";
					when "01001110010001101" => rgb <= "101000";
					when "01001110010001110" => rgb <= "101000";
					when "01001110010001111" => rgb <= "101000";
					when "01001110010010000" => rgb <= "101000";
					when "01001110010010001" => rgb <= "101000";
					when "01001110010010010" => rgb <= "101000";
					when "01001110010010011" => rgb <= "101000";
					when "01001110010010100" => rgb <= "101000";
					when "01001110010010101" => rgb <= "101000";
					when "01001110010010110" => rgb <= "101000";
					when "01001110010010111" => rgb <= "101000";
					when "01001110010011000" => rgb <= "101000";
					when "01001110010011001" => rgb <= "101000";
					when "01001110010011010" => rgb <= "101000";
					when "01001110010011011" => rgb <= "101000";
					when "01001110010011100" => rgb <= "101000";
					when "01001110010011101" => rgb <= "101000";
					when "01001110010011110" => rgb <= "101000";
					when "01001110010011111" => rgb <= "101000";
					when "01001110010100000" => rgb <= "101000";
					when "01001110010100001" => rgb <= "101000";
					when "01001110010100010" => rgb <= "101000";
					when "01001110010100011" => rgb <= "101000";
					when "01001110010100100" => rgb <= "101000";
					when "01001110010100101" => rgb <= "101000";
					when "01001110010100110" => rgb <= "101000";
					when "01001110010100111" => rgb <= "101000";
					when "01001110010101000" => rgb <= "101000";
					when "01001110010101001" => rgb <= "101000";
					when "01001110010101010" => rgb <= "101000";
					when "01001110010101011" => rgb <= "101000";
					when "01001110010101100" => rgb <= "101000";
					when "01001110010101101" => rgb <= "101000";
					when "01001110010101110" => rgb <= "101000";
					when "01001110010101111" => rgb <= "101000";
					when "01001110010110000" => rgb <= "101000";
					when "01001110010110001" => rgb <= "101000";
					when "01001110010110010" => rgb <= "101000";
					when "01001110010110011" => rgb <= "101000";
					when "01001110010110100" => rgb <= "101000";
					when "01001110010110101" => rgb <= "010100";
					when "01001110010110110" => rgb <= "000000";
					when "01001110010110111" => rgb <= "000000";
					when "01001110010111000" => rgb <= "000000";
					when "01001110010111001" => rgb <= "000000";
					when "01001110010111010" => rgb <= "000000";
					when "01001110010111011" => rgb <= "000000";
					when "01001110010111100" => rgb <= "000000";
					when "01001110010111101" => rgb <= "000000";
					when "01001110010111110" => rgb <= "000000";
					when "01001110010111111" => rgb <= "000000";
					when "01001110011000000" => rgb <= "000000";
					when "01001110011000001" => rgb <= "000000";
					when "01001110011000010" => rgb <= "000000";
					when "01001110011000011" => rgb <= "000000";
					when "01001110011000100" => rgb <= "000000";
					when "01001110011000101" => rgb <= "000000";
					when "01001110011000110" => rgb <= "000000";
					when "01001110011000111" => rgb <= "000000";
					when "01001110011001000" => rgb <= "000000";
					when "01001110011001001" => rgb <= "000000";
					when "01001110011001010" => rgb <= "000000";
					when "01001110011001011" => rgb <= "000000";
					when "01001110011001100" => rgb <= "000000";
					when "01001110011001101" => rgb <= "000000";
					when "01001110011001110" => rgb <= "000000";
					when "01001110011001111" => rgb <= "000000";
					when "01001110011010000" => rgb <= "000000";
					when "01001110011010001" => rgb <= "000000";
					when "01001110011010010" => rgb <= "000000";
					when "01001110011010011" => rgb <= "000000";
					when "01001110011010100" => rgb <= "000000";
					when "01001110011010101" => rgb <= "000000";
					when "01001110011010110" => rgb <= "000000";
					when "01001110011010111" => rgb <= "000000";
					when "01001110011011000" => rgb <= "000000";
					when "01001110011011001" => rgb <= "000000";
					when "01001110011011010" => rgb <= "000000";
					when "01001110011011011" => rgb <= "000000";
					when "01001110011011100" => rgb <= "000000";
					when "01001110011011101" => rgb <= "000000";
					when "01001110011011110" => rgb <= "000000";
					when "01001110011011111" => rgb <= "000000";
					when "01001110011100000" => rgb <= "000000";
					when "01001110011100001" => rgb <= "000000";
					when "01001110011100010" => rgb <= "000000";
					when "01001110011100011" => rgb <= "000000";
					when "01001110011100100" => rgb <= "000000";
					when "01001110011100101" => rgb <= "000000";
					when "01001110011100110" => rgb <= "000000";
					when "01001110011100111" => rgb <= "000000";
					when "01001110011101000" => rgb <= "000000";
					when "01001110011101001" => rgb <= "000000";
					when "01001110011101010" => rgb <= "000000";
					when "01001110011101011" => rgb <= "000000";
					when "01001110011101100" => rgb <= "000000";
					when "01001110011101101" => rgb <= "000000";
					when "01001110011101110" => rgb <= "000000";
					when "01001110011101111" => rgb <= "000000";
					when "01001110011110000" => rgb <= "000000";
					when "01001110011110001" => rgb <= "000000";
					when "01001110011110010" => rgb <= "000000";
					when "01001110011110011" => rgb <= "000000";
					when "01001110011110100" => rgb <= "000000";
					when "01001110011110101" => rgb <= "000000";
					when "01001110011110110" => rgb <= "000000";
					when "01001110011110111" => rgb <= "000000";
					when "01001110011111000" => rgb <= "000000";
					when "01001110011111001" => rgb <= "000000";
					when "01001110011111010" => rgb <= "000000";
					when "01001110011111011" => rgb <= "000000";
					when "01001110011111100" => rgb <= "000000";
					when "01001110011111101" => rgb <= "000000";
					when "01001110011111110" => rgb <= "000000";
					when "01001110011111111" => rgb <= "000000";
					when "01001110100000000" => rgb <= "000000";
					when "01001110100000001" => rgb <= "000000";
					when "01001110100000010" => rgb <= "000000";
					when "01001110100000011" => rgb <= "000000";
					when "01001110100000100" => rgb <= "000000";
					when "01001110100000101" => rgb <= "000000";
					when "01001110100000110" => rgb <= "000000";
					when "01001110100000111" => rgb <= "000000";
					when "01001110100001000" => rgb <= "000000";
					when "01001110100001001" => rgb <= "000000";
					when "01001110100001010" => rgb <= "000000";
					when "01001110100001011" => rgb <= "000000";
					when "01001110100001100" => rgb <= "000000";
					when "01001110100001101" => rgb <= "000000";
					when "01001110100001110" => rgb <= "000000";
					when "01001110100001111" => rgb <= "000000";
					when "01001110100010000" => rgb <= "000000";
					when "01001110100010001" => rgb <= "000000";
					when "01001110100010010" => rgb <= "000000";
					when "01001110100010011" => rgb <= "000000";
					when "01001110100010100" => rgb <= "000000";
					when "01001110100010101" => rgb <= "000000";
					when "01001110100010110" => rgb <= "000000";
					when "01001110100010111" => rgb <= "000000";
					when "01001110100011000" => rgb <= "000000";
					when "01001110100011001" => rgb <= "000000";
					when "01001110100011010" => rgb <= "000000";
					when "01001110100011011" => rgb <= "000000";
					when "01001110100011100" => rgb <= "000000";
					when "01001110100011101" => rgb <= "000000";
					when "01001110100011110" => rgb <= "000000";
					when "01001110100011111" => rgb <= "000000";
					when "01001110100100000" => rgb <= "000000";
					when "01001110100100001" => rgb <= "000000";
					when "01001110100100010" => rgb <= "000000";
					when "01001110100100011" => rgb <= "000000";
					when "01001110100100100" => rgb <= "000000";
					when "01001110100100101" => rgb <= "000000";
					when "01001110100100110" => rgb <= "000000";
					when "01001110100100111" => rgb <= "000000";
					when "01001110100101000" => rgb <= "000000";
					when "01001110100101001" => rgb <= "000000";
					when "01001110100101010" => rgb <= "000000";
					when "01001110100101011" => rgb <= "000000";
					when "01001110100101100" => rgb <= "000000";
					when "01001110100101101" => rgb <= "000000";
					when "01001110100101110" => rgb <= "000000";
					when "01001110100101111" => rgb <= "000000";
					when "01001110100110000" => rgb <= "000000";
					when "01001110100110001" => rgb <= "000000";
					when "01001110100110010" => rgb <= "000000";
					when "01001110100110011" => rgb <= "000000";
					when "01001110100110100" => rgb <= "000000";
					when "01001110100110101" => rgb <= "000000";
					when "01001110100110110" => rgb <= "000000";
					when "01001110100110111" => rgb <= "000000";
					when "01001110100111000" => rgb <= "000000";
					when "01001110100111001" => rgb <= "000000";
					when "01001110100111010" => rgb <= "000000";
					when "01001110100111011" => rgb <= "000000";
					when "01001110100111100" => rgb <= "000000";
					when "01001110100111101" => rgb <= "000000";
					when "01001110100111110" => rgb <= "000000";
					when "01001110100111111" => rgb <= "000000";
					when "01001111000000000" => rgb <= "000000";
					when "01001111000000001" => rgb <= "000000";
					when "01001111000000010" => rgb <= "000000";
					when "01001111000000011" => rgb <= "000000";
					when "01001111000000100" => rgb <= "000000";
					when "01001111000000101" => rgb <= "000000";
					when "01001111000000110" => rgb <= "000000";
					when "01001111000000111" => rgb <= "000000";
					when "01001111000001000" => rgb <= "000000";
					when "01001111000001001" => rgb <= "000000";
					when "01001111000001010" => rgb <= "000000";
					when "01001111000001011" => rgb <= "000000";
					when "01001111000001100" => rgb <= "000000";
					when "01001111000001101" => rgb <= "000000";
					when "01001111000001110" => rgb <= "000000";
					when "01001111000001111" => rgb <= "000000";
					when "01001111000010000" => rgb <= "000000";
					when "01001111000010001" => rgb <= "000000";
					when "01001111000010010" => rgb <= "000000";
					when "01001111000010011" => rgb <= "000000";
					when "01001111000010100" => rgb <= "000000";
					when "01001111000010101" => rgb <= "000000";
					when "01001111000010110" => rgb <= "000000";
					when "01001111000010111" => rgb <= "000000";
					when "01001111000011000" => rgb <= "000000";
					when "01001111000011001" => rgb <= "000000";
					when "01001111000011010" => rgb <= "000000";
					when "01001111000011011" => rgb <= "000000";
					when "01001111000011100" => rgb <= "000000";
					when "01001111000011101" => rgb <= "000000";
					when "01001111000011110" => rgb <= "000000";
					when "01001111000011111" => rgb <= "000000";
					when "01001111000100000" => rgb <= "000000";
					when "01001111000100001" => rgb <= "000000";
					when "01001111000100010" => rgb <= "000000";
					when "01001111000100011" => rgb <= "000000";
					when "01001111000100100" => rgb <= "000000";
					when "01001111000100101" => rgb <= "000000";
					when "01001111000100110" => rgb <= "000000";
					when "01001111000100111" => rgb <= "000000";
					when "01001111000101000" => rgb <= "000000";
					when "01001111000101001" => rgb <= "000000";
					when "01001111000101010" => rgb <= "000000";
					when "01001111000101011" => rgb <= "000000";
					when "01001111000101100" => rgb <= "000000";
					when "01001111000101101" => rgb <= "000000";
					when "01001111000101110" => rgb <= "000000";
					when "01001111000101111" => rgb <= "000000";
					when "01001111000110000" => rgb <= "000000";
					when "01001111000110001" => rgb <= "000000";
					when "01001111000110010" => rgb <= "000000";
					when "01001111000110011" => rgb <= "000000";
					when "01001111000110100" => rgb <= "000000";
					when "01001111000110101" => rgb <= "000000";
					when "01001111000110110" => rgb <= "000000";
					when "01001111000110111" => rgb <= "000000";
					when "01001111000111000" => rgb <= "000000";
					when "01001111000111001" => rgb <= "000000";
					when "01001111000111010" => rgb <= "000000";
					when "01001111000111011" => rgb <= "000000";
					when "01001111000111100" => rgb <= "000000";
					when "01001111000111101" => rgb <= "000000";
					when "01001111000111110" => rgb <= "000000";
					when "01001111000111111" => rgb <= "000000";
					when "01001111001000000" => rgb <= "000000";
					when "01001111001000001" => rgb <= "000000";
					when "01001111001000010" => rgb <= "000000";
					when "01001111001000011" => rgb <= "000000";
					when "01001111001000100" => rgb <= "000000";
					when "01001111001000101" => rgb <= "000000";
					when "01001111001000110" => rgb <= "000000";
					when "01001111001000111" => rgb <= "000000";
					when "01001111001001000" => rgb <= "000000";
					when "01001111001001001" => rgb <= "000000";
					when "01001111001001010" => rgb <= "000000";
					when "01001111001001011" => rgb <= "000000";
					when "01001111001001100" => rgb <= "000000";
					when "01001111001001101" => rgb <= "000000";
					when "01001111001001110" => rgb <= "000000";
					when "01001111001001111" => rgb <= "000000";
					when "01001111001010000" => rgb <= "000000";
					when "01001111001010001" => rgb <= "000000";
					when "01001111001010010" => rgb <= "000000";
					when "01001111001010011" => rgb <= "000000";
					when "01001111001010100" => rgb <= "000000";
					when "01001111001010101" => rgb <= "000000";
					when "01001111001010110" => rgb <= "000000";
					when "01001111001010111" => rgb <= "000000";
					when "01001111001011000" => rgb <= "000000";
					when "01001111001011001" => rgb <= "000000";
					when "01001111001011010" => rgb <= "000000";
					when "01001111001011011" => rgb <= "000000";
					when "01001111001011100" => rgb <= "000000";
					when "01001111001011101" => rgb <= "000000";
					when "01001111001011110" => rgb <= "000000";
					when "01001111001011111" => rgb <= "000000";
					when "01001111001100000" => rgb <= "000000";
					when "01001111001100001" => rgb <= "000000";
					when "01001111001100010" => rgb <= "000000";
					when "01001111001100011" => rgb <= "000000";
					when "01001111001100100" => rgb <= "000000";
					when "01001111001100101" => rgb <= "000000";
					when "01001111001100110" => rgb <= "000000";
					when "01001111001100111" => rgb <= "000000";
					when "01001111001101000" => rgb <= "000000";
					when "01001111001101001" => rgb <= "000000";
					when "01001111001101010" => rgb <= "000000";
					when "01001111001101011" => rgb <= "000000";
					when "01001111001101100" => rgb <= "000000";
					when "01001111001101101" => rgb <= "000000";
					when "01001111001101110" => rgb <= "000000";
					when "01001111001101111" => rgb <= "000000";
					when "01001111001110000" => rgb <= "000000";
					when "01001111001110001" => rgb <= "000000";
					when "01001111001110010" => rgb <= "000000";
					when "01001111001110011" => rgb <= "000000";
					when "01001111001110100" => rgb <= "000000";
					when "01001111001110101" => rgb <= "000000";
					when "01001111001110110" => rgb <= "000000";
					when "01001111001110111" => rgb <= "000000";
					when "01001111001111000" => rgb <= "000000";
					when "01001111001111001" => rgb <= "000000";
					when "01001111001111010" => rgb <= "000000";
					when "01001111001111011" => rgb <= "000000";
					when "01001111001111100" => rgb <= "000000";
					when "01001111001111101" => rgb <= "000000";
					when "01001111001111110" => rgb <= "000000";
					when "01001111001111111" => rgb <= "000000";
					when "01001111010000000" => rgb <= "000000";
					when "01001111010000001" => rgb <= "000000";
					when "01001111010000010" => rgb <= "000000";
					when "01001111010000011" => rgb <= "000000";
					when "01001111010000100" => rgb <= "000000";
					when "01001111010000101" => rgb <= "000000";
					when "01001111010000110" => rgb <= "000000";
					when "01001111010000111" => rgb <= "000000";
					when "01001111010001000" => rgb <= "100100";
					when "01001111010001001" => rgb <= "101000";
					when "01001111010001010" => rgb <= "101000";
					when "01001111010001011" => rgb <= "101000";
					when "01001111010001100" => rgb <= "101000";
					when "01001111010001101" => rgb <= "101000";
					when "01001111010001110" => rgb <= "101000";
					when "01001111010001111" => rgb <= "101000";
					when "01001111010010000" => rgb <= "101000";
					when "01001111010010001" => rgb <= "101000";
					when "01001111010010010" => rgb <= "101000";
					when "01001111010010011" => rgb <= "101000";
					when "01001111010010100" => rgb <= "101000";
					when "01001111010010101" => rgb <= "101000";
					when "01001111010010110" => rgb <= "101000";
					when "01001111010010111" => rgb <= "101000";
					when "01001111010011000" => rgb <= "101000";
					when "01001111010011001" => rgb <= "101000";
					when "01001111010011010" => rgb <= "101000";
					when "01001111010011011" => rgb <= "101000";
					when "01001111010011100" => rgb <= "101000";
					when "01001111010011101" => rgb <= "101000";
					when "01001111010011110" => rgb <= "101000";
					when "01001111010011111" => rgb <= "101000";
					when "01001111010100000" => rgb <= "101000";
					when "01001111010100001" => rgb <= "101000";
					when "01001111010100010" => rgb <= "101000";
					when "01001111010100011" => rgb <= "101000";
					when "01001111010100100" => rgb <= "101000";
					when "01001111010100101" => rgb <= "101000";
					when "01001111010100110" => rgb <= "101000";
					when "01001111010100111" => rgb <= "101000";
					when "01001111010101000" => rgb <= "101000";
					when "01001111010101001" => rgb <= "101000";
					when "01001111010101010" => rgb <= "101000";
					when "01001111010101011" => rgb <= "101000";
					when "01001111010101100" => rgb <= "101000";
					when "01001111010101101" => rgb <= "101000";
					when "01001111010101110" => rgb <= "101000";
					when "01001111010101111" => rgb <= "101000";
					when "01001111010110000" => rgb <= "101000";
					when "01001111010110001" => rgb <= "101000";
					when "01001111010110010" => rgb <= "101000";
					when "01001111010110011" => rgb <= "101000";
					when "01001111010110100" => rgb <= "101000";
					when "01001111010110101" => rgb <= "010100";
					when "01001111010110110" => rgb <= "000000";
					when "01001111010110111" => rgb <= "000000";
					when "01001111010111000" => rgb <= "000000";
					when "01001111010111001" => rgb <= "000000";
					when "01001111010111010" => rgb <= "000000";
					when "01001111010111011" => rgb <= "000000";
					when "01001111010111100" => rgb <= "000000";
					when "01001111010111101" => rgb <= "000000";
					when "01001111010111110" => rgb <= "000000";
					when "01001111010111111" => rgb <= "000000";
					when "01001111011000000" => rgb <= "000000";
					when "01001111011000001" => rgb <= "000000";
					when "01001111011000010" => rgb <= "000000";
					when "01001111011000011" => rgb <= "000000";
					when "01001111011000100" => rgb <= "000000";
					when "01001111011000101" => rgb <= "000000";
					when "01001111011000110" => rgb <= "000000";
					when "01001111011000111" => rgb <= "000000";
					when "01001111011001000" => rgb <= "000000";
					when "01001111011001001" => rgb <= "000000";
					when "01001111011001010" => rgb <= "000000";
					when "01001111011001011" => rgb <= "000000";
					when "01001111011001100" => rgb <= "000000";
					when "01001111011001101" => rgb <= "000000";
					when "01001111011001110" => rgb <= "000000";
					when "01001111011001111" => rgb <= "000000";
					when "01001111011010000" => rgb <= "000000";
					when "01001111011010001" => rgb <= "000000";
					when "01001111011010010" => rgb <= "000000";
					when "01001111011010011" => rgb <= "000000";
					when "01001111011010100" => rgb <= "000000";
					when "01001111011010101" => rgb <= "000000";
					when "01001111011010110" => rgb <= "000000";
					when "01001111011010111" => rgb <= "000000";
					when "01001111011011000" => rgb <= "000000";
					when "01001111011011001" => rgb <= "000000";
					when "01001111011011010" => rgb <= "000000";
					when "01001111011011011" => rgb <= "000000";
					when "01001111011011100" => rgb <= "000000";
					when "01001111011011101" => rgb <= "000000";
					when "01001111011011110" => rgb <= "000000";
					when "01001111011011111" => rgb <= "000000";
					when "01001111011100000" => rgb <= "000000";
					when "01001111011100001" => rgb <= "000000";
					when "01001111011100010" => rgb <= "000000";
					when "01001111011100011" => rgb <= "000000";
					when "01001111011100100" => rgb <= "000000";
					when "01001111011100101" => rgb <= "000000";
					when "01001111011100110" => rgb <= "000000";
					when "01001111011100111" => rgb <= "000000";
					when "01001111011101000" => rgb <= "000000";
					when "01001111011101001" => rgb <= "000000";
					when "01001111011101010" => rgb <= "000000";
					when "01001111011101011" => rgb <= "000000";
					when "01001111011101100" => rgb <= "000000";
					when "01001111011101101" => rgb <= "000000";
					when "01001111011101110" => rgb <= "000000";
					when "01001111011101111" => rgb <= "000000";
					when "01001111011110000" => rgb <= "000000";
					when "01001111011110001" => rgb <= "000000";
					when "01001111011110010" => rgb <= "000000";
					when "01001111011110011" => rgb <= "000000";
					when "01001111011110100" => rgb <= "000000";
					when "01001111011110101" => rgb <= "000000";
					when "01001111011110110" => rgb <= "000000";
					when "01001111011110111" => rgb <= "000000";
					when "01001111011111000" => rgb <= "000000";
					when "01001111011111001" => rgb <= "000000";
					when "01001111011111010" => rgb <= "000000";
					when "01001111011111011" => rgb <= "000000";
					when "01001111011111100" => rgb <= "000000";
					when "01001111011111101" => rgb <= "000000";
					when "01001111011111110" => rgb <= "000000";
					when "01001111011111111" => rgb <= "000000";
					when "01001111100000000" => rgb <= "000000";
					when "01001111100000001" => rgb <= "000000";
					when "01001111100000010" => rgb <= "000000";
					when "01001111100000011" => rgb <= "000000";
					when "01001111100000100" => rgb <= "000000";
					when "01001111100000101" => rgb <= "000000";
					when "01001111100000110" => rgb <= "000000";
					when "01001111100000111" => rgb <= "000000";
					when "01001111100001000" => rgb <= "000000";
					when "01001111100001001" => rgb <= "000000";
					when "01001111100001010" => rgb <= "000000";
					when "01001111100001011" => rgb <= "000000";
					when "01001111100001100" => rgb <= "000000";
					when "01001111100001101" => rgb <= "000000";
					when "01001111100001110" => rgb <= "000000";
					when "01001111100001111" => rgb <= "000000";
					when "01001111100010000" => rgb <= "000000";
					when "01001111100010001" => rgb <= "000000";
					when "01001111100010010" => rgb <= "000000";
					when "01001111100010011" => rgb <= "000000";
					when "01001111100010100" => rgb <= "000000";
					when "01001111100010101" => rgb <= "000000";
					when "01001111100010110" => rgb <= "000000";
					when "01001111100010111" => rgb <= "000000";
					when "01001111100011000" => rgb <= "000000";
					when "01001111100011001" => rgb <= "000000";
					when "01001111100011010" => rgb <= "000000";
					when "01001111100011011" => rgb <= "000000";
					when "01001111100011100" => rgb <= "000000";
					when "01001111100011101" => rgb <= "000000";
					when "01001111100011110" => rgb <= "000000";
					when "01001111100011111" => rgb <= "000000";
					when "01001111100100000" => rgb <= "000000";
					when "01001111100100001" => rgb <= "000000";
					when "01001111100100010" => rgb <= "000000";
					when "01001111100100011" => rgb <= "000000";
					when "01001111100100100" => rgb <= "000000";
					when "01001111100100101" => rgb <= "000000";
					when "01001111100100110" => rgb <= "000000";
					when "01001111100100111" => rgb <= "000000";
					when "01001111100101000" => rgb <= "000000";
					when "01001111100101001" => rgb <= "000000";
					when "01001111100101010" => rgb <= "000000";
					when "01001111100101011" => rgb <= "000000";
					when "01001111100101100" => rgb <= "000000";
					when "01001111100101101" => rgb <= "000000";
					when "01001111100101110" => rgb <= "000000";
					when "01001111100101111" => rgb <= "000000";
					when "01001111100110000" => rgb <= "000000";
					when "01001111100110001" => rgb <= "000000";
					when "01001111100110010" => rgb <= "000000";
					when "01001111100110011" => rgb <= "000000";
					when "01001111100110100" => rgb <= "000000";
					when "01001111100110101" => rgb <= "000000";
					when "01001111100110110" => rgb <= "000000";
					when "01001111100110111" => rgb <= "000000";
					when "01001111100111000" => rgb <= "000000";
					when "01001111100111001" => rgb <= "000000";
					when "01001111100111010" => rgb <= "000000";
					when "01001111100111011" => rgb <= "000000";
					when "01001111100111100" => rgb <= "000000";
					when "01001111100111101" => rgb <= "000000";
					when "01001111100111110" => rgb <= "000000";
					when "01001111100111111" => rgb <= "000000";
					when "01010000000000000" => rgb <= "000000";
					when "01010000000000001" => rgb <= "000000";
					when "01010000000000010" => rgb <= "000000";
					when "01010000000000011" => rgb <= "000000";
					when "01010000000000100" => rgb <= "000000";
					when "01010000000000101" => rgb <= "000000";
					when "01010000000000110" => rgb <= "000000";
					when "01010000000000111" => rgb <= "000000";
					when "01010000000001000" => rgb <= "000000";
					when "01010000000001001" => rgb <= "000000";
					when "01010000000001010" => rgb <= "000000";
					when "01010000000001011" => rgb <= "000000";
					when "01010000000001100" => rgb <= "000000";
					when "01010000000001101" => rgb <= "000000";
					when "01010000000001110" => rgb <= "000000";
					when "01010000000001111" => rgb <= "000000";
					when "01010000000010000" => rgb <= "000000";
					when "01010000000010001" => rgb <= "000000";
					when "01010000000010010" => rgb <= "000000";
					when "01010000000010011" => rgb <= "000000";
					when "01010000000010100" => rgb <= "000000";
					when "01010000000010101" => rgb <= "000000";
					when "01010000000010110" => rgb <= "000000";
					when "01010000000010111" => rgb <= "000000";
					when "01010000000011000" => rgb <= "000000";
					when "01010000000011001" => rgb <= "000000";
					when "01010000000011010" => rgb <= "000000";
					when "01010000000011011" => rgb <= "000000";
					when "01010000000011100" => rgb <= "000000";
					when "01010000000011101" => rgb <= "000000";
					when "01010000000011110" => rgb <= "000000";
					when "01010000000011111" => rgb <= "000000";
					when "01010000000100000" => rgb <= "000000";
					when "01010000000100001" => rgb <= "000000";
					when "01010000000100010" => rgb <= "000000";
					when "01010000000100011" => rgb <= "000000";
					when "01010000000100100" => rgb <= "000000";
					when "01010000000100101" => rgb <= "000000";
					when "01010000000100110" => rgb <= "000000";
					when "01010000000100111" => rgb <= "000000";
					when "01010000000101000" => rgb <= "000000";
					when "01010000000101001" => rgb <= "000000";
					when "01010000000101010" => rgb <= "000000";
					when "01010000000101011" => rgb <= "000000";
					when "01010000000101100" => rgb <= "000000";
					when "01010000000101101" => rgb <= "000000";
					when "01010000000101110" => rgb <= "000000";
					when "01010000000101111" => rgb <= "000000";
					when "01010000000110000" => rgb <= "000000";
					when "01010000000110001" => rgb <= "000000";
					when "01010000000110010" => rgb <= "000000";
					when "01010000000110011" => rgb <= "000000";
					when "01010000000110100" => rgb <= "000000";
					when "01010000000110101" => rgb <= "000000";
					when "01010000000110110" => rgb <= "000000";
					when "01010000000110111" => rgb <= "000000";
					when "01010000000111000" => rgb <= "000000";
					when "01010000000111001" => rgb <= "000000";
					when "01010000000111010" => rgb <= "000000";
					when "01010000000111011" => rgb <= "000000";
					when "01010000000111100" => rgb <= "000000";
					when "01010000000111101" => rgb <= "000000";
					when "01010000000111110" => rgb <= "000000";
					when "01010000000111111" => rgb <= "000000";
					when "01010000001000000" => rgb <= "000000";
					when "01010000001000001" => rgb <= "000000";
					when "01010000001000010" => rgb <= "000000";
					when "01010000001000011" => rgb <= "000000";
					when "01010000001000100" => rgb <= "000000";
					when "01010000001000101" => rgb <= "000000";
					when "01010000001000110" => rgb <= "000000";
					when "01010000001000111" => rgb <= "000000";
					when "01010000001001000" => rgb <= "000000";
					when "01010000001001001" => rgb <= "000000";
					when "01010000001001010" => rgb <= "000000";
					when "01010000001001011" => rgb <= "000000";
					when "01010000001001100" => rgb <= "000000";
					when "01010000001001101" => rgb <= "000000";
					when "01010000001001110" => rgb <= "000000";
					when "01010000001001111" => rgb <= "000000";
					when "01010000001010000" => rgb <= "000000";
					when "01010000001010001" => rgb <= "000000";
					when "01010000001010010" => rgb <= "000000";
					when "01010000001010011" => rgb <= "000000";
					when "01010000001010100" => rgb <= "000000";
					when "01010000001010101" => rgb <= "000000";
					when "01010000001010110" => rgb <= "000000";
					when "01010000001010111" => rgb <= "000000";
					when "01010000001011000" => rgb <= "000000";
					when "01010000001011001" => rgb <= "000000";
					when "01010000001011010" => rgb <= "000000";
					when "01010000001011011" => rgb <= "000000";
					when "01010000001011100" => rgb <= "000000";
					when "01010000001011101" => rgb <= "000000";
					when "01010000001011110" => rgb <= "000000";
					when "01010000001011111" => rgb <= "000000";
					when "01010000001100000" => rgb <= "000000";
					when "01010000001100001" => rgb <= "000000";
					when "01010000001100010" => rgb <= "000000";
					when "01010000001100011" => rgb <= "000000";
					when "01010000001100100" => rgb <= "000000";
					when "01010000001100101" => rgb <= "000000";
					when "01010000001100110" => rgb <= "000000";
					when "01010000001100111" => rgb <= "000000";
					when "01010000001101000" => rgb <= "000000";
					when "01010000001101001" => rgb <= "000000";
					when "01010000001101010" => rgb <= "000000";
					when "01010000001101011" => rgb <= "000000";
					when "01010000001101100" => rgb <= "000000";
					when "01010000001101101" => rgb <= "000000";
					when "01010000001101110" => rgb <= "000000";
					when "01010000001101111" => rgb <= "000000";
					when "01010000001110000" => rgb <= "000000";
					when "01010000001110001" => rgb <= "000000";
					when "01010000001110010" => rgb <= "000000";
					when "01010000001110011" => rgb <= "000000";
					when "01010000001110100" => rgb <= "000000";
					when "01010000001110101" => rgb <= "000000";
					when "01010000001110110" => rgb <= "000000";
					when "01010000001110111" => rgb <= "000000";
					when "01010000001111000" => rgb <= "000000";
					when "01010000001111001" => rgb <= "000000";
					when "01010000001111010" => rgb <= "000000";
					when "01010000001111011" => rgb <= "000000";
					when "01010000001111100" => rgb <= "000000";
					when "01010000001111101" => rgb <= "000000";
					when "01010000001111110" => rgb <= "000000";
					when "01010000001111111" => rgb <= "000000";
					when "01010000010000000" => rgb <= "000000";
					when "01010000010000001" => rgb <= "000000";
					when "01010000010000010" => rgb <= "000000";
					when "01010000010000011" => rgb <= "000000";
					when "01010000010000100" => rgb <= "000000";
					when "01010000010000101" => rgb <= "000000";
					when "01010000010000110" => rgb <= "000000";
					when "01010000010000111" => rgb <= "000000";
					when "01010000010001000" => rgb <= "100100";
					when "01010000010001001" => rgb <= "101000";
					when "01010000010001010" => rgb <= "101000";
					when "01010000010001011" => rgb <= "101000";
					when "01010000010001100" => rgb <= "101000";
					when "01010000010001101" => rgb <= "101000";
					when "01010000010001110" => rgb <= "101000";
					when "01010000010001111" => rgb <= "101000";
					when "01010000010010000" => rgb <= "101000";
					when "01010000010010001" => rgb <= "101001";
					when "01010000010010010" => rgb <= "101000";
					when "01010000010010011" => rgb <= "101000";
					when "01010000010010100" => rgb <= "101000";
					when "01010000010010101" => rgb <= "101000";
					when "01010000010010110" => rgb <= "101000";
					when "01010000010010111" => rgb <= "101000";
					when "01010000010011000" => rgb <= "101000";
					when "01010000010011001" => rgb <= "101000";
					when "01010000010011010" => rgb <= "101000";
					when "01010000010011011" => rgb <= "101000";
					when "01010000010011100" => rgb <= "101000";
					when "01010000010011101" => rgb <= "101000";
					when "01010000010011110" => rgb <= "101000";
					when "01010000010011111" => rgb <= "101000";
					when "01010000010100000" => rgb <= "101000";
					when "01010000010100001" => rgb <= "101000";
					when "01010000010100010" => rgb <= "101000";
					when "01010000010100011" => rgb <= "101000";
					when "01010000010100100" => rgb <= "101000";
					when "01010000010100101" => rgb <= "101000";
					when "01010000010100110" => rgb <= "101000";
					when "01010000010100111" => rgb <= "101000";
					when "01010000010101000" => rgb <= "101000";
					when "01010000010101001" => rgb <= "101001";
					when "01010000010101010" => rgb <= "101000";
					when "01010000010101011" => rgb <= "101000";
					when "01010000010101100" => rgb <= "101000";
					when "01010000010101101" => rgb <= "101000";
					when "01010000010101110" => rgb <= "101000";
					when "01010000010101111" => rgb <= "101000";
					when "01010000010110000" => rgb <= "101000";
					when "01010000010110001" => rgb <= "101000";
					when "01010000010110010" => rgb <= "101000";
					when "01010000010110011" => rgb <= "101000";
					when "01010000010110100" => rgb <= "101000";
					when "01010000010110101" => rgb <= "010100";
					when "01010000010110110" => rgb <= "000000";
					when "01010000010110111" => rgb <= "000000";
					when "01010000010111000" => rgb <= "000000";
					when "01010000010111001" => rgb <= "000000";
					when "01010000010111010" => rgb <= "000000";
					when "01010000010111011" => rgb <= "000000";
					when "01010000010111100" => rgb <= "000000";
					when "01010000010111101" => rgb <= "000000";
					when "01010000010111110" => rgb <= "000000";
					when "01010000010111111" => rgb <= "000000";
					when "01010000011000000" => rgb <= "000000";
					when "01010000011000001" => rgb <= "000000";
					when "01010000011000010" => rgb <= "000000";
					when "01010000011000011" => rgb <= "000000";
					when "01010000011000100" => rgb <= "000000";
					when "01010000011000101" => rgb <= "000000";
					when "01010000011000110" => rgb <= "000000";
					when "01010000011000111" => rgb <= "000000";
					when "01010000011001000" => rgb <= "000000";
					when "01010000011001001" => rgb <= "000000";
					when "01010000011001010" => rgb <= "000000";
					when "01010000011001011" => rgb <= "000000";
					when "01010000011001100" => rgb <= "000000";
					when "01010000011001101" => rgb <= "000000";
					when "01010000011001110" => rgb <= "000000";
					when "01010000011001111" => rgb <= "000000";
					when "01010000011010000" => rgb <= "000000";
					when "01010000011010001" => rgb <= "000000";
					when "01010000011010010" => rgb <= "000000";
					when "01010000011010011" => rgb <= "000000";
					when "01010000011010100" => rgb <= "000000";
					when "01010000011010101" => rgb <= "000000";
					when "01010000011010110" => rgb <= "000000";
					when "01010000011010111" => rgb <= "000000";
					when "01010000011011000" => rgb <= "000000";
					when "01010000011011001" => rgb <= "000000";
					when "01010000011011010" => rgb <= "000000";
					when "01010000011011011" => rgb <= "000000";
					when "01010000011011100" => rgb <= "000000";
					when "01010000011011101" => rgb <= "000000";
					when "01010000011011110" => rgb <= "000000";
					when "01010000011011111" => rgb <= "000000";
					when "01010000011100000" => rgb <= "000000";
					when "01010000011100001" => rgb <= "000000";
					when "01010000011100010" => rgb <= "000000";
					when "01010000011100011" => rgb <= "000000";
					when "01010000011100100" => rgb <= "000000";
					when "01010000011100101" => rgb <= "000000";
					when "01010000011100110" => rgb <= "000000";
					when "01010000011100111" => rgb <= "000000";
					when "01010000011101000" => rgb <= "000000";
					when "01010000011101001" => rgb <= "000000";
					when "01010000011101010" => rgb <= "000000";
					when "01010000011101011" => rgb <= "000000";
					when "01010000011101100" => rgb <= "000000";
					when "01010000011101101" => rgb <= "000000";
					when "01010000011101110" => rgb <= "000000";
					when "01010000011101111" => rgb <= "000000";
					when "01010000011110000" => rgb <= "000000";
					when "01010000011110001" => rgb <= "000000";
					when "01010000011110010" => rgb <= "000000";
					when "01010000011110011" => rgb <= "000000";
					when "01010000011110100" => rgb <= "000000";
					when "01010000011110101" => rgb <= "000000";
					when "01010000011110110" => rgb <= "000000";
					when "01010000011110111" => rgb <= "000000";
					when "01010000011111000" => rgb <= "000000";
					when "01010000011111001" => rgb <= "000000";
					when "01010000011111010" => rgb <= "000000";
					when "01010000011111011" => rgb <= "000000";
					when "01010000011111100" => rgb <= "000000";
					when "01010000011111101" => rgb <= "000000";
					when "01010000011111110" => rgb <= "000000";
					when "01010000011111111" => rgb <= "000000";
					when "01010000100000000" => rgb <= "000000";
					when "01010000100000001" => rgb <= "000000";
					when "01010000100000010" => rgb <= "000000";
					when "01010000100000011" => rgb <= "000000";
					when "01010000100000100" => rgb <= "000000";
					when "01010000100000101" => rgb <= "000000";
					when "01010000100000110" => rgb <= "000000";
					when "01010000100000111" => rgb <= "000000";
					when "01010000100001000" => rgb <= "000000";
					when "01010000100001001" => rgb <= "000000";
					when "01010000100001010" => rgb <= "000000";
					when "01010000100001011" => rgb <= "000000";
					when "01010000100001100" => rgb <= "000000";
					when "01010000100001101" => rgb <= "000000";
					when "01010000100001110" => rgb <= "000000";
					when "01010000100001111" => rgb <= "000000";
					when "01010000100010000" => rgb <= "000000";
					when "01010000100010001" => rgb <= "000000";
					when "01010000100010010" => rgb <= "000000";
					when "01010000100010011" => rgb <= "000000";
					when "01010000100010100" => rgb <= "000000";
					when "01010000100010101" => rgb <= "000000";
					when "01010000100010110" => rgb <= "000000";
					when "01010000100010111" => rgb <= "000000";
					when "01010000100011000" => rgb <= "000000";
					when "01010000100011001" => rgb <= "000000";
					when "01010000100011010" => rgb <= "000000";
					when "01010000100011011" => rgb <= "000000";
					when "01010000100011100" => rgb <= "000000";
					when "01010000100011101" => rgb <= "000000";
					when "01010000100011110" => rgb <= "000000";
					when "01010000100011111" => rgb <= "000000";
					when "01010000100100000" => rgb <= "000000";
					when "01010000100100001" => rgb <= "000000";
					when "01010000100100010" => rgb <= "000000";
					when "01010000100100011" => rgb <= "000000";
					when "01010000100100100" => rgb <= "000000";
					when "01010000100100101" => rgb <= "000000";
					when "01010000100100110" => rgb <= "000000";
					when "01010000100100111" => rgb <= "000000";
					when "01010000100101000" => rgb <= "000000";
					when "01010000100101001" => rgb <= "000000";
					when "01010000100101010" => rgb <= "000000";
					when "01010000100101011" => rgb <= "000000";
					when "01010000100101100" => rgb <= "000000";
					when "01010000100101101" => rgb <= "000000";
					when "01010000100101110" => rgb <= "000000";
					when "01010000100101111" => rgb <= "000000";
					when "01010000100110000" => rgb <= "000000";
					when "01010000100110001" => rgb <= "000000";
					when "01010000100110010" => rgb <= "000000";
					when "01010000100110011" => rgb <= "000000";
					when "01010000100110100" => rgb <= "000000";
					when "01010000100110101" => rgb <= "000000";
					when "01010000100110110" => rgb <= "000000";
					when "01010000100110111" => rgb <= "000000";
					when "01010000100111000" => rgb <= "000000";
					when "01010000100111001" => rgb <= "000000";
					when "01010000100111010" => rgb <= "000000";
					when "01010000100111011" => rgb <= "000000";
					when "01010000100111100" => rgb <= "000000";
					when "01010000100111101" => rgb <= "000000";
					when "01010000100111110" => rgb <= "000000";
					when "01010000100111111" => rgb <= "000000";
					when "01010001000000000" => rgb <= "000000";
					when "01010001000000001" => rgb <= "000000";
					when "01010001000000010" => rgb <= "000000";
					when "01010001000000011" => rgb <= "000000";
					when "01010001000000100" => rgb <= "000000";
					when "01010001000000101" => rgb <= "000000";
					when "01010001000000110" => rgb <= "000000";
					when "01010001000000111" => rgb <= "000000";
					when "01010001000001000" => rgb <= "000000";
					when "01010001000001001" => rgb <= "000000";
					when "01010001000001010" => rgb <= "000000";
					when "01010001000001011" => rgb <= "000000";
					when "01010001000001100" => rgb <= "000000";
					when "01010001000001101" => rgb <= "000000";
					when "01010001000001110" => rgb <= "000000";
					when "01010001000001111" => rgb <= "000000";
					when "01010001000010000" => rgb <= "000000";
					when "01010001000010001" => rgb <= "000000";
					when "01010001000010010" => rgb <= "000000";
					when "01010001000010011" => rgb <= "000000";
					when "01010001000010100" => rgb <= "000000";
					when "01010001000010101" => rgb <= "000000";
					when "01010001000010110" => rgb <= "000000";
					when "01010001000010111" => rgb <= "000000";
					when "01010001000011000" => rgb <= "000000";
					when "01010001000011001" => rgb <= "000000";
					when "01010001000011010" => rgb <= "000000";
					when "01010001000011011" => rgb <= "000000";
					when "01010001000011100" => rgb <= "000000";
					when "01010001000011101" => rgb <= "000000";
					when "01010001000011110" => rgb <= "000000";
					when "01010001000011111" => rgb <= "000000";
					when "01010001000100000" => rgb <= "000000";
					when "01010001000100001" => rgb <= "000000";
					when "01010001000100010" => rgb <= "000000";
					when "01010001000100011" => rgb <= "000000";
					when "01010001000100100" => rgb <= "000000";
					when "01010001000100101" => rgb <= "000000";
					when "01010001000100110" => rgb <= "000000";
					when "01010001000100111" => rgb <= "000000";
					when "01010001000101000" => rgb <= "000000";
					when "01010001000101001" => rgb <= "000000";
					when "01010001000101010" => rgb <= "000000";
					when "01010001000101011" => rgb <= "000000";
					when "01010001000101100" => rgb <= "000000";
					when "01010001000101101" => rgb <= "000000";
					when "01010001000101110" => rgb <= "000000";
					when "01010001000101111" => rgb <= "000000";
					when "01010001000110000" => rgb <= "000000";
					when "01010001000110001" => rgb <= "000000";
					when "01010001000110010" => rgb <= "000000";
					when "01010001000110011" => rgb <= "000000";
					when "01010001000110100" => rgb <= "000000";
					when "01010001000110101" => rgb <= "000000";
					when "01010001000110110" => rgb <= "000000";
					when "01010001000110111" => rgb <= "000000";
					when "01010001000111000" => rgb <= "000000";
					when "01010001000111001" => rgb <= "000000";
					when "01010001000111010" => rgb <= "000000";
					when "01010001000111011" => rgb <= "000000";
					when "01010001000111100" => rgb <= "000000";
					when "01010001000111101" => rgb <= "000000";
					when "01010001000111110" => rgb <= "000000";
					when "01010001000111111" => rgb <= "000000";
					when "01010001001000000" => rgb <= "000000";
					when "01010001001000001" => rgb <= "000000";
					when "01010001001000010" => rgb <= "000000";
					when "01010001001000011" => rgb <= "000000";
					when "01010001001000100" => rgb <= "000000";
					when "01010001001000101" => rgb <= "000000";
					when "01010001001000110" => rgb <= "000000";
					when "01010001001000111" => rgb <= "000000";
					when "01010001001001000" => rgb <= "000000";
					when "01010001001001001" => rgb <= "000000";
					when "01010001001001010" => rgb <= "000000";
					when "01010001001001011" => rgb <= "000000";
					when "01010001001001100" => rgb <= "000000";
					when "01010001001001101" => rgb <= "000000";
					when "01010001001001110" => rgb <= "000000";
					when "01010001001001111" => rgb <= "000000";
					when "01010001001010000" => rgb <= "000000";
					when "01010001001010001" => rgb <= "000000";
					when "01010001001010010" => rgb <= "000000";
					when "01010001001010011" => rgb <= "000000";
					when "01010001001010100" => rgb <= "000000";
					when "01010001001010101" => rgb <= "000000";
					when "01010001001010110" => rgb <= "000000";
					when "01010001001010111" => rgb <= "000000";
					when "01010001001011000" => rgb <= "000000";
					when "01010001001011001" => rgb <= "000000";
					when "01010001001011010" => rgb <= "000000";
					when "01010001001011011" => rgb <= "000000";
					when "01010001001011100" => rgb <= "000000";
					when "01010001001011101" => rgb <= "000000";
					when "01010001001011110" => rgb <= "000000";
					when "01010001001011111" => rgb <= "000000";
					when "01010001001100000" => rgb <= "000000";
					when "01010001001100001" => rgb <= "000000";
					when "01010001001100010" => rgb <= "000000";
					when "01010001001100011" => rgb <= "000000";
					when "01010001001100100" => rgb <= "000000";
					when "01010001001100101" => rgb <= "000000";
					when "01010001001100110" => rgb <= "000000";
					when "01010001001100111" => rgb <= "000000";
					when "01010001001101000" => rgb <= "000000";
					when "01010001001101001" => rgb <= "000000";
					when "01010001001101010" => rgb <= "000000";
					when "01010001001101011" => rgb <= "000000";
					when "01010001001101100" => rgb <= "000000";
					when "01010001001101101" => rgb <= "000000";
					when "01010001001101110" => rgb <= "000000";
					when "01010001001101111" => rgb <= "000000";
					when "01010001001110000" => rgb <= "000000";
					when "01010001001110001" => rgb <= "000000";
					when "01010001001110010" => rgb <= "000000";
					when "01010001001110011" => rgb <= "000000";
					when "01010001001110100" => rgb <= "000000";
					when "01010001001110101" => rgb <= "000000";
					when "01010001001110110" => rgb <= "000000";
					when "01010001001110111" => rgb <= "000000";
					when "01010001001111000" => rgb <= "000000";
					when "01010001001111001" => rgb <= "000000";
					when "01010001001111010" => rgb <= "000000";
					when "01010001001111011" => rgb <= "000000";
					when "01010001001111100" => rgb <= "000000";
					when "01010001001111101" => rgb <= "000000";
					when "01010001001111110" => rgb <= "000000";
					when "01010001001111111" => rgb <= "000000";
					when "01010001010000000" => rgb <= "000000";
					when "01010001010000001" => rgb <= "000000";
					when "01010001010000010" => rgb <= "000000";
					when "01010001010000011" => rgb <= "000000";
					when "01010001010000100" => rgb <= "000000";
					when "01010001010000101" => rgb <= "000000";
					when "01010001010000110" => rgb <= "000000";
					when "01010001010000111" => rgb <= "000000";
					when "01010001010001000" => rgb <= "100100";
					when "01010001010001001" => rgb <= "101000";
					when "01010001010001010" => rgb <= "101000";
					when "01010001010001011" => rgb <= "101000";
					when "01010001010001100" => rgb <= "101000";
					when "01010001010001101" => rgb <= "101000";
					when "01010001010001110" => rgb <= "101000";
					when "01010001010001111" => rgb <= "101000";
					when "01010001010010000" => rgb <= "101000";
					when "01010001010010001" => rgb <= "101000";
					when "01010001010010010" => rgb <= "101000";
					when "01010001010010011" => rgb <= "101000";
					when "01010001010010100" => rgb <= "101000";
					when "01010001010010101" => rgb <= "101000";
					when "01010001010010110" => rgb <= "101000";
					when "01010001010010111" => rgb <= "101000";
					when "01010001010011000" => rgb <= "101000";
					when "01010001010011001" => rgb <= "101000";
					when "01010001010011010" => rgb <= "101000";
					when "01010001010011011" => rgb <= "101000";
					when "01010001010011100" => rgb <= "101000";
					when "01010001010011101" => rgb <= "101000";
					when "01010001010011110" => rgb <= "101000";
					when "01010001010011111" => rgb <= "101000";
					when "01010001010100000" => rgb <= "101000";
					when "01010001010100001" => rgb <= "101000";
					when "01010001010100010" => rgb <= "101000";
					when "01010001010100011" => rgb <= "101000";
					when "01010001010100100" => rgb <= "101000";
					when "01010001010100101" => rgb <= "101000";
					when "01010001010100110" => rgb <= "101000";
					when "01010001010100111" => rgb <= "101000";
					when "01010001010101000" => rgb <= "101000";
					when "01010001010101001" => rgb <= "101000";
					when "01010001010101010" => rgb <= "101000";
					when "01010001010101011" => rgb <= "101000";
					when "01010001010101100" => rgb <= "101000";
					when "01010001010101101" => rgb <= "101000";
					when "01010001010101110" => rgb <= "101000";
					when "01010001010101111" => rgb <= "101000";
					when "01010001010110000" => rgb <= "101000";
					when "01010001010110001" => rgb <= "101000";
					when "01010001010110010" => rgb <= "101000";
					when "01010001010110011" => rgb <= "101000";
					when "01010001010110100" => rgb <= "101000";
					when "01010001010110101" => rgb <= "010100";
					when "01010001010110110" => rgb <= "000000";
					when "01010001010110111" => rgb <= "000000";
					when "01010001010111000" => rgb <= "000000";
					when "01010001010111001" => rgb <= "000000";
					when "01010001010111010" => rgb <= "000000";
					when "01010001010111011" => rgb <= "000000";
					when "01010001010111100" => rgb <= "000000";
					when "01010001010111101" => rgb <= "000000";
					when "01010001010111110" => rgb <= "000000";
					when "01010001010111111" => rgb <= "000000";
					when "01010001011000000" => rgb <= "000000";
					when "01010001011000001" => rgb <= "000000";
					when "01010001011000010" => rgb <= "000000";
					when "01010001011000011" => rgb <= "000000";
					when "01010001011000100" => rgb <= "000000";
					when "01010001011000101" => rgb <= "000000";
					when "01010001011000110" => rgb <= "000000";
					when "01010001011000111" => rgb <= "000000";
					when "01010001011001000" => rgb <= "000000";
					when "01010001011001001" => rgb <= "000000";
					when "01010001011001010" => rgb <= "000000";
					when "01010001011001011" => rgb <= "000000";
					when "01010001011001100" => rgb <= "000000";
					when "01010001011001101" => rgb <= "000000";
					when "01010001011001110" => rgb <= "000000";
					when "01010001011001111" => rgb <= "000000";
					when "01010001011010000" => rgb <= "000000";
					when "01010001011010001" => rgb <= "000000";
					when "01010001011010010" => rgb <= "000000";
					when "01010001011010011" => rgb <= "000000";
					when "01010001011010100" => rgb <= "000000";
					when "01010001011010101" => rgb <= "000000";
					when "01010001011010110" => rgb <= "000000";
					when "01010001011010111" => rgb <= "000000";
					when "01010001011011000" => rgb <= "000000";
					when "01010001011011001" => rgb <= "000000";
					when "01010001011011010" => rgb <= "000000";
					when "01010001011011011" => rgb <= "000000";
					when "01010001011011100" => rgb <= "000000";
					when "01010001011011101" => rgb <= "000000";
					when "01010001011011110" => rgb <= "000000";
					when "01010001011011111" => rgb <= "000000";
					when "01010001011100000" => rgb <= "000000";
					when "01010001011100001" => rgb <= "000000";
					when "01010001011100010" => rgb <= "000000";
					when "01010001011100011" => rgb <= "000000";
					when "01010001011100100" => rgb <= "000000";
					when "01010001011100101" => rgb <= "000000";
					when "01010001011100110" => rgb <= "000000";
					when "01010001011100111" => rgb <= "000000";
					when "01010001011101000" => rgb <= "000000";
					when "01010001011101001" => rgb <= "000000";
					when "01010001011101010" => rgb <= "000000";
					when "01010001011101011" => rgb <= "000000";
					when "01010001011101100" => rgb <= "000000";
					when "01010001011101101" => rgb <= "000000";
					when "01010001011101110" => rgb <= "000000";
					when "01010001011101111" => rgb <= "000000";
					when "01010001011110000" => rgb <= "000000";
					when "01010001011110001" => rgb <= "000000";
					when "01010001011110010" => rgb <= "000000";
					when "01010001011110011" => rgb <= "000000";
					when "01010001011110100" => rgb <= "000000";
					when "01010001011110101" => rgb <= "000000";
					when "01010001011110110" => rgb <= "000000";
					when "01010001011110111" => rgb <= "000000";
					when "01010001011111000" => rgb <= "000000";
					when "01010001011111001" => rgb <= "000000";
					when "01010001011111010" => rgb <= "000000";
					when "01010001011111011" => rgb <= "000000";
					when "01010001011111100" => rgb <= "000000";
					when "01010001011111101" => rgb <= "000000";
					when "01010001011111110" => rgb <= "000000";
					when "01010001011111111" => rgb <= "000000";
					when "01010001100000000" => rgb <= "000000";
					when "01010001100000001" => rgb <= "000000";
					when "01010001100000010" => rgb <= "000000";
					when "01010001100000011" => rgb <= "000000";
					when "01010001100000100" => rgb <= "000000";
					when "01010001100000101" => rgb <= "000000";
					when "01010001100000110" => rgb <= "000000";
					when "01010001100000111" => rgb <= "000000";
					when "01010001100001000" => rgb <= "000000";
					when "01010001100001001" => rgb <= "000000";
					when "01010001100001010" => rgb <= "000000";
					when "01010001100001011" => rgb <= "000000";
					when "01010001100001100" => rgb <= "000000";
					when "01010001100001101" => rgb <= "000000";
					when "01010001100001110" => rgb <= "000000";
					when "01010001100001111" => rgb <= "000000";
					when "01010001100010000" => rgb <= "000000";
					when "01010001100010001" => rgb <= "000000";
					when "01010001100010010" => rgb <= "000000";
					when "01010001100010011" => rgb <= "000000";
					when "01010001100010100" => rgb <= "000000";
					when "01010001100010101" => rgb <= "000000";
					when "01010001100010110" => rgb <= "000000";
					when "01010001100010111" => rgb <= "000000";
					when "01010001100011000" => rgb <= "000000";
					when "01010001100011001" => rgb <= "000000";
					when "01010001100011010" => rgb <= "000000";
					when "01010001100011011" => rgb <= "000000";
					when "01010001100011100" => rgb <= "000000";
					when "01010001100011101" => rgb <= "000000";
					when "01010001100011110" => rgb <= "000000";
					when "01010001100011111" => rgb <= "000000";
					when "01010001100100000" => rgb <= "000000";
					when "01010001100100001" => rgb <= "000000";
					when "01010001100100010" => rgb <= "000000";
					when "01010001100100011" => rgb <= "000000";
					when "01010001100100100" => rgb <= "000000";
					when "01010001100100101" => rgb <= "000000";
					when "01010001100100110" => rgb <= "000000";
					when "01010001100100111" => rgb <= "000000";
					when "01010001100101000" => rgb <= "000000";
					when "01010001100101001" => rgb <= "000000";
					when "01010001100101010" => rgb <= "000000";
					when "01010001100101011" => rgb <= "000000";
					when "01010001100101100" => rgb <= "000000";
					when "01010001100101101" => rgb <= "000000";
					when "01010001100101110" => rgb <= "000000";
					when "01010001100101111" => rgb <= "000000";
					when "01010001100110000" => rgb <= "000000";
					when "01010001100110001" => rgb <= "000000";
					when "01010001100110010" => rgb <= "000000";
					when "01010001100110011" => rgb <= "000000";
					when "01010001100110100" => rgb <= "000000";
					when "01010001100110101" => rgb <= "000000";
					when "01010001100110110" => rgb <= "000000";
					when "01010001100110111" => rgb <= "000000";
					when "01010001100111000" => rgb <= "000000";
					when "01010001100111001" => rgb <= "000000";
					when "01010001100111010" => rgb <= "000000";
					when "01010001100111011" => rgb <= "000000";
					when "01010001100111100" => rgb <= "000000";
					when "01010001100111101" => rgb <= "000000";
					when "01010001100111110" => rgb <= "000000";
					when "01010001100111111" => rgb <= "000000";
					when "01010010000000000" => rgb <= "000000";
					when "01010010000000001" => rgb <= "000000";
					when "01010010000000010" => rgb <= "000000";
					when "01010010000000011" => rgb <= "000000";
					when "01010010000000100" => rgb <= "000000";
					when "01010010000000101" => rgb <= "000000";
					when "01010010000000110" => rgb <= "000000";
					when "01010010000000111" => rgb <= "000000";
					when "01010010000001000" => rgb <= "000000";
					when "01010010000001001" => rgb <= "000000";
					when "01010010000001010" => rgb <= "000000";
					when "01010010000001011" => rgb <= "000000";
					when "01010010000001100" => rgb <= "000000";
					when "01010010000001101" => rgb <= "000000";
					when "01010010000001110" => rgb <= "000000";
					when "01010010000001111" => rgb <= "000000";
					when "01010010000010000" => rgb <= "000000";
					when "01010010000010001" => rgb <= "000000";
					when "01010010000010010" => rgb <= "000000";
					when "01010010000010011" => rgb <= "000000";
					when "01010010000010100" => rgb <= "000000";
					when "01010010000010101" => rgb <= "000000";
					when "01010010000010110" => rgb <= "000000";
					when "01010010000010111" => rgb <= "000000";
					when "01010010000011000" => rgb <= "000000";
					when "01010010000011001" => rgb <= "000000";
					when "01010010000011010" => rgb <= "000000";
					when "01010010000011011" => rgb <= "000000";
					when "01010010000011100" => rgb <= "000000";
					when "01010010000011101" => rgb <= "000000";
					when "01010010000011110" => rgb <= "000000";
					when "01010010000011111" => rgb <= "000000";
					when "01010010000100000" => rgb <= "000000";
					when "01010010000100001" => rgb <= "000000";
					when "01010010000100010" => rgb <= "000000";
					when "01010010000100011" => rgb <= "000000";
					when "01010010000100100" => rgb <= "000000";
					when "01010010000100101" => rgb <= "000000";
					when "01010010000100110" => rgb <= "000000";
					when "01010010000100111" => rgb <= "000000";
					when "01010010000101000" => rgb <= "000000";
					when "01010010000101001" => rgb <= "000000";
					when "01010010000101010" => rgb <= "000000";
					when "01010010000101011" => rgb <= "000000";
					when "01010010000101100" => rgb <= "000000";
					when "01010010000101101" => rgb <= "000000";
					when "01010010000101110" => rgb <= "000000";
					when "01010010000101111" => rgb <= "000000";
					when "01010010000110000" => rgb <= "000000";
					when "01010010000110001" => rgb <= "000000";
					when "01010010000110010" => rgb <= "000000";
					when "01010010000110011" => rgb <= "000000";
					when "01010010000110100" => rgb <= "000000";
					when "01010010000110101" => rgb <= "000000";
					when "01010010000110110" => rgb <= "000000";
					when "01010010000110111" => rgb <= "000000";
					when "01010010000111000" => rgb <= "000000";
					when "01010010000111001" => rgb <= "000000";
					when "01010010000111010" => rgb <= "000000";
					when "01010010000111011" => rgb <= "000000";
					when "01010010000111100" => rgb <= "000000";
					when "01010010000111101" => rgb <= "000000";
					when "01010010000111110" => rgb <= "000000";
					when "01010010000111111" => rgb <= "000000";
					when "01010010001000000" => rgb <= "000000";
					when "01010010001000001" => rgb <= "000000";
					when "01010010001000010" => rgb <= "000000";
					when "01010010001000011" => rgb <= "000000";
					when "01010010001000100" => rgb <= "000000";
					when "01010010001000101" => rgb <= "000000";
					when "01010010001000110" => rgb <= "000000";
					when "01010010001000111" => rgb <= "000000";
					when "01010010001001000" => rgb <= "000000";
					when "01010010001001001" => rgb <= "000000";
					when "01010010001001010" => rgb <= "000000";
					when "01010010001001011" => rgb <= "000000";
					when "01010010001001100" => rgb <= "000000";
					when "01010010001001101" => rgb <= "000000";
					when "01010010001001110" => rgb <= "000000";
					when "01010010001001111" => rgb <= "000000";
					when "01010010001010000" => rgb <= "000000";
					when "01010010001010001" => rgb <= "000000";
					when "01010010001010010" => rgb <= "000000";
					when "01010010001010011" => rgb <= "000000";
					when "01010010001010100" => rgb <= "000000";
					when "01010010001010101" => rgb <= "000000";
					when "01010010001010110" => rgb <= "000000";
					when "01010010001010111" => rgb <= "000000";
					when "01010010001011000" => rgb <= "000000";
					when "01010010001011001" => rgb <= "000000";
					when "01010010001011010" => rgb <= "000000";
					when "01010010001011011" => rgb <= "000000";
					when "01010010001011100" => rgb <= "000000";
					when "01010010001011101" => rgb <= "000000";
					when "01010010001011110" => rgb <= "000000";
					when "01010010001011111" => rgb <= "000000";
					when "01010010001100000" => rgb <= "000000";
					when "01010010001100001" => rgb <= "000000";
					when "01010010001100010" => rgb <= "000000";
					when "01010010001100011" => rgb <= "000000";
					when "01010010001100100" => rgb <= "000000";
					when "01010010001100101" => rgb <= "000000";
					when "01010010001100110" => rgb <= "000000";
					when "01010010001100111" => rgb <= "000000";
					when "01010010001101000" => rgb <= "000000";
					when "01010010001101001" => rgb <= "000000";
					when "01010010001101010" => rgb <= "000000";
					when "01010010001101011" => rgb <= "000000";
					when "01010010001101100" => rgb <= "000000";
					when "01010010001101101" => rgb <= "000000";
					when "01010010001101110" => rgb <= "000000";
					when "01010010001101111" => rgb <= "000000";
					when "01010010001110000" => rgb <= "000000";
					when "01010010001110001" => rgb <= "000000";
					when "01010010001110010" => rgb <= "000000";
					when "01010010001110011" => rgb <= "000000";
					when "01010010001110100" => rgb <= "000000";
					when "01010010001110101" => rgb <= "000000";
					when "01010010001110110" => rgb <= "000000";
					when "01010010001110111" => rgb <= "000000";
					when "01010010001111000" => rgb <= "000000";
					when "01010010001111001" => rgb <= "000000";
					when "01010010001111010" => rgb <= "000000";
					when "01010010001111011" => rgb <= "000000";
					when "01010010001111100" => rgb <= "000000";
					when "01010010001111101" => rgb <= "000000";
					when "01010010001111110" => rgb <= "000000";
					when "01010010001111111" => rgb <= "000000";
					when "01010010010000000" => rgb <= "000000";
					when "01010010010000001" => rgb <= "000000";
					when "01010010010000010" => rgb <= "000000";
					when "01010010010000011" => rgb <= "000000";
					when "01010010010000100" => rgb <= "000000";
					when "01010010010000101" => rgb <= "000000";
					when "01010010010000110" => rgb <= "000000";
					when "01010010010000111" => rgb <= "000000";
					when "01010010010001000" => rgb <= "100100";
					when "01010010010001001" => rgb <= "101000";
					when "01010010010001010" => rgb <= "101000";
					when "01010010010001011" => rgb <= "101000";
					when "01010010010001100" => rgb <= "101000";
					when "01010010010001101" => rgb <= "101000";
					when "01010010010001110" => rgb <= "101000";
					when "01010010010001111" => rgb <= "101000";
					when "01010010010010000" => rgb <= "101000";
					when "01010010010010001" => rgb <= "101000";
					when "01010010010010010" => rgb <= "101000";
					when "01010010010010011" => rgb <= "101000";
					when "01010010010010100" => rgb <= "101000";
					when "01010010010010101" => rgb <= "101000";
					when "01010010010010110" => rgb <= "101000";
					when "01010010010010111" => rgb <= "111000";
					when "01010010010011000" => rgb <= "101000";
					when "01010010010011001" => rgb <= "101000";
					when "01010010010011010" => rgb <= "101000";
					when "01010010010011011" => rgb <= "101000";
					when "01010010010011100" => rgb <= "101000";
					when "01010010010011101" => rgb <= "101000";
					when "01010010010011110" => rgb <= "101000";
					when "01010010010011111" => rgb <= "101000";
					when "01010010010100000" => rgb <= "101000";
					when "01010010010100001" => rgb <= "101000";
					when "01010010010100010" => rgb <= "101000";
					when "01010010010100011" => rgb <= "101000";
					when "01010010010100100" => rgb <= "101000";
					when "01010010010100101" => rgb <= "101000";
					when "01010010010100110" => rgb <= "101000";
					when "01010010010100111" => rgb <= "101000";
					when "01010010010101000" => rgb <= "101000";
					when "01010010010101001" => rgb <= "101000";
					when "01010010010101010" => rgb <= "101000";
					when "01010010010101011" => rgb <= "101000";
					when "01010010010101100" => rgb <= "101000";
					when "01010010010101101" => rgb <= "101000";
					when "01010010010101110" => rgb <= "101000";
					when "01010010010101111" => rgb <= "101000";
					when "01010010010110000" => rgb <= "101000";
					when "01010010010110001" => rgb <= "101000";
					when "01010010010110010" => rgb <= "101000";
					when "01010010010110011" => rgb <= "101000";
					when "01010010010110100" => rgb <= "101000";
					when "01010010010110101" => rgb <= "010100";
					when "01010010010110110" => rgb <= "000000";
					when "01010010010110111" => rgb <= "000000";
					when "01010010010111000" => rgb <= "000000";
					when "01010010010111001" => rgb <= "000000";
					when "01010010010111010" => rgb <= "000000";
					when "01010010010111011" => rgb <= "000000";
					when "01010010010111100" => rgb <= "000000";
					when "01010010010111101" => rgb <= "000000";
					when "01010010010111110" => rgb <= "000000";
					when "01010010010111111" => rgb <= "000000";
					when "01010010011000000" => rgb <= "000000";
					when "01010010011000001" => rgb <= "000000";
					when "01010010011000010" => rgb <= "000000";
					when "01010010011000011" => rgb <= "000000";
					when "01010010011000100" => rgb <= "000000";
					when "01010010011000101" => rgb <= "000000";
					when "01010010011000110" => rgb <= "000000";
					when "01010010011000111" => rgb <= "000000";
					when "01010010011001000" => rgb <= "000000";
					when "01010010011001001" => rgb <= "000000";
					when "01010010011001010" => rgb <= "000000";
					when "01010010011001011" => rgb <= "000000";
					when "01010010011001100" => rgb <= "000000";
					when "01010010011001101" => rgb <= "000000";
					when "01010010011001110" => rgb <= "000000";
					when "01010010011001111" => rgb <= "000000";
					when "01010010011010000" => rgb <= "000000";
					when "01010010011010001" => rgb <= "000000";
					when "01010010011010010" => rgb <= "000000";
					when "01010010011010011" => rgb <= "000000";
					when "01010010011010100" => rgb <= "000000";
					when "01010010011010101" => rgb <= "000000";
					when "01010010011010110" => rgb <= "000000";
					when "01010010011010111" => rgb <= "000000";
					when "01010010011011000" => rgb <= "000000";
					when "01010010011011001" => rgb <= "000000";
					when "01010010011011010" => rgb <= "000000";
					when "01010010011011011" => rgb <= "000000";
					when "01010010011011100" => rgb <= "000000";
					when "01010010011011101" => rgb <= "000000";
					when "01010010011011110" => rgb <= "000000";
					when "01010010011011111" => rgb <= "000000";
					when "01010010011100000" => rgb <= "000000";
					when "01010010011100001" => rgb <= "000000";
					when "01010010011100010" => rgb <= "000000";
					when "01010010011100011" => rgb <= "000000";
					when "01010010011100100" => rgb <= "000000";
					when "01010010011100101" => rgb <= "000000";
					when "01010010011100110" => rgb <= "000000";
					when "01010010011100111" => rgb <= "000000";
					when "01010010011101000" => rgb <= "000000";
					when "01010010011101001" => rgb <= "000000";
					when "01010010011101010" => rgb <= "000000";
					when "01010010011101011" => rgb <= "000000";
					when "01010010011101100" => rgb <= "000000";
					when "01010010011101101" => rgb <= "000000";
					when "01010010011101110" => rgb <= "000000";
					when "01010010011101111" => rgb <= "000000";
					when "01010010011110000" => rgb <= "000000";
					when "01010010011110001" => rgb <= "000000";
					when "01010010011110010" => rgb <= "000000";
					when "01010010011110011" => rgb <= "000000";
					when "01010010011110100" => rgb <= "000000";
					when "01010010011110101" => rgb <= "000000";
					when "01010010011110110" => rgb <= "000000";
					when "01010010011110111" => rgb <= "000000";
					when "01010010011111000" => rgb <= "000000";
					when "01010010011111001" => rgb <= "000000";
					when "01010010011111010" => rgb <= "000000";
					when "01010010011111011" => rgb <= "000000";
					when "01010010011111100" => rgb <= "000000";
					when "01010010011111101" => rgb <= "000000";
					when "01010010011111110" => rgb <= "000000";
					when "01010010011111111" => rgb <= "000000";
					when "01010010100000000" => rgb <= "000000";
					when "01010010100000001" => rgb <= "000000";
					when "01010010100000010" => rgb <= "000000";
					when "01010010100000011" => rgb <= "000000";
					when "01010010100000100" => rgb <= "000000";
					when "01010010100000101" => rgb <= "000000";
					when "01010010100000110" => rgb <= "000000";
					when "01010010100000111" => rgb <= "000000";
					when "01010010100001000" => rgb <= "000000";
					when "01010010100001001" => rgb <= "000000";
					when "01010010100001010" => rgb <= "000000";
					when "01010010100001011" => rgb <= "000000";
					when "01010010100001100" => rgb <= "000000";
					when "01010010100001101" => rgb <= "000000";
					when "01010010100001110" => rgb <= "000000";
					when "01010010100001111" => rgb <= "000000";
					when "01010010100010000" => rgb <= "000000";
					when "01010010100010001" => rgb <= "000000";
					when "01010010100010010" => rgb <= "000000";
					when "01010010100010011" => rgb <= "000000";
					when "01010010100010100" => rgb <= "000000";
					when "01010010100010101" => rgb <= "000000";
					when "01010010100010110" => rgb <= "000000";
					when "01010010100010111" => rgb <= "000000";
					when "01010010100011000" => rgb <= "000000";
					when "01010010100011001" => rgb <= "000000";
					when "01010010100011010" => rgb <= "000000";
					when "01010010100011011" => rgb <= "000000";
					when "01010010100011100" => rgb <= "000000";
					when "01010010100011101" => rgb <= "000000";
					when "01010010100011110" => rgb <= "000000";
					when "01010010100011111" => rgb <= "000000";
					when "01010010100100000" => rgb <= "000000";
					when "01010010100100001" => rgb <= "000000";
					when "01010010100100010" => rgb <= "000000";
					when "01010010100100011" => rgb <= "000000";
					when "01010010100100100" => rgb <= "000000";
					when "01010010100100101" => rgb <= "000000";
					when "01010010100100110" => rgb <= "000000";
					when "01010010100100111" => rgb <= "000000";
					when "01010010100101000" => rgb <= "000000";
					when "01010010100101001" => rgb <= "000000";
					when "01010010100101010" => rgb <= "000000";
					when "01010010100101011" => rgb <= "000000";
					when "01010010100101100" => rgb <= "000000";
					when "01010010100101101" => rgb <= "000000";
					when "01010010100101110" => rgb <= "000000";
					when "01010010100101111" => rgb <= "000000";
					when "01010010100110000" => rgb <= "000000";
					when "01010010100110001" => rgb <= "000000";
					when "01010010100110010" => rgb <= "000000";
					when "01010010100110011" => rgb <= "000000";
					when "01010010100110100" => rgb <= "000000";
					when "01010010100110101" => rgb <= "000000";
					when "01010010100110110" => rgb <= "000000";
					when "01010010100110111" => rgb <= "000000";
					when "01010010100111000" => rgb <= "000000";
					when "01010010100111001" => rgb <= "000000";
					when "01010010100111010" => rgb <= "000000";
					when "01010010100111011" => rgb <= "000000";
					when "01010010100111100" => rgb <= "000000";
					when "01010010100111101" => rgb <= "000000";
					when "01010010100111110" => rgb <= "000000";
					when "01010010100111111" => rgb <= "000000";
					when "01010011000000000" => rgb <= "000000";
					when "01010011000000001" => rgb <= "000000";
					when "01010011000000010" => rgb <= "000000";
					when "01010011000000011" => rgb <= "000000";
					when "01010011000000100" => rgb <= "000000";
					when "01010011000000101" => rgb <= "000000";
					when "01010011000000110" => rgb <= "000000";
					when "01010011000000111" => rgb <= "000000";
					when "01010011000001000" => rgb <= "000000";
					when "01010011000001001" => rgb <= "000000";
					when "01010011000001010" => rgb <= "000000";
					when "01010011000001011" => rgb <= "000000";
					when "01010011000001100" => rgb <= "000000";
					when "01010011000001101" => rgb <= "000000";
					when "01010011000001110" => rgb <= "000000";
					when "01010011000001111" => rgb <= "000000";
					when "01010011000010000" => rgb <= "000000";
					when "01010011000010001" => rgb <= "000000";
					when "01010011000010010" => rgb <= "000000";
					when "01010011000010011" => rgb <= "000000";
					when "01010011000010100" => rgb <= "000000";
					when "01010011000010101" => rgb <= "000000";
					when "01010011000010110" => rgb <= "000000";
					when "01010011000010111" => rgb <= "000000";
					when "01010011000011000" => rgb <= "000000";
					when "01010011000011001" => rgb <= "000000";
					when "01010011000011010" => rgb <= "000000";
					when "01010011000011011" => rgb <= "000000";
					when "01010011000011100" => rgb <= "000000";
					when "01010011000011101" => rgb <= "000000";
					when "01010011000011110" => rgb <= "000000";
					when "01010011000011111" => rgb <= "000000";
					when "01010011000100000" => rgb <= "000000";
					when "01010011000100001" => rgb <= "000000";
					when "01010011000100010" => rgb <= "000000";
					when "01010011000100011" => rgb <= "000000";
					when "01010011000100100" => rgb <= "000000";
					when "01010011000100101" => rgb <= "000000";
					when "01010011000100110" => rgb <= "000000";
					when "01010011000100111" => rgb <= "000000";
					when "01010011000101000" => rgb <= "000000";
					when "01010011000101001" => rgb <= "000000";
					when "01010011000101010" => rgb <= "000000";
					when "01010011000101011" => rgb <= "000000";
					when "01010011000101100" => rgb <= "000000";
					when "01010011000101101" => rgb <= "000000";
					when "01010011000101110" => rgb <= "000000";
					when "01010011000101111" => rgb <= "000000";
					when "01010011000110000" => rgb <= "000000";
					when "01010011000110001" => rgb <= "000000";
					when "01010011000110010" => rgb <= "000000";
					when "01010011000110011" => rgb <= "000000";
					when "01010011000110100" => rgb <= "000000";
					when "01010011000110101" => rgb <= "000000";
					when "01010011000110110" => rgb <= "000000";
					when "01010011000110111" => rgb <= "000000";
					when "01010011000111000" => rgb <= "000000";
					when "01010011000111001" => rgb <= "000000";
					when "01010011000111010" => rgb <= "000000";
					when "01010011000111011" => rgb <= "000000";
					when "01010011000111100" => rgb <= "000000";
					when "01010011000111101" => rgb <= "000000";
					when "01010011000111110" => rgb <= "000000";
					when "01010011000111111" => rgb <= "000000";
					when "01010011001000000" => rgb <= "000000";
					when "01010011001000001" => rgb <= "000000";
					when "01010011001000010" => rgb <= "000000";
					when "01010011001000011" => rgb <= "000000";
					when "01010011001000100" => rgb <= "000000";
					when "01010011001000101" => rgb <= "000000";
					when "01010011001000110" => rgb <= "000000";
					when "01010011001000111" => rgb <= "000000";
					when "01010011001001000" => rgb <= "000000";
					when "01010011001001001" => rgb <= "000000";
					when "01010011001001010" => rgb <= "000000";
					when "01010011001001011" => rgb <= "000000";
					when "01010011001001100" => rgb <= "000000";
					when "01010011001001101" => rgb <= "000000";
					when "01010011001001110" => rgb <= "000000";
					when "01010011001001111" => rgb <= "000000";
					when "01010011001010000" => rgb <= "000000";
					when "01010011001010001" => rgb <= "000000";
					when "01010011001010010" => rgb <= "000000";
					when "01010011001010011" => rgb <= "000000";
					when "01010011001010100" => rgb <= "000000";
					when "01010011001010101" => rgb <= "000000";
					when "01010011001010110" => rgb <= "000000";
					when "01010011001010111" => rgb <= "000000";
					when "01010011001011000" => rgb <= "000000";
					when "01010011001011001" => rgb <= "000000";
					when "01010011001011010" => rgb <= "000000";
					when "01010011001011011" => rgb <= "000000";
					when "01010011001011100" => rgb <= "000000";
					when "01010011001011101" => rgb <= "000000";
					when "01010011001011110" => rgb <= "000000";
					when "01010011001011111" => rgb <= "000000";
					when "01010011001100000" => rgb <= "000000";
					when "01010011001100001" => rgb <= "000000";
					when "01010011001100010" => rgb <= "000000";
					when "01010011001100011" => rgb <= "000000";
					when "01010011001100100" => rgb <= "000000";
					when "01010011001100101" => rgb <= "000000";
					when "01010011001100110" => rgb <= "000000";
					when "01010011001100111" => rgb <= "000000";
					when "01010011001101000" => rgb <= "000000";
					when "01010011001101001" => rgb <= "000000";
					when "01010011001101010" => rgb <= "000000";
					when "01010011001101011" => rgb <= "000000";
					when "01010011001101100" => rgb <= "000000";
					when "01010011001101101" => rgb <= "000000";
					when "01010011001101110" => rgb <= "000000";
					when "01010011001101111" => rgb <= "000000";
					when "01010011001110000" => rgb <= "000000";
					when "01010011001110001" => rgb <= "000000";
					when "01010011001110010" => rgb <= "000000";
					when "01010011001110011" => rgb <= "000000";
					when "01010011001110100" => rgb <= "000000";
					when "01010011001110101" => rgb <= "000000";
					when "01010011001110110" => rgb <= "000000";
					when "01010011001110111" => rgb <= "000000";
					when "01010011001111000" => rgb <= "000000";
					when "01010011001111001" => rgb <= "000000";
					when "01010011001111010" => rgb <= "000000";
					when "01010011001111011" => rgb <= "000000";
					when "01010011001111100" => rgb <= "000000";
					when "01010011001111101" => rgb <= "000000";
					when "01010011001111110" => rgb <= "000000";
					when "01010011001111111" => rgb <= "000000";
					when "01010011010000000" => rgb <= "000000";
					when "01010011010000001" => rgb <= "000000";
					when "01010011010000010" => rgb <= "000000";
					when "01010011010000011" => rgb <= "000000";
					when "01010011010000100" => rgb <= "000000";
					when "01010011010000101" => rgb <= "000000";
					when "01010011010000110" => rgb <= "000000";
					when "01010011010000111" => rgb <= "000000";
					when "01010011010001000" => rgb <= "100100";
					when "01010011010001001" => rgb <= "101000";
					when "01010011010001010" => rgb <= "101000";
					when "01010011010001011" => rgb <= "101000";
					when "01010011010001100" => rgb <= "101000";
					when "01010011010001101" => rgb <= "101000";
					when "01010011010001110" => rgb <= "101000";
					when "01010011010001111" => rgb <= "101000";
					when "01010011010010000" => rgb <= "111001";
					when "01010011010010001" => rgb <= "101000";
					when "01010011010010010" => rgb <= "101000";
					when "01010011010010011" => rgb <= "101000";
					when "01010011010010100" => rgb <= "101000";
					when "01010011010010101" => rgb <= "101000";
					when "01010011010010110" => rgb <= "101000";
					when "01010011010010111" => rgb <= "101000";
					when "01010011010011000" => rgb <= "101000";
					when "01010011010011001" => rgb <= "101000";
					when "01010011010011010" => rgb <= "101000";
					when "01010011010011011" => rgb <= "101000";
					when "01010011010011100" => rgb <= "101000";
					when "01010011010011101" => rgb <= "101000";
					when "01010011010011110" => rgb <= "101000";
					when "01010011010011111" => rgb <= "101000";
					when "01010011010100000" => rgb <= "101000";
					when "01010011010100001" => rgb <= "101000";
					when "01010011010100010" => rgb <= "101000";
					when "01010011010100011" => rgb <= "101000";
					when "01010011010100100" => rgb <= "101000";
					when "01010011010100101" => rgb <= "101000";
					when "01010011010100110" => rgb <= "101000";
					when "01010011010100111" => rgb <= "101000";
					when "01010011010101000" => rgb <= "101000";
					when "01010011010101001" => rgb <= "101000";
					when "01010011010101010" => rgb <= "101000";
					when "01010011010101011" => rgb <= "101000";
					when "01010011010101100" => rgb <= "101000";
					when "01010011010101101" => rgb <= "101000";
					when "01010011010101110" => rgb <= "101000";
					when "01010011010101111" => rgb <= "101000";
					when "01010011010110000" => rgb <= "101000";
					when "01010011010110001" => rgb <= "101000";
					when "01010011010110010" => rgb <= "101000";
					when "01010011010110011" => rgb <= "101000";
					when "01010011010110100" => rgb <= "101000";
					when "01010011010110101" => rgb <= "010100";
					when "01010011010110110" => rgb <= "000000";
					when "01010011010110111" => rgb <= "000000";
					when "01010011010111000" => rgb <= "000000";
					when "01010011010111001" => rgb <= "000000";
					when "01010011010111010" => rgb <= "000000";
					when "01010011010111011" => rgb <= "000000";
					when "01010011010111100" => rgb <= "000000";
					when "01010011010111101" => rgb <= "000000";
					when "01010011010111110" => rgb <= "000000";
					when "01010011010111111" => rgb <= "000000";
					when "01010011011000000" => rgb <= "000000";
					when "01010011011000001" => rgb <= "000000";
					when "01010011011000010" => rgb <= "000000";
					when "01010011011000011" => rgb <= "000000";
					when "01010011011000100" => rgb <= "000000";
					when "01010011011000101" => rgb <= "000000";
					when "01010011011000110" => rgb <= "000000";
					when "01010011011000111" => rgb <= "000000";
					when "01010011011001000" => rgb <= "000000";
					when "01010011011001001" => rgb <= "000000";
					when "01010011011001010" => rgb <= "000000";
					when "01010011011001011" => rgb <= "000000";
					when "01010011011001100" => rgb <= "000000";
					when "01010011011001101" => rgb <= "000000";
					when "01010011011001110" => rgb <= "000000";
					when "01010011011001111" => rgb <= "000000";
					when "01010011011010000" => rgb <= "000000";
					when "01010011011010001" => rgb <= "000000";
					when "01010011011010010" => rgb <= "000000";
					when "01010011011010011" => rgb <= "000000";
					when "01010011011010100" => rgb <= "000000";
					when "01010011011010101" => rgb <= "000000";
					when "01010011011010110" => rgb <= "000000";
					when "01010011011010111" => rgb <= "000000";
					when "01010011011011000" => rgb <= "000000";
					when "01010011011011001" => rgb <= "000000";
					when "01010011011011010" => rgb <= "000000";
					when "01010011011011011" => rgb <= "000000";
					when "01010011011011100" => rgb <= "000000";
					when "01010011011011101" => rgb <= "000000";
					when "01010011011011110" => rgb <= "000000";
					when "01010011011011111" => rgb <= "000000";
					when "01010011011100000" => rgb <= "000000";
					when "01010011011100001" => rgb <= "000000";
					when "01010011011100010" => rgb <= "000000";
					when "01010011011100011" => rgb <= "000000";
					when "01010011011100100" => rgb <= "000000";
					when "01010011011100101" => rgb <= "000000";
					when "01010011011100110" => rgb <= "000000";
					when "01010011011100111" => rgb <= "000000";
					when "01010011011101000" => rgb <= "000000";
					when "01010011011101001" => rgb <= "000000";
					when "01010011011101010" => rgb <= "000000";
					when "01010011011101011" => rgb <= "000000";
					when "01010011011101100" => rgb <= "000000";
					when "01010011011101101" => rgb <= "000000";
					when "01010011011101110" => rgb <= "000000";
					when "01010011011101111" => rgb <= "000000";
					when "01010011011110000" => rgb <= "000000";
					when "01010011011110001" => rgb <= "000000";
					when "01010011011110010" => rgb <= "000000";
					when "01010011011110011" => rgb <= "000000";
					when "01010011011110100" => rgb <= "000000";
					when "01010011011110101" => rgb <= "000000";
					when "01010011011110110" => rgb <= "000000";
					when "01010011011110111" => rgb <= "000000";
					when "01010011011111000" => rgb <= "000000";
					when "01010011011111001" => rgb <= "000000";
					when "01010011011111010" => rgb <= "000000";
					when "01010011011111011" => rgb <= "000000";
					when "01010011011111100" => rgb <= "000000";
					when "01010011011111101" => rgb <= "000000";
					when "01010011011111110" => rgb <= "000000";
					when "01010011011111111" => rgb <= "000000";
					when "01010011100000000" => rgb <= "000000";
					when "01010011100000001" => rgb <= "000000";
					when "01010011100000010" => rgb <= "000000";
					when "01010011100000011" => rgb <= "000000";
					when "01010011100000100" => rgb <= "000000";
					when "01010011100000101" => rgb <= "000000";
					when "01010011100000110" => rgb <= "000000";
					when "01010011100000111" => rgb <= "000000";
					when "01010011100001000" => rgb <= "000000";
					when "01010011100001001" => rgb <= "000000";
					when "01010011100001010" => rgb <= "000000";
					when "01010011100001011" => rgb <= "000000";
					when "01010011100001100" => rgb <= "000000";
					when "01010011100001101" => rgb <= "000000";
					when "01010011100001110" => rgb <= "000000";
					when "01010011100001111" => rgb <= "000000";
					when "01010011100010000" => rgb <= "000000";
					when "01010011100010001" => rgb <= "000000";
					when "01010011100010010" => rgb <= "000000";
					when "01010011100010011" => rgb <= "000000";
					when "01010011100010100" => rgb <= "000000";
					when "01010011100010101" => rgb <= "000000";
					when "01010011100010110" => rgb <= "000000";
					when "01010011100010111" => rgb <= "000000";
					when "01010011100011000" => rgb <= "000000";
					when "01010011100011001" => rgb <= "000000";
					when "01010011100011010" => rgb <= "000000";
					when "01010011100011011" => rgb <= "000000";
					when "01010011100011100" => rgb <= "000000";
					when "01010011100011101" => rgb <= "000000";
					when "01010011100011110" => rgb <= "000000";
					when "01010011100011111" => rgb <= "000000";
					when "01010011100100000" => rgb <= "000000";
					when "01010011100100001" => rgb <= "000000";
					when "01010011100100010" => rgb <= "000000";
					when "01010011100100011" => rgb <= "000000";
					when "01010011100100100" => rgb <= "000000";
					when "01010011100100101" => rgb <= "000000";
					when "01010011100100110" => rgb <= "000000";
					when "01010011100100111" => rgb <= "000000";
					when "01010011100101000" => rgb <= "000000";
					when "01010011100101001" => rgb <= "000000";
					when "01010011100101010" => rgb <= "000000";
					when "01010011100101011" => rgb <= "000000";
					when "01010011100101100" => rgb <= "000000";
					when "01010011100101101" => rgb <= "000000";
					when "01010011100101110" => rgb <= "000000";
					when "01010011100101111" => rgb <= "000000";
					when "01010011100110000" => rgb <= "000000";
					when "01010011100110001" => rgb <= "000000";
					when "01010011100110010" => rgb <= "000000";
					when "01010011100110011" => rgb <= "000000";
					when "01010011100110100" => rgb <= "000000";
					when "01010011100110101" => rgb <= "000000";
					when "01010011100110110" => rgb <= "000000";
					when "01010011100110111" => rgb <= "000000";
					when "01010011100111000" => rgb <= "000000";
					when "01010011100111001" => rgb <= "000000";
					when "01010011100111010" => rgb <= "000000";
					when "01010011100111011" => rgb <= "000000";
					when "01010011100111100" => rgb <= "000000";
					when "01010011100111101" => rgb <= "000000";
					when "01010011100111110" => rgb <= "000000";
					when "01010011100111111" => rgb <= "000000";
					when "01010100000000000" => rgb <= "000000";
					when "01010100000000001" => rgb <= "000000";
					when "01010100000000010" => rgb <= "000000";
					when "01010100000000011" => rgb <= "000000";
					when "01010100000000100" => rgb <= "000000";
					when "01010100000000101" => rgb <= "000000";
					when "01010100000000110" => rgb <= "000000";
					when "01010100000000111" => rgb <= "000000";
					when "01010100000001000" => rgb <= "000000";
					when "01010100000001001" => rgb <= "000000";
					when "01010100000001010" => rgb <= "000000";
					when "01010100000001011" => rgb <= "000000";
					when "01010100000001100" => rgb <= "000000";
					when "01010100000001101" => rgb <= "000000";
					when "01010100000001110" => rgb <= "000000";
					when "01010100000001111" => rgb <= "000000";
					when "01010100000010000" => rgb <= "000000";
					when "01010100000010001" => rgb <= "000000";
					when "01010100000010010" => rgb <= "000000";
					when "01010100000010011" => rgb <= "000000";
					when "01010100000010100" => rgb <= "000000";
					when "01010100000010101" => rgb <= "000000";
					when "01010100000010110" => rgb <= "000000";
					when "01010100000010111" => rgb <= "000000";
					when "01010100000011000" => rgb <= "000000";
					when "01010100000011001" => rgb <= "000000";
					when "01010100000011010" => rgb <= "000000";
					when "01010100000011011" => rgb <= "000000";
					when "01010100000011100" => rgb <= "000000";
					when "01010100000011101" => rgb <= "000000";
					when "01010100000011110" => rgb <= "000000";
					when "01010100000011111" => rgb <= "000000";
					when "01010100000100000" => rgb <= "000000";
					when "01010100000100001" => rgb <= "000000";
					when "01010100000100010" => rgb <= "000000";
					when "01010100000100011" => rgb <= "000000";
					when "01010100000100100" => rgb <= "000000";
					when "01010100000100101" => rgb <= "000000";
					when "01010100000100110" => rgb <= "000000";
					when "01010100000100111" => rgb <= "000000";
					when "01010100000101000" => rgb <= "000000";
					when "01010100000101001" => rgb <= "000000";
					when "01010100000101010" => rgb <= "000000";
					when "01010100000101011" => rgb <= "000000";
					when "01010100000101100" => rgb <= "000000";
					when "01010100000101101" => rgb <= "000000";
					when "01010100000101110" => rgb <= "000000";
					when "01010100000101111" => rgb <= "000000";
					when "01010100000110000" => rgb <= "000000";
					when "01010100000110001" => rgb <= "000000";
					when "01010100000110010" => rgb <= "000000";
					when "01010100000110011" => rgb <= "000000";
					when "01010100000110100" => rgb <= "000000";
					when "01010100000110101" => rgb <= "000000";
					when "01010100000110110" => rgb <= "000000";
					when "01010100000110111" => rgb <= "000000";
					when "01010100000111000" => rgb <= "000000";
					when "01010100000111001" => rgb <= "000000";
					when "01010100000111010" => rgb <= "000000";
					when "01010100000111011" => rgb <= "000000";
					when "01010100000111100" => rgb <= "000000";
					when "01010100000111101" => rgb <= "000000";
					when "01010100000111110" => rgb <= "000000";
					when "01010100000111111" => rgb <= "000000";
					when "01010100001000000" => rgb <= "000000";
					when "01010100001000001" => rgb <= "000000";
					when "01010100001000010" => rgb <= "000000";
					when "01010100001000011" => rgb <= "000000";
					when "01010100001000100" => rgb <= "000000";
					when "01010100001000101" => rgb <= "000000";
					when "01010100001000110" => rgb <= "000000";
					when "01010100001000111" => rgb <= "000000";
					when "01010100001001000" => rgb <= "000000";
					when "01010100001001001" => rgb <= "000000";
					when "01010100001001010" => rgb <= "000000";
					when "01010100001001011" => rgb <= "000000";
					when "01010100001001100" => rgb <= "000000";
					when "01010100001001101" => rgb <= "000000";
					when "01010100001001110" => rgb <= "000000";
					when "01010100001001111" => rgb <= "000000";
					when "01010100001010000" => rgb <= "000000";
					when "01010100001010001" => rgb <= "000000";
					when "01010100001010010" => rgb <= "000000";
					when "01010100001010011" => rgb <= "000000";
					when "01010100001010100" => rgb <= "000000";
					when "01010100001010101" => rgb <= "000000";
					when "01010100001010110" => rgb <= "000000";
					when "01010100001010111" => rgb <= "000000";
					when "01010100001011000" => rgb <= "000000";
					when "01010100001011001" => rgb <= "000000";
					when "01010100001011010" => rgb <= "000000";
					when "01010100001011011" => rgb <= "000000";
					when "01010100001011100" => rgb <= "000000";
					when "01010100001011101" => rgb <= "000000";
					when "01010100001011110" => rgb <= "000000";
					when "01010100001011111" => rgb <= "000000";
					when "01010100001100000" => rgb <= "000000";
					when "01010100001100001" => rgb <= "000000";
					when "01010100001100010" => rgb <= "000000";
					when "01010100001100011" => rgb <= "000000";
					when "01010100001100100" => rgb <= "000000";
					when "01010100001100101" => rgb <= "000000";
					when "01010100001100110" => rgb <= "000000";
					when "01010100001100111" => rgb <= "000000";
					when "01010100001101000" => rgb <= "000000";
					when "01010100001101001" => rgb <= "000000";
					when "01010100001101010" => rgb <= "000000";
					when "01010100001101011" => rgb <= "000000";
					when "01010100001101100" => rgb <= "000000";
					when "01010100001101101" => rgb <= "000000";
					when "01010100001101110" => rgb <= "000000";
					when "01010100001101111" => rgb <= "000000";
					when "01010100001110000" => rgb <= "000000";
					when "01010100001110001" => rgb <= "000000";
					when "01010100001110010" => rgb <= "000000";
					when "01010100001110011" => rgb <= "000000";
					when "01010100001110100" => rgb <= "000000";
					when "01010100001110101" => rgb <= "000000";
					when "01010100001110110" => rgb <= "000000";
					when "01010100001110111" => rgb <= "000000";
					when "01010100001111000" => rgb <= "000000";
					when "01010100001111001" => rgb <= "000000";
					when "01010100001111010" => rgb <= "000000";
					when "01010100001111011" => rgb <= "000000";
					when "01010100001111100" => rgb <= "000000";
					when "01010100001111101" => rgb <= "000000";
					when "01010100001111110" => rgb <= "000000";
					when "01010100001111111" => rgb <= "000000";
					when "01010100010000000" => rgb <= "000000";
					when "01010100010000001" => rgb <= "000000";
					when "01010100010000010" => rgb <= "000000";
					when "01010100010000011" => rgb <= "000000";
					when "01010100010000100" => rgb <= "000000";
					when "01010100010000101" => rgb <= "000000";
					when "01010100010000110" => rgb <= "000000";
					when "01010100010000111" => rgb <= "000000";
					when "01010100010001000" => rgb <= "100100";
					when "01010100010001001" => rgb <= "101000";
					when "01010100010001010" => rgb <= "101000";
					when "01010100010001011" => rgb <= "101000";
					when "01010100010001100" => rgb <= "101000";
					when "01010100010001101" => rgb <= "101000";
					when "01010100010001110" => rgb <= "101000";
					when "01010100010001111" => rgb <= "101000";
					when "01010100010010000" => rgb <= "101000";
					when "01010100010010001" => rgb <= "101000";
					when "01010100010010010" => rgb <= "101000";
					when "01010100010010011" => rgb <= "101000";
					when "01010100010010100" => rgb <= "101000";
					when "01010100010010101" => rgb <= "101000";
					when "01010100010010110" => rgb <= "101000";
					when "01010100010010111" => rgb <= "101000";
					when "01010100010011000" => rgb <= "101000";
					when "01010100010011001" => rgb <= "101000";
					when "01010100010011010" => rgb <= "101000";
					when "01010100010011011" => rgb <= "101000";
					when "01010100010011100" => rgb <= "101000";
					when "01010100010011101" => rgb <= "101000";
					when "01010100010011110" => rgb <= "101000";
					when "01010100010011111" => rgb <= "101000";
					when "01010100010100000" => rgb <= "101000";
					when "01010100010100001" => rgb <= "101000";
					when "01010100010100010" => rgb <= "101000";
					when "01010100010100011" => rgb <= "101000";
					when "01010100010100100" => rgb <= "101000";
					when "01010100010100101" => rgb <= "101000";
					when "01010100010100110" => rgb <= "101000";
					when "01010100010100111" => rgb <= "101000";
					when "01010100010101000" => rgb <= "101000";
					when "01010100010101001" => rgb <= "101000";
					when "01010100010101010" => rgb <= "101000";
					when "01010100010101011" => rgb <= "101000";
					when "01010100010101100" => rgb <= "101000";
					when "01010100010101101" => rgb <= "101000";
					when "01010100010101110" => rgb <= "101000";
					when "01010100010101111" => rgb <= "101000";
					when "01010100010110000" => rgb <= "101000";
					when "01010100010110001" => rgb <= "101000";
					when "01010100010110010" => rgb <= "101000";
					when "01010100010110011" => rgb <= "101000";
					when "01010100010110100" => rgb <= "101000";
					when "01010100010110101" => rgb <= "010100";
					when "01010100010110110" => rgb <= "000000";
					when "01010100010110111" => rgb <= "000000";
					when "01010100010111000" => rgb <= "000000";
					when "01010100010111001" => rgb <= "000000";
					when "01010100010111010" => rgb <= "000000";
					when "01010100010111011" => rgb <= "000000";
					when "01010100010111100" => rgb <= "000000";
					when "01010100010111101" => rgb <= "000000";
					when "01010100010111110" => rgb <= "000000";
					when "01010100010111111" => rgb <= "000000";
					when "01010100011000000" => rgb <= "000000";
					when "01010100011000001" => rgb <= "000000";
					when "01010100011000010" => rgb <= "000000";
					when "01010100011000011" => rgb <= "000000";
					when "01010100011000100" => rgb <= "000000";
					when "01010100011000101" => rgb <= "000000";
					when "01010100011000110" => rgb <= "000000";
					when "01010100011000111" => rgb <= "000000";
					when "01010100011001000" => rgb <= "000000";
					when "01010100011001001" => rgb <= "000000";
					when "01010100011001010" => rgb <= "000000";
					when "01010100011001011" => rgb <= "000000";
					when "01010100011001100" => rgb <= "000000";
					when "01010100011001101" => rgb <= "000000";
					when "01010100011001110" => rgb <= "000000";
					when "01010100011001111" => rgb <= "000000";
					when "01010100011010000" => rgb <= "000000";
					when "01010100011010001" => rgb <= "000000";
					when "01010100011010010" => rgb <= "000000";
					when "01010100011010011" => rgb <= "000000";
					when "01010100011010100" => rgb <= "000000";
					when "01010100011010101" => rgb <= "000000";
					when "01010100011010110" => rgb <= "000000";
					when "01010100011010111" => rgb <= "000000";
					when "01010100011011000" => rgb <= "000000";
					when "01010100011011001" => rgb <= "000000";
					when "01010100011011010" => rgb <= "000000";
					when "01010100011011011" => rgb <= "000000";
					when "01010100011011100" => rgb <= "000000";
					when "01010100011011101" => rgb <= "000000";
					when "01010100011011110" => rgb <= "000000";
					when "01010100011011111" => rgb <= "000000";
					when "01010100011100000" => rgb <= "000000";
					when "01010100011100001" => rgb <= "000000";
					when "01010100011100010" => rgb <= "000000";
					when "01010100011100011" => rgb <= "000000";
					when "01010100011100100" => rgb <= "000000";
					when "01010100011100101" => rgb <= "000000";
					when "01010100011100110" => rgb <= "000000";
					when "01010100011100111" => rgb <= "000000";
					when "01010100011101000" => rgb <= "000000";
					when "01010100011101001" => rgb <= "000000";
					when "01010100011101010" => rgb <= "000000";
					when "01010100011101011" => rgb <= "000000";
					when "01010100011101100" => rgb <= "000000";
					when "01010100011101101" => rgb <= "000000";
					when "01010100011101110" => rgb <= "000000";
					when "01010100011101111" => rgb <= "000000";
					when "01010100011110000" => rgb <= "000000";
					when "01010100011110001" => rgb <= "000000";
					when "01010100011110010" => rgb <= "000000";
					when "01010100011110011" => rgb <= "000000";
					when "01010100011110100" => rgb <= "000000";
					when "01010100011110101" => rgb <= "000000";
					when "01010100011110110" => rgb <= "000000";
					when "01010100011110111" => rgb <= "000000";
					when "01010100011111000" => rgb <= "000000";
					when "01010100011111001" => rgb <= "000000";
					when "01010100011111010" => rgb <= "000000";
					when "01010100011111011" => rgb <= "000000";
					when "01010100011111100" => rgb <= "000000";
					when "01010100011111101" => rgb <= "000000";
					when "01010100011111110" => rgb <= "000000";
					when "01010100011111111" => rgb <= "000000";
					when "01010100100000000" => rgb <= "000000";
					when "01010100100000001" => rgb <= "000000";
					when "01010100100000010" => rgb <= "000000";
					when "01010100100000011" => rgb <= "000000";
					when "01010100100000100" => rgb <= "000000";
					when "01010100100000101" => rgb <= "000000";
					when "01010100100000110" => rgb <= "000000";
					when "01010100100000111" => rgb <= "000000";
					when "01010100100001000" => rgb <= "000000";
					when "01010100100001001" => rgb <= "000000";
					when "01010100100001010" => rgb <= "000000";
					when "01010100100001011" => rgb <= "000000";
					when "01010100100001100" => rgb <= "000000";
					when "01010100100001101" => rgb <= "000000";
					when "01010100100001110" => rgb <= "000000";
					when "01010100100001111" => rgb <= "000000";
					when "01010100100010000" => rgb <= "000000";
					when "01010100100010001" => rgb <= "000000";
					when "01010100100010010" => rgb <= "000000";
					when "01010100100010011" => rgb <= "000000";
					when "01010100100010100" => rgb <= "000000";
					when "01010100100010101" => rgb <= "000000";
					when "01010100100010110" => rgb <= "000000";
					when "01010100100010111" => rgb <= "000000";
					when "01010100100011000" => rgb <= "000000";
					when "01010100100011001" => rgb <= "000000";
					when "01010100100011010" => rgb <= "000000";
					when "01010100100011011" => rgb <= "000000";
					when "01010100100011100" => rgb <= "000000";
					when "01010100100011101" => rgb <= "000000";
					when "01010100100011110" => rgb <= "000000";
					when "01010100100011111" => rgb <= "000000";
					when "01010100100100000" => rgb <= "000000";
					when "01010100100100001" => rgb <= "000000";
					when "01010100100100010" => rgb <= "000000";
					when "01010100100100011" => rgb <= "000000";
					when "01010100100100100" => rgb <= "000000";
					when "01010100100100101" => rgb <= "000000";
					when "01010100100100110" => rgb <= "000000";
					when "01010100100100111" => rgb <= "000000";
					when "01010100100101000" => rgb <= "000000";
					when "01010100100101001" => rgb <= "000000";
					when "01010100100101010" => rgb <= "000000";
					when "01010100100101011" => rgb <= "000000";
					when "01010100100101100" => rgb <= "000000";
					when "01010100100101101" => rgb <= "000000";
					when "01010100100101110" => rgb <= "000000";
					when "01010100100101111" => rgb <= "000000";
					when "01010100100110000" => rgb <= "000000";
					when "01010100100110001" => rgb <= "000000";
					when "01010100100110010" => rgb <= "000000";
					when "01010100100110011" => rgb <= "000000";
					when "01010100100110100" => rgb <= "000000";
					when "01010100100110101" => rgb <= "000000";
					when "01010100100110110" => rgb <= "000000";
					when "01010100100110111" => rgb <= "000000";
					when "01010100100111000" => rgb <= "000000";
					when "01010100100111001" => rgb <= "000000";
					when "01010100100111010" => rgb <= "000000";
					when "01010100100111011" => rgb <= "000000";
					when "01010100100111100" => rgb <= "000000";
					when "01010100100111101" => rgb <= "000000";
					when "01010100100111110" => rgb <= "000000";
					when "01010100100111111" => rgb <= "000000";
					when "01010101000000000" => rgb <= "000000";
					when "01010101000000001" => rgb <= "000000";
					when "01010101000000010" => rgb <= "000000";
					when "01010101000000011" => rgb <= "000000";
					when "01010101000000100" => rgb <= "000000";
					when "01010101000000101" => rgb <= "000000";
					when "01010101000000110" => rgb <= "000000";
					when "01010101000000111" => rgb <= "000000";
					when "01010101000001000" => rgb <= "000000";
					when "01010101000001001" => rgb <= "000000";
					when "01010101000001010" => rgb <= "000000";
					when "01010101000001011" => rgb <= "000000";
					when "01010101000001100" => rgb <= "000000";
					when "01010101000001101" => rgb <= "000000";
					when "01010101000001110" => rgb <= "000000";
					when "01010101000001111" => rgb <= "000000";
					when "01010101000010000" => rgb <= "000000";
					when "01010101000010001" => rgb <= "000000";
					when "01010101000010010" => rgb <= "000000";
					when "01010101000010011" => rgb <= "000000";
					when "01010101000010100" => rgb <= "000000";
					when "01010101000010101" => rgb <= "000000";
					when "01010101000010110" => rgb <= "000000";
					when "01010101000010111" => rgb <= "000000";
					when "01010101000011000" => rgb <= "000000";
					when "01010101000011001" => rgb <= "000000";
					when "01010101000011010" => rgb <= "000000";
					when "01010101000011011" => rgb <= "000000";
					when "01010101000011100" => rgb <= "000000";
					when "01010101000011101" => rgb <= "000000";
					when "01010101000011110" => rgb <= "000000";
					when "01010101000011111" => rgb <= "000000";
					when "01010101000100000" => rgb <= "000000";
					when "01010101000100001" => rgb <= "000000";
					when "01010101000100010" => rgb <= "000000";
					when "01010101000100011" => rgb <= "000000";
					when "01010101000100100" => rgb <= "000000";
					when "01010101000100101" => rgb <= "000000";
					when "01010101000100110" => rgb <= "000000";
					when "01010101000100111" => rgb <= "000000";
					when "01010101000101000" => rgb <= "000000";
					when "01010101000101001" => rgb <= "000000";
					when "01010101000101010" => rgb <= "000000";
					when "01010101000101011" => rgb <= "000000";
					when "01010101000101100" => rgb <= "000000";
					when "01010101000101101" => rgb <= "000000";
					when "01010101000101110" => rgb <= "000000";
					when "01010101000101111" => rgb <= "000000";
					when "01010101000110000" => rgb <= "000000";
					when "01010101000110001" => rgb <= "000000";
					when "01010101000110010" => rgb <= "000000";
					when "01010101000110011" => rgb <= "000000";
					when "01010101000110100" => rgb <= "000000";
					when "01010101000110101" => rgb <= "000000";
					when "01010101000110110" => rgb <= "000000";
					when "01010101000110111" => rgb <= "000000";
					when "01010101000111000" => rgb <= "000000";
					when "01010101000111001" => rgb <= "000000";
					when "01010101000111010" => rgb <= "000000";
					when "01010101000111011" => rgb <= "000000";
					when "01010101000111100" => rgb <= "000000";
					when "01010101000111101" => rgb <= "000000";
					when "01010101000111110" => rgb <= "000000";
					when "01010101000111111" => rgb <= "000000";
					when "01010101001000000" => rgb <= "000000";
					when "01010101001000001" => rgb <= "000000";
					when "01010101001000010" => rgb <= "000000";
					when "01010101001000011" => rgb <= "000000";
					when "01010101001000100" => rgb <= "000000";
					when "01010101001000101" => rgb <= "000000";
					when "01010101001000110" => rgb <= "000000";
					when "01010101001000111" => rgb <= "000000";
					when "01010101001001000" => rgb <= "000000";
					when "01010101001001001" => rgb <= "000000";
					when "01010101001001010" => rgb <= "000000";
					when "01010101001001011" => rgb <= "000000";
					when "01010101001001100" => rgb <= "000000";
					when "01010101001001101" => rgb <= "000000";
					when "01010101001001110" => rgb <= "000000";
					when "01010101001001111" => rgb <= "000000";
					when "01010101001010000" => rgb <= "000000";
					when "01010101001010001" => rgb <= "000000";
					when "01010101001010010" => rgb <= "000000";
					when "01010101001010011" => rgb <= "000000";
					when "01010101001010100" => rgb <= "000000";
					when "01010101001010101" => rgb <= "000000";
					when "01010101001010110" => rgb <= "000000";
					when "01010101001010111" => rgb <= "000000";
					when "01010101001011000" => rgb <= "000000";
					when "01010101001011001" => rgb <= "000000";
					when "01010101001011010" => rgb <= "000000";
					when "01010101001011011" => rgb <= "000000";
					when "01010101001011100" => rgb <= "000000";
					when "01010101001011101" => rgb <= "000000";
					when "01010101001011110" => rgb <= "000000";
					when "01010101001011111" => rgb <= "000000";
					when "01010101001100000" => rgb <= "000000";
					when "01010101001100001" => rgb <= "000000";
					when "01010101001100010" => rgb <= "000000";
					when "01010101001100011" => rgb <= "000000";
					when "01010101001100100" => rgb <= "000000";
					when "01010101001100101" => rgb <= "000000";
					when "01010101001100110" => rgb <= "000000";
					when "01010101001100111" => rgb <= "000000";
					when "01010101001101000" => rgb <= "000000";
					when "01010101001101001" => rgb <= "000000";
					when "01010101001101010" => rgb <= "000000";
					when "01010101001101011" => rgb <= "000000";
					when "01010101001101100" => rgb <= "000000";
					when "01010101001101101" => rgb <= "000000";
					when "01010101001101110" => rgb <= "000000";
					when "01010101001101111" => rgb <= "000000";
					when "01010101001110000" => rgb <= "000000";
					when "01010101001110001" => rgb <= "000000";
					when "01010101001110010" => rgb <= "000000";
					when "01010101001110011" => rgb <= "000000";
					when "01010101001110100" => rgb <= "000000";
					when "01010101001110101" => rgb <= "000000";
					when "01010101001110110" => rgb <= "000000";
					when "01010101001110111" => rgb <= "000000";
					when "01010101001111000" => rgb <= "000000";
					when "01010101001111001" => rgb <= "000000";
					when "01010101001111010" => rgb <= "000000";
					when "01010101001111011" => rgb <= "000000";
					when "01010101001111100" => rgb <= "000000";
					when "01010101001111101" => rgb <= "000000";
					when "01010101001111110" => rgb <= "000000";
					when "01010101001111111" => rgb <= "000000";
					when "01010101010000000" => rgb <= "000000";
					when "01010101010000001" => rgb <= "000000";
					when "01010101010000010" => rgb <= "000000";
					when "01010101010000011" => rgb <= "000000";
					when "01010101010000100" => rgb <= "000000";
					when "01010101010000101" => rgb <= "000000";
					when "01010101010000110" => rgb <= "000000";
					when "01010101010000111" => rgb <= "000000";
					when "01010101010001000" => rgb <= "000000";
					when "01010101010001001" => rgb <= "000000";
					when "01010101010001010" => rgb <= "000000";
					when "01010101010001011" => rgb <= "000000";
					when "01010101010001100" => rgb <= "000000";
					when "01010101010001101" => rgb <= "000000";
					when "01010101010001110" => rgb <= "000000";
					when "01010101010001111" => rgb <= "000000";
					when "01010101010010000" => rgb <= "000000";
					when "01010101010010001" => rgb <= "000000";
					when "01010101010010010" => rgb <= "000000";
					when "01010101010010011" => rgb <= "010100";
					when "01010101010010100" => rgb <= "101000";
					when "01010101010010101" => rgb <= "101000";
					when "01010101010010110" => rgb <= "101000";
					when "01010101010010111" => rgb <= "101000";
					when "01010101010011000" => rgb <= "101000";
					when "01010101010011001" => rgb <= "101000";
					when "01010101010011010" => rgb <= "101000";
					when "01010101010011011" => rgb <= "101000";
					when "01010101010011100" => rgb <= "101000";
					when "01010101010011101" => rgb <= "101000";
					when "01010101010011110" => rgb <= "101000";
					when "01010101010011111" => rgb <= "101000";
					when "01010101010100000" => rgb <= "101000";
					when "01010101010100001" => rgb <= "101000";
					when "01010101010100010" => rgb <= "101000";
					when "01010101010100011" => rgb <= "101000";
					when "01010101010100100" => rgb <= "101000";
					when "01010101010100101" => rgb <= "101000";
					when "01010101010100110" => rgb <= "101000";
					when "01010101010100111" => rgb <= "101000";
					when "01010101010101000" => rgb <= "101000";
					when "01010101010101001" => rgb <= "101000";
					when "01010101010101010" => rgb <= "010100";
					when "01010101010101011" => rgb <= "000000";
					when "01010101010101100" => rgb <= "000000";
					when "01010101010101101" => rgb <= "000000";
					when "01010101010101110" => rgb <= "000000";
					when "01010101010101111" => rgb <= "000000";
					when "01010101010110000" => rgb <= "000000";
					when "01010101010110001" => rgb <= "000000";
					when "01010101010110010" => rgb <= "000000";
					when "01010101010110011" => rgb <= "000000";
					when "01010101010110100" => rgb <= "000000";
					when "01010101010110101" => rgb <= "000000";
					when "01010101010110110" => rgb <= "000000";
					when "01010101010110111" => rgb <= "000000";
					when "01010101010111000" => rgb <= "000000";
					when "01010101010111001" => rgb <= "000000";
					when "01010101010111010" => rgb <= "000000";
					when "01010101010111011" => rgb <= "000000";
					when "01010101010111100" => rgb <= "000000";
					when "01010101010111101" => rgb <= "000000";
					when "01010101010111110" => rgb <= "000000";
					when "01010101010111111" => rgb <= "000000";
					when "01010101011000000" => rgb <= "000000";
					when "01010101011000001" => rgb <= "000000";
					when "01010101011000010" => rgb <= "000000";
					when "01010101011000011" => rgb <= "000000";
					when "01010101011000100" => rgb <= "000000";
					when "01010101011000101" => rgb <= "000000";
					when "01010101011000110" => rgb <= "000000";
					when "01010101011000111" => rgb <= "000000";
					when "01010101011001000" => rgb <= "000000";
					when "01010101011001001" => rgb <= "000000";
					when "01010101011001010" => rgb <= "000000";
					when "01010101011001011" => rgb <= "000000";
					when "01010101011001100" => rgb <= "000000";
					when "01010101011001101" => rgb <= "000000";
					when "01010101011001110" => rgb <= "000000";
					when "01010101011001111" => rgb <= "000000";
					when "01010101011010000" => rgb <= "000000";
					when "01010101011010001" => rgb <= "000000";
					when "01010101011010010" => rgb <= "000000";
					when "01010101011010011" => rgb <= "000000";
					when "01010101011010100" => rgb <= "000000";
					when "01010101011010101" => rgb <= "000000";
					when "01010101011010110" => rgb <= "000000";
					when "01010101011010111" => rgb <= "000000";
					when "01010101011011000" => rgb <= "000000";
					when "01010101011011001" => rgb <= "000000";
					when "01010101011011010" => rgb <= "000000";
					when "01010101011011011" => rgb <= "000000";
					when "01010101011011100" => rgb <= "000000";
					when "01010101011011101" => rgb <= "000000";
					when "01010101011011110" => rgb <= "000000";
					when "01010101011011111" => rgb <= "000000";
					when "01010101011100000" => rgb <= "000000";
					when "01010101011100001" => rgb <= "000000";
					when "01010101011100010" => rgb <= "000000";
					when "01010101011100011" => rgb <= "000000";
					when "01010101011100100" => rgb <= "000000";
					when "01010101011100101" => rgb <= "000000";
					when "01010101011100110" => rgb <= "000000";
					when "01010101011100111" => rgb <= "000000";
					when "01010101011101000" => rgb <= "000000";
					when "01010101011101001" => rgb <= "000000";
					when "01010101011101010" => rgb <= "000000";
					when "01010101011101011" => rgb <= "000000";
					when "01010101011101100" => rgb <= "000000";
					when "01010101011101101" => rgb <= "000000";
					when "01010101011101110" => rgb <= "000000";
					when "01010101011101111" => rgb <= "000000";
					when "01010101011110000" => rgb <= "000000";
					when "01010101011110001" => rgb <= "000000";
					when "01010101011110010" => rgb <= "000000";
					when "01010101011110011" => rgb <= "000000";
					when "01010101011110100" => rgb <= "000000";
					when "01010101011110101" => rgb <= "000000";
					when "01010101011110110" => rgb <= "000000";
					when "01010101011110111" => rgb <= "000000";
					when "01010101011111000" => rgb <= "000000";
					when "01010101011111001" => rgb <= "000000";
					when "01010101011111010" => rgb <= "000000";
					when "01010101011111011" => rgb <= "000000";
					when "01010101011111100" => rgb <= "000000";
					when "01010101011111101" => rgb <= "000000";
					when "01010101011111110" => rgb <= "000000";
					when "01010101011111111" => rgb <= "000000";
					when "01010101100000000" => rgb <= "000000";
					when "01010101100000001" => rgb <= "000000";
					when "01010101100000010" => rgb <= "000000";
					when "01010101100000011" => rgb <= "000000";
					when "01010101100000100" => rgb <= "000000";
					when "01010101100000101" => rgb <= "000000";
					when "01010101100000110" => rgb <= "000000";
					when "01010101100000111" => rgb <= "000000";
					when "01010101100001000" => rgb <= "000000";
					when "01010101100001001" => rgb <= "000000";
					when "01010101100001010" => rgb <= "000000";
					when "01010101100001011" => rgb <= "000000";
					when "01010101100001100" => rgb <= "000000";
					when "01010101100001101" => rgb <= "000000";
					when "01010101100001110" => rgb <= "000000";
					when "01010101100001111" => rgb <= "000000";
					when "01010101100010000" => rgb <= "000000";
					when "01010101100010001" => rgb <= "000000";
					when "01010101100010010" => rgb <= "000000";
					when "01010101100010011" => rgb <= "000000";
					when "01010101100010100" => rgb <= "000000";
					when "01010101100010101" => rgb <= "000000";
					when "01010101100010110" => rgb <= "000000";
					when "01010101100010111" => rgb <= "000000";
					when "01010101100011000" => rgb <= "000000";
					when "01010101100011001" => rgb <= "000000";
					when "01010101100011010" => rgb <= "000000";
					when "01010101100011011" => rgb <= "000000";
					when "01010101100011100" => rgb <= "000000";
					when "01010101100011101" => rgb <= "000000";
					when "01010101100011110" => rgb <= "000000";
					when "01010101100011111" => rgb <= "000000";
					when "01010101100100000" => rgb <= "000000";
					when "01010101100100001" => rgb <= "000000";
					when "01010101100100010" => rgb <= "000000";
					when "01010101100100011" => rgb <= "000000";
					when "01010101100100100" => rgb <= "000000";
					when "01010101100100101" => rgb <= "000000";
					when "01010101100100110" => rgb <= "000000";
					when "01010101100100111" => rgb <= "000000";
					when "01010101100101000" => rgb <= "000000";
					when "01010101100101001" => rgb <= "000000";
					when "01010101100101010" => rgb <= "000000";
					when "01010101100101011" => rgb <= "000000";
					when "01010101100101100" => rgb <= "000000";
					when "01010101100101101" => rgb <= "000000";
					when "01010101100101110" => rgb <= "000000";
					when "01010101100101111" => rgb <= "000000";
					when "01010101100110000" => rgb <= "000000";
					when "01010101100110001" => rgb <= "000000";
					when "01010101100110010" => rgb <= "000000";
					when "01010101100110011" => rgb <= "000000";
					when "01010101100110100" => rgb <= "000000";
					when "01010101100110101" => rgb <= "000000";
					when "01010101100110110" => rgb <= "000000";
					when "01010101100110111" => rgb <= "000000";
					when "01010101100111000" => rgb <= "000000";
					when "01010101100111001" => rgb <= "000000";
					when "01010101100111010" => rgb <= "000000";
					when "01010101100111011" => rgb <= "000000";
					when "01010101100111100" => rgb <= "000000";
					when "01010101100111101" => rgb <= "000000";
					when "01010101100111110" => rgb <= "000000";
					when "01010101100111111" => rgb <= "000000";
					when "01010110000000000" => rgb <= "000000";
					when "01010110000000001" => rgb <= "000000";
					when "01010110000000010" => rgb <= "000000";
					when "01010110000000011" => rgb <= "000000";
					when "01010110000000100" => rgb <= "000000";
					when "01010110000000101" => rgb <= "000000";
					when "01010110000000110" => rgb <= "000000";
					when "01010110000000111" => rgb <= "000000";
					when "01010110000001000" => rgb <= "000000";
					when "01010110000001001" => rgb <= "000000";
					when "01010110000001010" => rgb <= "000000";
					when "01010110000001011" => rgb <= "000000";
					when "01010110000001100" => rgb <= "000000";
					when "01010110000001101" => rgb <= "000000";
					when "01010110000001110" => rgb <= "000000";
					when "01010110000001111" => rgb <= "000000";
					when "01010110000010000" => rgb <= "000000";
					when "01010110000010001" => rgb <= "000000";
					when "01010110000010010" => rgb <= "000000";
					when "01010110000010011" => rgb <= "000000";
					when "01010110000010100" => rgb <= "000000";
					when "01010110000010101" => rgb <= "000000";
					when "01010110000010110" => rgb <= "000000";
					when "01010110000010111" => rgb <= "000000";
					when "01010110000011000" => rgb <= "000000";
					when "01010110000011001" => rgb <= "000000";
					when "01010110000011010" => rgb <= "000000";
					when "01010110000011011" => rgb <= "000000";
					when "01010110000011100" => rgb <= "000000";
					when "01010110000011101" => rgb <= "000000";
					when "01010110000011110" => rgb <= "000000";
					when "01010110000011111" => rgb <= "000000";
					when "01010110000100000" => rgb <= "000000";
					when "01010110000100001" => rgb <= "000000";
					when "01010110000100010" => rgb <= "000000";
					when "01010110000100011" => rgb <= "000000";
					when "01010110000100100" => rgb <= "000000";
					when "01010110000100101" => rgb <= "000000";
					when "01010110000100110" => rgb <= "000000";
					when "01010110000100111" => rgb <= "000000";
					when "01010110000101000" => rgb <= "000000";
					when "01010110000101001" => rgb <= "000000";
					when "01010110000101010" => rgb <= "000000";
					when "01010110000101011" => rgb <= "000000";
					when "01010110000101100" => rgb <= "000000";
					when "01010110000101101" => rgb <= "000000";
					when "01010110000101110" => rgb <= "000000";
					when "01010110000101111" => rgb <= "000000";
					when "01010110000110000" => rgb <= "000000";
					when "01010110000110001" => rgb <= "000000";
					when "01010110000110010" => rgb <= "000000";
					when "01010110000110011" => rgb <= "000000";
					when "01010110000110100" => rgb <= "000000";
					when "01010110000110101" => rgb <= "000000";
					when "01010110000110110" => rgb <= "000000";
					when "01010110000110111" => rgb <= "000000";
					when "01010110000111000" => rgb <= "000000";
					when "01010110000111001" => rgb <= "000000";
					when "01010110000111010" => rgb <= "000000";
					when "01010110000111011" => rgb <= "000000";
					when "01010110000111100" => rgb <= "000000";
					when "01010110000111101" => rgb <= "000000";
					when "01010110000111110" => rgb <= "000000";
					when "01010110000111111" => rgb <= "000000";
					when "01010110001000000" => rgb <= "000000";
					when "01010110001000001" => rgb <= "000000";
					when "01010110001000010" => rgb <= "000000";
					when "01010110001000011" => rgb <= "000000";
					when "01010110001000100" => rgb <= "000000";
					when "01010110001000101" => rgb <= "000000";
					when "01010110001000110" => rgb <= "000000";
					when "01010110001000111" => rgb <= "000000";
					when "01010110001001000" => rgb <= "000000";
					when "01010110001001001" => rgb <= "000000";
					when "01010110001001010" => rgb <= "000000";
					when "01010110001001011" => rgb <= "000000";
					when "01010110001001100" => rgb <= "000000";
					when "01010110001001101" => rgb <= "000000";
					when "01010110001001110" => rgb <= "000000";
					when "01010110001001111" => rgb <= "000000";
					when "01010110001010000" => rgb <= "000000";
					when "01010110001010001" => rgb <= "000000";
					when "01010110001010010" => rgb <= "000000";
					when "01010110001010011" => rgb <= "000000";
					when "01010110001010100" => rgb <= "000000";
					when "01010110001010101" => rgb <= "000000";
					when "01010110001010110" => rgb <= "000000";
					when "01010110001010111" => rgb <= "000000";
					when "01010110001011000" => rgb <= "000000";
					when "01010110001011001" => rgb <= "000000";
					when "01010110001011010" => rgb <= "000000";
					when "01010110001011011" => rgb <= "000000";
					when "01010110001011100" => rgb <= "000000";
					when "01010110001011101" => rgb <= "000000";
					when "01010110001011110" => rgb <= "000000";
					when "01010110001011111" => rgb <= "000000";
					when "01010110001100000" => rgb <= "000000";
					when "01010110001100001" => rgb <= "000000";
					when "01010110001100010" => rgb <= "000000";
					when "01010110001100011" => rgb <= "000000";
					when "01010110001100100" => rgb <= "000000";
					when "01010110001100101" => rgb <= "000000";
					when "01010110001100110" => rgb <= "000000";
					when "01010110001100111" => rgb <= "000000";
					when "01010110001101000" => rgb <= "000000";
					when "01010110001101001" => rgb <= "000000";
					when "01010110001101010" => rgb <= "000000";
					when "01010110001101011" => rgb <= "000000";
					when "01010110001101100" => rgb <= "000000";
					when "01010110001101101" => rgb <= "000000";
					when "01010110001101110" => rgb <= "000000";
					when "01010110001101111" => rgb <= "000000";
					when "01010110001110000" => rgb <= "000000";
					when "01010110001110001" => rgb <= "000000";
					when "01010110001110010" => rgb <= "000000";
					when "01010110001110011" => rgb <= "000000";
					when "01010110001110100" => rgb <= "000000";
					when "01010110001110101" => rgb <= "000000";
					when "01010110001110110" => rgb <= "000000";
					when "01010110001110111" => rgb <= "000000";
					when "01010110001111000" => rgb <= "000000";
					when "01010110001111001" => rgb <= "000000";
					when "01010110001111010" => rgb <= "000000";
					when "01010110001111011" => rgb <= "000000";
					when "01010110001111100" => rgb <= "000000";
					when "01010110001111101" => rgb <= "000000";
					when "01010110001111110" => rgb <= "000000";
					when "01010110001111111" => rgb <= "000000";
					when "01010110010000000" => rgb <= "000000";
					when "01010110010000001" => rgb <= "000000";
					when "01010110010000010" => rgb <= "000000";
					when "01010110010000011" => rgb <= "000000";
					when "01010110010000100" => rgb <= "000000";
					when "01010110010000101" => rgb <= "000000";
					when "01010110010000110" => rgb <= "000000";
					when "01010110010000111" => rgb <= "000000";
					when "01010110010001000" => rgb <= "000000";
					when "01010110010001001" => rgb <= "000000";
					when "01010110010001010" => rgb <= "000000";
					when "01010110010001011" => rgb <= "000000";
					when "01010110010001100" => rgb <= "000000";
					when "01010110010001101" => rgb <= "000000";
					when "01010110010001110" => rgb <= "000000";
					when "01010110010001111" => rgb <= "000000";
					when "01010110010010000" => rgb <= "000000";
					when "01010110010010001" => rgb <= "000000";
					when "01010110010010010" => rgb <= "000000";
					when "01010110010010011" => rgb <= "010000";
					when "01010110010010100" => rgb <= "101000";
					when "01010110010010101" => rgb <= "101000";
					when "01010110010010110" => rgb <= "101000";
					when "01010110010010111" => rgb <= "101000";
					when "01010110010011000" => rgb <= "101000";
					when "01010110010011001" => rgb <= "101000";
					when "01010110010011010" => rgb <= "101000";
					when "01010110010011011" => rgb <= "101000";
					when "01010110010011100" => rgb <= "101000";
					when "01010110010011101" => rgb <= "101000";
					when "01010110010011110" => rgb <= "101000";
					when "01010110010011111" => rgb <= "101000";
					when "01010110010100000" => rgb <= "101000";
					when "01010110010100001" => rgb <= "101000";
					when "01010110010100010" => rgb <= "101000";
					when "01010110010100011" => rgb <= "101000";
					when "01010110010100100" => rgb <= "101000";
					when "01010110010100101" => rgb <= "101000";
					when "01010110010100110" => rgb <= "101000";
					when "01010110010100111" => rgb <= "101000";
					when "01010110010101000" => rgb <= "101000";
					when "01010110010101001" => rgb <= "101000";
					when "01010110010101010" => rgb <= "000000";
					when "01010110010101011" => rgb <= "000000";
					when "01010110010101100" => rgb <= "000000";
					when "01010110010101101" => rgb <= "000000";
					when "01010110010101110" => rgb <= "000000";
					when "01010110010101111" => rgb <= "000000";
					when "01010110010110000" => rgb <= "000000";
					when "01010110010110001" => rgb <= "000000";
					when "01010110010110010" => rgb <= "000000";
					when "01010110010110011" => rgb <= "000000";
					when "01010110010110100" => rgb <= "000000";
					when "01010110010110101" => rgb <= "000000";
					when "01010110010110110" => rgb <= "000000";
					when "01010110010110111" => rgb <= "000000";
					when "01010110010111000" => rgb <= "000000";
					when "01010110010111001" => rgb <= "000000";
					when "01010110010111010" => rgb <= "000000";
					when "01010110010111011" => rgb <= "000000";
					when "01010110010111100" => rgb <= "000000";
					when "01010110010111101" => rgb <= "000000";
					when "01010110010111110" => rgb <= "000000";
					when "01010110010111111" => rgb <= "000000";
					when "01010110011000000" => rgb <= "000000";
					when "01010110011000001" => rgb <= "000000";
					when "01010110011000010" => rgb <= "000000";
					when "01010110011000011" => rgb <= "000000";
					when "01010110011000100" => rgb <= "000000";
					when "01010110011000101" => rgb <= "000000";
					when "01010110011000110" => rgb <= "000000";
					when "01010110011000111" => rgb <= "000000";
					when "01010110011001000" => rgb <= "000000";
					when "01010110011001001" => rgb <= "000000";
					when "01010110011001010" => rgb <= "000000";
					when "01010110011001011" => rgb <= "000000";
					when "01010110011001100" => rgb <= "000000";
					when "01010110011001101" => rgb <= "000000";
					when "01010110011001110" => rgb <= "000000";
					when "01010110011001111" => rgb <= "000000";
					when "01010110011010000" => rgb <= "000000";
					when "01010110011010001" => rgb <= "000000";
					when "01010110011010010" => rgb <= "000000";
					when "01010110011010011" => rgb <= "000000";
					when "01010110011010100" => rgb <= "000000";
					when "01010110011010101" => rgb <= "000000";
					when "01010110011010110" => rgb <= "000000";
					when "01010110011010111" => rgb <= "000000";
					when "01010110011011000" => rgb <= "000000";
					when "01010110011011001" => rgb <= "000000";
					when "01010110011011010" => rgb <= "000000";
					when "01010110011011011" => rgb <= "000000";
					when "01010110011011100" => rgb <= "000000";
					when "01010110011011101" => rgb <= "000000";
					when "01010110011011110" => rgb <= "000000";
					when "01010110011011111" => rgb <= "000000";
					when "01010110011100000" => rgb <= "000000";
					when "01010110011100001" => rgb <= "000000";
					when "01010110011100010" => rgb <= "000000";
					when "01010110011100011" => rgb <= "000000";
					when "01010110011100100" => rgb <= "000000";
					when "01010110011100101" => rgb <= "000000";
					when "01010110011100110" => rgb <= "000000";
					when "01010110011100111" => rgb <= "000000";
					when "01010110011101000" => rgb <= "000000";
					when "01010110011101001" => rgb <= "000000";
					when "01010110011101010" => rgb <= "000000";
					when "01010110011101011" => rgb <= "000000";
					when "01010110011101100" => rgb <= "000000";
					when "01010110011101101" => rgb <= "000000";
					when "01010110011101110" => rgb <= "000000";
					when "01010110011101111" => rgb <= "000000";
					when "01010110011110000" => rgb <= "000000";
					when "01010110011110001" => rgb <= "000000";
					when "01010110011110010" => rgb <= "000000";
					when "01010110011110011" => rgb <= "000000";
					when "01010110011110100" => rgb <= "000000";
					when "01010110011110101" => rgb <= "000000";
					when "01010110011110110" => rgb <= "000000";
					when "01010110011110111" => rgb <= "000000";
					when "01010110011111000" => rgb <= "000000";
					when "01010110011111001" => rgb <= "000000";
					when "01010110011111010" => rgb <= "000000";
					when "01010110011111011" => rgb <= "000000";
					when "01010110011111100" => rgb <= "000000";
					when "01010110011111101" => rgb <= "000000";
					when "01010110011111110" => rgb <= "000000";
					when "01010110011111111" => rgb <= "000000";
					when "01010110100000000" => rgb <= "000000";
					when "01010110100000001" => rgb <= "000000";
					when "01010110100000010" => rgb <= "000000";
					when "01010110100000011" => rgb <= "000000";
					when "01010110100000100" => rgb <= "000000";
					when "01010110100000101" => rgb <= "000000";
					when "01010110100000110" => rgb <= "000000";
					when "01010110100000111" => rgb <= "000000";
					when "01010110100001000" => rgb <= "000000";
					when "01010110100001001" => rgb <= "000000";
					when "01010110100001010" => rgb <= "000000";
					when "01010110100001011" => rgb <= "000000";
					when "01010110100001100" => rgb <= "000000";
					when "01010110100001101" => rgb <= "000000";
					when "01010110100001110" => rgb <= "000000";
					when "01010110100001111" => rgb <= "000000";
					when "01010110100010000" => rgb <= "000000";
					when "01010110100010001" => rgb <= "000000";
					when "01010110100010010" => rgb <= "000000";
					when "01010110100010011" => rgb <= "000000";
					when "01010110100010100" => rgb <= "000000";
					when "01010110100010101" => rgb <= "000000";
					when "01010110100010110" => rgb <= "000000";
					when "01010110100010111" => rgb <= "000000";
					when "01010110100011000" => rgb <= "000000";
					when "01010110100011001" => rgb <= "000000";
					when "01010110100011010" => rgb <= "000000";
					when "01010110100011011" => rgb <= "000000";
					when "01010110100011100" => rgb <= "000000";
					when "01010110100011101" => rgb <= "000000";
					when "01010110100011110" => rgb <= "000000";
					when "01010110100011111" => rgb <= "000000";
					when "01010110100100000" => rgb <= "000000";
					when "01010110100100001" => rgb <= "000000";
					when "01010110100100010" => rgb <= "000000";
					when "01010110100100011" => rgb <= "000000";
					when "01010110100100100" => rgb <= "000000";
					when "01010110100100101" => rgb <= "000000";
					when "01010110100100110" => rgb <= "000000";
					when "01010110100100111" => rgb <= "000000";
					when "01010110100101000" => rgb <= "000000";
					when "01010110100101001" => rgb <= "000000";
					when "01010110100101010" => rgb <= "000000";
					when "01010110100101011" => rgb <= "000000";
					when "01010110100101100" => rgb <= "000000";
					when "01010110100101101" => rgb <= "000000";
					when "01010110100101110" => rgb <= "000000";
					when "01010110100101111" => rgb <= "000000";
					when "01010110100110000" => rgb <= "000000";
					when "01010110100110001" => rgb <= "000000";
					when "01010110100110010" => rgb <= "000000";
					when "01010110100110011" => rgb <= "000000";
					when "01010110100110100" => rgb <= "000000";
					when "01010110100110101" => rgb <= "000000";
					when "01010110100110110" => rgb <= "000000";
					when "01010110100110111" => rgb <= "000000";
					when "01010110100111000" => rgb <= "000000";
					when "01010110100111001" => rgb <= "000000";
					when "01010110100111010" => rgb <= "000000";
					when "01010110100111011" => rgb <= "000000";
					when "01010110100111100" => rgb <= "000000";
					when "01010110100111101" => rgb <= "000000";
					when "01010110100111110" => rgb <= "000000";
					when "01010110100111111" => rgb <= "000000";
					when "01010111000000000" => rgb <= "000000";
					when "01010111000000001" => rgb <= "000000";
					when "01010111000000010" => rgb <= "000000";
					when "01010111000000011" => rgb <= "000000";
					when "01010111000000100" => rgb <= "000000";
					when "01010111000000101" => rgb <= "000000";
					when "01010111000000110" => rgb <= "000000";
					when "01010111000000111" => rgb <= "000000";
					when "01010111000001000" => rgb <= "000000";
					when "01010111000001001" => rgb <= "000000";
					when "01010111000001010" => rgb <= "000000";
					when "01010111000001011" => rgb <= "000000";
					when "01010111000001100" => rgb <= "000000";
					when "01010111000001101" => rgb <= "000000";
					when "01010111000001110" => rgb <= "000000";
					when "01010111000001111" => rgb <= "000000";
					when "01010111000010000" => rgb <= "000000";
					when "01010111000010001" => rgb <= "000000";
					when "01010111000010010" => rgb <= "000000";
					when "01010111000010011" => rgb <= "000000";
					when "01010111000010100" => rgb <= "000000";
					when "01010111000010101" => rgb <= "000000";
					when "01010111000010110" => rgb <= "000000";
					when "01010111000010111" => rgb <= "000000";
					when "01010111000011000" => rgb <= "000000";
					when "01010111000011001" => rgb <= "000000";
					when "01010111000011010" => rgb <= "000000";
					when "01010111000011011" => rgb <= "000000";
					when "01010111000011100" => rgb <= "000000";
					when "01010111000011101" => rgb <= "000000";
					when "01010111000011110" => rgb <= "000000";
					when "01010111000011111" => rgb <= "000000";
					when "01010111000100000" => rgb <= "000000";
					when "01010111000100001" => rgb <= "000000";
					when "01010111000100010" => rgb <= "000000";
					when "01010111000100011" => rgb <= "000000";
					when "01010111000100100" => rgb <= "000000";
					when "01010111000100101" => rgb <= "000000";
					when "01010111000100110" => rgb <= "000000";
					when "01010111000100111" => rgb <= "000000";
					when "01010111000101000" => rgb <= "000000";
					when "01010111000101001" => rgb <= "000000";
					when "01010111000101010" => rgb <= "000000";
					when "01010111000101011" => rgb <= "000000";
					when "01010111000101100" => rgb <= "000000";
					when "01010111000101101" => rgb <= "000000";
					when "01010111000101110" => rgb <= "000000";
					when "01010111000101111" => rgb <= "000000";
					when "01010111000110000" => rgb <= "000000";
					when "01010111000110001" => rgb <= "000000";
					when "01010111000110010" => rgb <= "000000";
					when "01010111000110011" => rgb <= "000000";
					when "01010111000110100" => rgb <= "000000";
					when "01010111000110101" => rgb <= "000000";
					when "01010111000110110" => rgb <= "000000";
					when "01010111000110111" => rgb <= "000000";
					when "01010111000111000" => rgb <= "000000";
					when "01010111000111001" => rgb <= "000000";
					when "01010111000111010" => rgb <= "000000";
					when "01010111000111011" => rgb <= "000000";
					when "01010111000111100" => rgb <= "000000";
					when "01010111000111101" => rgb <= "000000";
					when "01010111000111110" => rgb <= "000000";
					when "01010111000111111" => rgb <= "000000";
					when "01010111001000000" => rgb <= "000000";
					when "01010111001000001" => rgb <= "000000";
					when "01010111001000010" => rgb <= "000000";
					when "01010111001000011" => rgb <= "000000";
					when "01010111001000100" => rgb <= "000000";
					when "01010111001000101" => rgb <= "000000";
					when "01010111001000110" => rgb <= "000000";
					when "01010111001000111" => rgb <= "000000";
					when "01010111001001000" => rgb <= "000000";
					when "01010111001001001" => rgb <= "000000";
					when "01010111001001010" => rgb <= "000000";
					when "01010111001001011" => rgb <= "000000";
					when "01010111001001100" => rgb <= "000000";
					when "01010111001001101" => rgb <= "000000";
					when "01010111001001110" => rgb <= "000000";
					when "01010111001001111" => rgb <= "000000";
					when "01010111001010000" => rgb <= "000000";
					when "01010111001010001" => rgb <= "000000";
					when "01010111001010010" => rgb <= "000000";
					when "01010111001010011" => rgb <= "000000";
					when "01010111001010100" => rgb <= "000000";
					when "01010111001010101" => rgb <= "000000";
					when "01010111001010110" => rgb <= "000000";
					when "01010111001010111" => rgb <= "000000";
					when "01010111001011000" => rgb <= "000000";
					when "01010111001011001" => rgb <= "000000";
					when "01010111001011010" => rgb <= "000000";
					when "01010111001011011" => rgb <= "000000";
					when "01010111001011100" => rgb <= "000000";
					when "01010111001011101" => rgb <= "000000";
					when "01010111001011110" => rgb <= "000000";
					when "01010111001011111" => rgb <= "000000";
					when "01010111001100000" => rgb <= "000000";
					when "01010111001100001" => rgb <= "000000";
					when "01010111001100010" => rgb <= "000000";
					when "01010111001100011" => rgb <= "000000";
					when "01010111001100100" => rgb <= "000000";
					when "01010111001100101" => rgb <= "000000";
					when "01010111001100110" => rgb <= "000000";
					when "01010111001100111" => rgb <= "000000";
					when "01010111001101000" => rgb <= "000000";
					when "01010111001101001" => rgb <= "000000";
					when "01010111001101010" => rgb <= "000000";
					when "01010111001101011" => rgb <= "000000";
					when "01010111001101100" => rgb <= "000000";
					when "01010111001101101" => rgb <= "000000";
					when "01010111001101110" => rgb <= "000000";
					when "01010111001101111" => rgb <= "000000";
					when "01010111001110000" => rgb <= "000000";
					when "01010111001110001" => rgb <= "000000";
					when "01010111001110010" => rgb <= "000000";
					when "01010111001110011" => rgb <= "000000";
					when "01010111001110100" => rgb <= "000000";
					when "01010111001110101" => rgb <= "000000";
					when "01010111001110110" => rgb <= "000000";
					when "01010111001110111" => rgb <= "000000";
					when "01010111001111000" => rgb <= "000000";
					when "01010111001111001" => rgb <= "000000";
					when "01010111001111010" => rgb <= "000000";
					when "01010111001111011" => rgb <= "000000";
					when "01010111001111100" => rgb <= "000000";
					when "01010111001111101" => rgb <= "000000";
					when "01010111001111110" => rgb <= "000000";
					when "01010111001111111" => rgb <= "000000";
					when "01010111010000000" => rgb <= "000000";
					when "01010111010000001" => rgb <= "000000";
					when "01010111010000010" => rgb <= "000000";
					when "01010111010000011" => rgb <= "000000";
					when "01010111010000100" => rgb <= "000000";
					when "01010111010000101" => rgb <= "000000";
					when "01010111010000110" => rgb <= "000000";
					when "01010111010000111" => rgb <= "000000";
					when "01010111010001000" => rgb <= "000000";
					when "01010111010001001" => rgb <= "000000";
					when "01010111010001010" => rgb <= "000000";
					when "01010111010001011" => rgb <= "000000";
					when "01010111010001100" => rgb <= "000000";
					when "01010111010001101" => rgb <= "000000";
					when "01010111010001110" => rgb <= "000000";
					when "01010111010001111" => rgb <= "000000";
					when "01010111010010000" => rgb <= "000000";
					when "01010111010010001" => rgb <= "000000";
					when "01010111010010010" => rgb <= "000000";
					when "01010111010010011" => rgb <= "010100";
					when "01010111010010100" => rgb <= "101000";
					when "01010111010010101" => rgb <= "101000";
					when "01010111010010110" => rgb <= "101000";
					when "01010111010010111" => rgb <= "101000";
					when "01010111010011000" => rgb <= "101000";
					when "01010111010011001" => rgb <= "101000";
					when "01010111010011010" => rgb <= "101000";
					when "01010111010011011" => rgb <= "101000";
					when "01010111010011100" => rgb <= "101000";
					when "01010111010011101" => rgb <= "101000";
					when "01010111010011110" => rgb <= "101000";
					when "01010111010011111" => rgb <= "101000";
					when "01010111010100000" => rgb <= "101000";
					when "01010111010100001" => rgb <= "101000";
					when "01010111010100010" => rgb <= "101000";
					when "01010111010100011" => rgb <= "101000";
					when "01010111010100100" => rgb <= "101000";
					when "01010111010100101" => rgb <= "101000";
					when "01010111010100110" => rgb <= "101000";
					when "01010111010100111" => rgb <= "101000";
					when "01010111010101000" => rgb <= "101000";
					when "01010111010101001" => rgb <= "101000";
					when "01010111010101010" => rgb <= "010000";
					when "01010111010101011" => rgb <= "000000";
					when "01010111010101100" => rgb <= "000000";
					when "01010111010101101" => rgb <= "000000";
					when "01010111010101110" => rgb <= "000000";
					when "01010111010101111" => rgb <= "000000";
					when "01010111010110000" => rgb <= "000000";
					when "01010111010110001" => rgb <= "000000";
					when "01010111010110010" => rgb <= "000000";
					when "01010111010110011" => rgb <= "000000";
					when "01010111010110100" => rgb <= "000000";
					when "01010111010110101" => rgb <= "000000";
					when "01010111010110110" => rgb <= "000000";
					when "01010111010110111" => rgb <= "000000";
					when "01010111010111000" => rgb <= "000000";
					when "01010111010111001" => rgb <= "000000";
					when "01010111010111010" => rgb <= "000000";
					when "01010111010111011" => rgb <= "000000";
					when "01010111010111100" => rgb <= "000000";
					when "01010111010111101" => rgb <= "000000";
					when "01010111010111110" => rgb <= "000000";
					when "01010111010111111" => rgb <= "000000";
					when "01010111011000000" => rgb <= "000000";
					when "01010111011000001" => rgb <= "000000";
					when "01010111011000010" => rgb <= "000000";
					when "01010111011000011" => rgb <= "000000";
					when "01010111011000100" => rgb <= "000000";
					when "01010111011000101" => rgb <= "000000";
					when "01010111011000110" => rgb <= "000000";
					when "01010111011000111" => rgb <= "000000";
					when "01010111011001000" => rgb <= "000000";
					when "01010111011001001" => rgb <= "000000";
					when "01010111011001010" => rgb <= "000000";
					when "01010111011001011" => rgb <= "000000";
					when "01010111011001100" => rgb <= "000000";
					when "01010111011001101" => rgb <= "000000";
					when "01010111011001110" => rgb <= "000000";
					when "01010111011001111" => rgb <= "000000";
					when "01010111011010000" => rgb <= "000000";
					when "01010111011010001" => rgb <= "000000";
					when "01010111011010010" => rgb <= "000000";
					when "01010111011010011" => rgb <= "000000";
					when "01010111011010100" => rgb <= "000000";
					when "01010111011010101" => rgb <= "000000";
					when "01010111011010110" => rgb <= "000000";
					when "01010111011010111" => rgb <= "000000";
					when "01010111011011000" => rgb <= "000000";
					when "01010111011011001" => rgb <= "000000";
					when "01010111011011010" => rgb <= "000000";
					when "01010111011011011" => rgb <= "000000";
					when "01010111011011100" => rgb <= "000000";
					when "01010111011011101" => rgb <= "000000";
					when "01010111011011110" => rgb <= "000000";
					when "01010111011011111" => rgb <= "000000";
					when "01010111011100000" => rgb <= "000000";
					when "01010111011100001" => rgb <= "000000";
					when "01010111011100010" => rgb <= "000000";
					when "01010111011100011" => rgb <= "000000";
					when "01010111011100100" => rgb <= "000000";
					when "01010111011100101" => rgb <= "000000";
					when "01010111011100110" => rgb <= "000000";
					when "01010111011100111" => rgb <= "000000";
					when "01010111011101000" => rgb <= "000000";
					when "01010111011101001" => rgb <= "000000";
					when "01010111011101010" => rgb <= "000000";
					when "01010111011101011" => rgb <= "000000";
					when "01010111011101100" => rgb <= "000000";
					when "01010111011101101" => rgb <= "000000";
					when "01010111011101110" => rgb <= "000000";
					when "01010111011101111" => rgb <= "000000";
					when "01010111011110000" => rgb <= "000000";
					when "01010111011110001" => rgb <= "000000";
					when "01010111011110010" => rgb <= "000000";
					when "01010111011110011" => rgb <= "000000";
					when "01010111011110100" => rgb <= "000000";
					when "01010111011110101" => rgb <= "000000";
					when "01010111011110110" => rgb <= "000000";
					when "01010111011110111" => rgb <= "000000";
					when "01010111011111000" => rgb <= "000000";
					when "01010111011111001" => rgb <= "000000";
					when "01010111011111010" => rgb <= "000000";
					when "01010111011111011" => rgb <= "000000";
					when "01010111011111100" => rgb <= "000000";
					when "01010111011111101" => rgb <= "000000";
					when "01010111011111110" => rgb <= "000000";
					when "01010111011111111" => rgb <= "000000";
					when "01010111100000000" => rgb <= "000000";
					when "01010111100000001" => rgb <= "000000";
					when "01010111100000010" => rgb <= "000000";
					when "01010111100000011" => rgb <= "000000";
					when "01010111100000100" => rgb <= "000000";
					when "01010111100000101" => rgb <= "000000";
					when "01010111100000110" => rgb <= "000000";
					when "01010111100000111" => rgb <= "000000";
					when "01010111100001000" => rgb <= "000000";
					when "01010111100001001" => rgb <= "000000";
					when "01010111100001010" => rgb <= "000000";
					when "01010111100001011" => rgb <= "000000";
					when "01010111100001100" => rgb <= "000000";
					when "01010111100001101" => rgb <= "000000";
					when "01010111100001110" => rgb <= "000000";
					when "01010111100001111" => rgb <= "000000";
					when "01010111100010000" => rgb <= "000000";
					when "01010111100010001" => rgb <= "000000";
					when "01010111100010010" => rgb <= "000000";
					when "01010111100010011" => rgb <= "000000";
					when "01010111100010100" => rgb <= "000000";
					when "01010111100010101" => rgb <= "000000";
					when "01010111100010110" => rgb <= "000000";
					when "01010111100010111" => rgb <= "000000";
					when "01010111100011000" => rgb <= "000000";
					when "01010111100011001" => rgb <= "000000";
					when "01010111100011010" => rgb <= "000000";
					when "01010111100011011" => rgb <= "000000";
					when "01010111100011100" => rgb <= "000000";
					when "01010111100011101" => rgb <= "000000";
					when "01010111100011110" => rgb <= "000000";
					when "01010111100011111" => rgb <= "000000";
					when "01010111100100000" => rgb <= "000000";
					when "01010111100100001" => rgb <= "000000";
					when "01010111100100010" => rgb <= "000000";
					when "01010111100100011" => rgb <= "000000";
					when "01010111100100100" => rgb <= "000000";
					when "01010111100100101" => rgb <= "000000";
					when "01010111100100110" => rgb <= "000000";
					when "01010111100100111" => rgb <= "000000";
					when "01010111100101000" => rgb <= "000000";
					when "01010111100101001" => rgb <= "000000";
					when "01010111100101010" => rgb <= "000000";
					when "01010111100101011" => rgb <= "000000";
					when "01010111100101100" => rgb <= "000000";
					when "01010111100101101" => rgb <= "000000";
					when "01010111100101110" => rgb <= "000000";
					when "01010111100101111" => rgb <= "000000";
					when "01010111100110000" => rgb <= "000000";
					when "01010111100110001" => rgb <= "000000";
					when "01010111100110010" => rgb <= "000000";
					when "01010111100110011" => rgb <= "000000";
					when "01010111100110100" => rgb <= "000000";
					when "01010111100110101" => rgb <= "000000";
					when "01010111100110110" => rgb <= "000000";
					when "01010111100110111" => rgb <= "000000";
					when "01010111100111000" => rgb <= "000000";
					when "01010111100111001" => rgb <= "000000";
					when "01010111100111010" => rgb <= "000000";
					when "01010111100111011" => rgb <= "000000";
					when "01010111100111100" => rgb <= "000000";
					when "01010111100111101" => rgb <= "000000";
					when "01010111100111110" => rgb <= "000000";
					when "01010111100111111" => rgb <= "000000";
					when "01011000000000000" => rgb <= "000000";
					when "01011000000000001" => rgb <= "000000";
					when "01011000000000010" => rgb <= "000000";
					when "01011000000000011" => rgb <= "000000";
					when "01011000000000100" => rgb <= "000000";
					when "01011000000000101" => rgb <= "000000";
					when "01011000000000110" => rgb <= "000000";
					when "01011000000000111" => rgb <= "000000";
					when "01011000000001000" => rgb <= "000000";
					when "01011000000001001" => rgb <= "000000";
					when "01011000000001010" => rgb <= "000000";
					when "01011000000001011" => rgb <= "000000";
					when "01011000000001100" => rgb <= "000000";
					when "01011000000001101" => rgb <= "000000";
					when "01011000000001110" => rgb <= "000000";
					when "01011000000001111" => rgb <= "000000";
					when "01011000000010000" => rgb <= "000000";
					when "01011000000010001" => rgb <= "000000";
					when "01011000000010010" => rgb <= "000000";
					when "01011000000010011" => rgb <= "000000";
					when "01011000000010100" => rgb <= "000000";
					when "01011000000010101" => rgb <= "000000";
					when "01011000000010110" => rgb <= "000000";
					when "01011000000010111" => rgb <= "000000";
					when "01011000000011000" => rgb <= "000000";
					when "01011000000011001" => rgb <= "000000";
					when "01011000000011010" => rgb <= "000000";
					when "01011000000011011" => rgb <= "000000";
					when "01011000000011100" => rgb <= "000000";
					when "01011000000011101" => rgb <= "000000";
					when "01011000000011110" => rgb <= "000000";
					when "01011000000011111" => rgb <= "000000";
					when "01011000000100000" => rgb <= "000000";
					when "01011000000100001" => rgb <= "000000";
					when "01011000000100010" => rgb <= "000000";
					when "01011000000100011" => rgb <= "000000";
					when "01011000000100100" => rgb <= "000000";
					when "01011000000100101" => rgb <= "000000";
					when "01011000000100110" => rgb <= "000000";
					when "01011000000100111" => rgb <= "000000";
					when "01011000000101000" => rgb <= "000000";
					when "01011000000101001" => rgb <= "000000";
					when "01011000000101010" => rgb <= "000000";
					when "01011000000101011" => rgb <= "000000";
					when "01011000000101100" => rgb <= "000000";
					when "01011000000101101" => rgb <= "000000";
					when "01011000000101110" => rgb <= "000000";
					when "01011000000101111" => rgb <= "000000";
					when "01011000000110000" => rgb <= "000000";
					when "01011000000110001" => rgb <= "000000";
					when "01011000000110010" => rgb <= "000000";
					when "01011000000110011" => rgb <= "000000";
					when "01011000000110100" => rgb <= "000000";
					when "01011000000110101" => rgb <= "000000";
					when "01011000000110110" => rgb <= "000000";
					when "01011000000110111" => rgb <= "000000";
					when "01011000000111000" => rgb <= "000000";
					when "01011000000111001" => rgb <= "000000";
					when "01011000000111010" => rgb <= "000000";
					when "01011000000111011" => rgb <= "000000";
					when "01011000000111100" => rgb <= "000000";
					when "01011000000111101" => rgb <= "000000";
					when "01011000000111110" => rgb <= "000000";
					when "01011000000111111" => rgb <= "000000";
					when "01011000001000000" => rgb <= "000000";
					when "01011000001000001" => rgb <= "000000";
					when "01011000001000010" => rgb <= "000000";
					when "01011000001000011" => rgb <= "000000";
					when "01011000001000100" => rgb <= "000000";
					when "01011000001000101" => rgb <= "000000";
					when "01011000001000110" => rgb <= "000000";
					when "01011000001000111" => rgb <= "000000";
					when "01011000001001000" => rgb <= "000000";
					when "01011000001001001" => rgb <= "000000";
					when "01011000001001010" => rgb <= "000000";
					when "01011000001001011" => rgb <= "000000";
					when "01011000001001100" => rgb <= "000000";
					when "01011000001001101" => rgb <= "000000";
					when "01011000001001110" => rgb <= "000000";
					when "01011000001001111" => rgb <= "000000";
					when "01011000001010000" => rgb <= "000000";
					when "01011000001010001" => rgb <= "000000";
					when "01011000001010010" => rgb <= "000000";
					when "01011000001010011" => rgb <= "000000";
					when "01011000001010100" => rgb <= "000000";
					when "01011000001010101" => rgb <= "000000";
					when "01011000001010110" => rgb <= "000000";
					when "01011000001010111" => rgb <= "000000";
					when "01011000001011000" => rgb <= "000000";
					when "01011000001011001" => rgb <= "000000";
					when "01011000001011010" => rgb <= "000000";
					when "01011000001011011" => rgb <= "000000";
					when "01011000001011100" => rgb <= "000000";
					when "01011000001011101" => rgb <= "000000";
					when "01011000001011110" => rgb <= "000000";
					when "01011000001011111" => rgb <= "000000";
					when "01011000001100000" => rgb <= "000000";
					when "01011000001100001" => rgb <= "000000";
					when "01011000001100010" => rgb <= "000000";
					when "01011000001100011" => rgb <= "000000";
					when "01011000001100100" => rgb <= "000000";
					when "01011000001100101" => rgb <= "000000";
					when "01011000001100110" => rgb <= "000000";
					when "01011000001100111" => rgb <= "000000";
					when "01011000001101000" => rgb <= "000000";
					when "01011000001101001" => rgb <= "000000";
					when "01011000001101010" => rgb <= "000000";
					when "01011000001101011" => rgb <= "000000";
					when "01011000001101100" => rgb <= "000000";
					when "01011000001101101" => rgb <= "000000";
					when "01011000001101110" => rgb <= "000000";
					when "01011000001101111" => rgb <= "000000";
					when "01011000001110000" => rgb <= "000000";
					when "01011000001110001" => rgb <= "000000";
					when "01011000001110010" => rgb <= "000000";
					when "01011000001110011" => rgb <= "000000";
					when "01011000001110100" => rgb <= "000000";
					when "01011000001110101" => rgb <= "000000";
					when "01011000001110110" => rgb <= "000000";
					when "01011000001110111" => rgb <= "000000";
					when "01011000001111000" => rgb <= "000000";
					when "01011000001111001" => rgb <= "000000";
					when "01011000001111010" => rgb <= "000000";
					when "01011000001111011" => rgb <= "000000";
					when "01011000001111100" => rgb <= "000000";
					when "01011000001111101" => rgb <= "000000";
					when "01011000001111110" => rgb <= "000000";
					when "01011000001111111" => rgb <= "000000";
					when "01011000010000000" => rgb <= "000000";
					when "01011000010000001" => rgb <= "000000";
					when "01011000010000010" => rgb <= "000000";
					when "01011000010000011" => rgb <= "000000";
					when "01011000010000100" => rgb <= "000000";
					when "01011000010000101" => rgb <= "000000";
					when "01011000010000110" => rgb <= "000000";
					when "01011000010000111" => rgb <= "000000";
					when "01011000010001000" => rgb <= "000000";
					when "01011000010001001" => rgb <= "000000";
					when "01011000010001010" => rgb <= "000000";
					when "01011000010001011" => rgb <= "000000";
					when "01011000010001100" => rgb <= "000000";
					when "01011000010001101" => rgb <= "000000";
					when "01011000010001110" => rgb <= "000000";
					when "01011000010001111" => rgb <= "000000";
					when "01011000010010000" => rgb <= "000000";
					when "01011000010010001" => rgb <= "000000";
					when "01011000010010010" => rgb <= "000000";
					when "01011000010010011" => rgb <= "010100";
					when "01011000010010100" => rgb <= "111000";
					when "01011000010010101" => rgb <= "101000";
					when "01011000010010110" => rgb <= "101000";
					when "01011000010010111" => rgb <= "101000";
					when "01011000010011000" => rgb <= "101000";
					when "01011000010011001" => rgb <= "101000";
					when "01011000010011010" => rgb <= "101000";
					when "01011000010011011" => rgb <= "101000";
					when "01011000010011100" => rgb <= "101000";
					when "01011000010011101" => rgb <= "101000";
					when "01011000010011110" => rgb <= "101000";
					when "01011000010011111" => rgb <= "101000";
					when "01011000010100000" => rgb <= "101000";
					when "01011000010100001" => rgb <= "101000";
					when "01011000010100010" => rgb <= "101000";
					when "01011000010100011" => rgb <= "101000";
					when "01011000010100100" => rgb <= "101000";
					when "01011000010100101" => rgb <= "101000";
					when "01011000010100110" => rgb <= "101000";
					when "01011000010100111" => rgb <= "101000";
					when "01011000010101000" => rgb <= "101000";
					when "01011000010101001" => rgb <= "101000";
					when "01011000010101010" => rgb <= "010000";
					when "01011000010101011" => rgb <= "000000";
					when "01011000010101100" => rgb <= "000000";
					when "01011000010101101" => rgb <= "000000";
					when "01011000010101110" => rgb <= "000000";
					when "01011000010101111" => rgb <= "000000";
					when "01011000010110000" => rgb <= "000000";
					when "01011000010110001" => rgb <= "000000";
					when "01011000010110010" => rgb <= "000000";
					when "01011000010110011" => rgb <= "000000";
					when "01011000010110100" => rgb <= "000000";
					when "01011000010110101" => rgb <= "000000";
					when "01011000010110110" => rgb <= "000000";
					when "01011000010110111" => rgb <= "000000";
					when "01011000010111000" => rgb <= "000000";
					when "01011000010111001" => rgb <= "000000";
					when "01011000010111010" => rgb <= "000000";
					when "01011000010111011" => rgb <= "000000";
					when "01011000010111100" => rgb <= "000000";
					when "01011000010111101" => rgb <= "000000";
					when "01011000010111110" => rgb <= "000000";
					when "01011000010111111" => rgb <= "000000";
					when "01011000011000000" => rgb <= "000000";
					when "01011000011000001" => rgb <= "000000";
					when "01011000011000010" => rgb <= "000000";
					when "01011000011000011" => rgb <= "000000";
					when "01011000011000100" => rgb <= "000000";
					when "01011000011000101" => rgb <= "000000";
					when "01011000011000110" => rgb <= "000000";
					when "01011000011000111" => rgb <= "000000";
					when "01011000011001000" => rgb <= "000000";
					when "01011000011001001" => rgb <= "000000";
					when "01011000011001010" => rgb <= "000000";
					when "01011000011001011" => rgb <= "000000";
					when "01011000011001100" => rgb <= "000000";
					when "01011000011001101" => rgb <= "000000";
					when "01011000011001110" => rgb <= "000000";
					when "01011000011001111" => rgb <= "000000";
					when "01011000011010000" => rgb <= "000000";
					when "01011000011010001" => rgb <= "000000";
					when "01011000011010010" => rgb <= "000000";
					when "01011000011010011" => rgb <= "000000";
					when "01011000011010100" => rgb <= "000000";
					when "01011000011010101" => rgb <= "000000";
					when "01011000011010110" => rgb <= "000000";
					when "01011000011010111" => rgb <= "000000";
					when "01011000011011000" => rgb <= "000000";
					when "01011000011011001" => rgb <= "000000";
					when "01011000011011010" => rgb <= "000000";
					when "01011000011011011" => rgb <= "000000";
					when "01011000011011100" => rgb <= "000000";
					when "01011000011011101" => rgb <= "000000";
					when "01011000011011110" => rgb <= "000000";
					when "01011000011011111" => rgb <= "000000";
					when "01011000011100000" => rgb <= "000000";
					when "01011000011100001" => rgb <= "000000";
					when "01011000011100010" => rgb <= "000000";
					when "01011000011100011" => rgb <= "000000";
					when "01011000011100100" => rgb <= "000000";
					when "01011000011100101" => rgb <= "000000";
					when "01011000011100110" => rgb <= "000000";
					when "01011000011100111" => rgb <= "000000";
					when "01011000011101000" => rgb <= "000000";
					when "01011000011101001" => rgb <= "000000";
					when "01011000011101010" => rgb <= "000000";
					when "01011000011101011" => rgb <= "000000";
					when "01011000011101100" => rgb <= "000000";
					when "01011000011101101" => rgb <= "000000";
					when "01011000011101110" => rgb <= "000000";
					when "01011000011101111" => rgb <= "000000";
					when "01011000011110000" => rgb <= "000000";
					when "01011000011110001" => rgb <= "000000";
					when "01011000011110010" => rgb <= "000000";
					when "01011000011110011" => rgb <= "000000";
					when "01011000011110100" => rgb <= "000000";
					when "01011000011110101" => rgb <= "000000";
					when "01011000011110110" => rgb <= "000000";
					when "01011000011110111" => rgb <= "000000";
					when "01011000011111000" => rgb <= "000000";
					when "01011000011111001" => rgb <= "000000";
					when "01011000011111010" => rgb <= "000000";
					when "01011000011111011" => rgb <= "000000";
					when "01011000011111100" => rgb <= "000000";
					when "01011000011111101" => rgb <= "000000";
					when "01011000011111110" => rgb <= "000000";
					when "01011000011111111" => rgb <= "000000";
					when "01011000100000000" => rgb <= "000000";
					when "01011000100000001" => rgb <= "000000";
					when "01011000100000010" => rgb <= "000000";
					when "01011000100000011" => rgb <= "000000";
					when "01011000100000100" => rgb <= "000000";
					when "01011000100000101" => rgb <= "000000";
					when "01011000100000110" => rgb <= "000000";
					when "01011000100000111" => rgb <= "000000";
					when "01011000100001000" => rgb <= "000000";
					when "01011000100001001" => rgb <= "000000";
					when "01011000100001010" => rgb <= "000000";
					when "01011000100001011" => rgb <= "000000";
					when "01011000100001100" => rgb <= "000000";
					when "01011000100001101" => rgb <= "000000";
					when "01011000100001110" => rgb <= "000000";
					when "01011000100001111" => rgb <= "000000";
					when "01011000100010000" => rgb <= "000000";
					when "01011000100010001" => rgb <= "000000";
					when "01011000100010010" => rgb <= "000000";
					when "01011000100010011" => rgb <= "000000";
					when "01011000100010100" => rgb <= "000000";
					when "01011000100010101" => rgb <= "000000";
					when "01011000100010110" => rgb <= "000000";
					when "01011000100010111" => rgb <= "000000";
					when "01011000100011000" => rgb <= "000000";
					when "01011000100011001" => rgb <= "000000";
					when "01011000100011010" => rgb <= "000000";
					when "01011000100011011" => rgb <= "000000";
					when "01011000100011100" => rgb <= "000000";
					when "01011000100011101" => rgb <= "000000";
					when "01011000100011110" => rgb <= "000000";
					when "01011000100011111" => rgb <= "000000";
					when "01011000100100000" => rgb <= "000000";
					when "01011000100100001" => rgb <= "000000";
					when "01011000100100010" => rgb <= "000000";
					when "01011000100100011" => rgb <= "000000";
					when "01011000100100100" => rgb <= "000000";
					when "01011000100100101" => rgb <= "000000";
					when "01011000100100110" => rgb <= "000000";
					when "01011000100100111" => rgb <= "000000";
					when "01011000100101000" => rgb <= "000000";
					when "01011000100101001" => rgb <= "000000";
					when "01011000100101010" => rgb <= "000000";
					when "01011000100101011" => rgb <= "000000";
					when "01011000100101100" => rgb <= "000000";
					when "01011000100101101" => rgb <= "000000";
					when "01011000100101110" => rgb <= "000000";
					when "01011000100101111" => rgb <= "000000";
					when "01011000100110000" => rgb <= "000000";
					when "01011000100110001" => rgb <= "000000";
					when "01011000100110010" => rgb <= "000000";
					when "01011000100110011" => rgb <= "000000";
					when "01011000100110100" => rgb <= "000000";
					when "01011000100110101" => rgb <= "000000";
					when "01011000100110110" => rgb <= "000000";
					when "01011000100110111" => rgb <= "000000";
					when "01011000100111000" => rgb <= "000000";
					when "01011000100111001" => rgb <= "000000";
					when "01011000100111010" => rgb <= "000000";
					when "01011000100111011" => rgb <= "000000";
					when "01011000100111100" => rgb <= "000000";
					when "01011000100111101" => rgb <= "000000";
					when "01011000100111110" => rgb <= "000000";
					when "01011000100111111" => rgb <= "000000";
					when "01011001000000000" => rgb <= "000000";
					when "01011001000000001" => rgb <= "000000";
					when "01011001000000010" => rgb <= "000000";
					when "01011001000000011" => rgb <= "000000";
					when "01011001000000100" => rgb <= "000000";
					when "01011001000000101" => rgb <= "000000";
					when "01011001000000110" => rgb <= "000000";
					when "01011001000000111" => rgb <= "000000";
					when "01011001000001000" => rgb <= "000000";
					when "01011001000001001" => rgb <= "000000";
					when "01011001000001010" => rgb <= "000000";
					when "01011001000001011" => rgb <= "000000";
					when "01011001000001100" => rgb <= "000000";
					when "01011001000001101" => rgb <= "000000";
					when "01011001000001110" => rgb <= "000000";
					when "01011001000001111" => rgb <= "000000";
					when "01011001000010000" => rgb <= "000000";
					when "01011001000010001" => rgb <= "000000";
					when "01011001000010010" => rgb <= "000000";
					when "01011001000010011" => rgb <= "000000";
					when "01011001000010100" => rgb <= "000000";
					when "01011001000010101" => rgb <= "000000";
					when "01011001000010110" => rgb <= "000000";
					when "01011001000010111" => rgb <= "000000";
					when "01011001000011000" => rgb <= "000000";
					when "01011001000011001" => rgb <= "000000";
					when "01011001000011010" => rgb <= "000000";
					when "01011001000011011" => rgb <= "000000";
					when "01011001000011100" => rgb <= "000000";
					when "01011001000011101" => rgb <= "000000";
					when "01011001000011110" => rgb <= "000000";
					when "01011001000011111" => rgb <= "000000";
					when "01011001000100000" => rgb <= "000000";
					when "01011001000100001" => rgb <= "000000";
					when "01011001000100010" => rgb <= "000000";
					when "01011001000100011" => rgb <= "000000";
					when "01011001000100100" => rgb <= "000000";
					when "01011001000100101" => rgb <= "000000";
					when "01011001000100110" => rgb <= "000000";
					when "01011001000100111" => rgb <= "000000";
					when "01011001000101000" => rgb <= "000000";
					when "01011001000101001" => rgb <= "000000";
					when "01011001000101010" => rgb <= "000000";
					when "01011001000101011" => rgb <= "000000";
					when "01011001000101100" => rgb <= "000000";
					when "01011001000101101" => rgb <= "000000";
					when "01011001000101110" => rgb <= "000000";
					when "01011001000101111" => rgb <= "000000";
					when "01011001000110000" => rgb <= "000000";
					when "01011001000110001" => rgb <= "000000";
					when "01011001000110010" => rgb <= "000000";
					when "01011001000110011" => rgb <= "000000";
					when "01011001000110100" => rgb <= "000000";
					when "01011001000110101" => rgb <= "000000";
					when "01011001000110110" => rgb <= "000000";
					when "01011001000110111" => rgb <= "000000";
					when "01011001000111000" => rgb <= "000000";
					when "01011001000111001" => rgb <= "000000";
					when "01011001000111010" => rgb <= "000000";
					when "01011001000111011" => rgb <= "000000";
					when "01011001000111100" => rgb <= "000000";
					when "01011001000111101" => rgb <= "000000";
					when "01011001000111110" => rgb <= "000000";
					when "01011001000111111" => rgb <= "000000";
					when "01011001001000000" => rgb <= "000000";
					when "01011001001000001" => rgb <= "000000";
					when "01011001001000010" => rgb <= "000000";
					when "01011001001000011" => rgb <= "000000";
					when "01011001001000100" => rgb <= "000000";
					when "01011001001000101" => rgb <= "000000";
					when "01011001001000110" => rgb <= "000000";
					when "01011001001000111" => rgb <= "000000";
					when "01011001001001000" => rgb <= "000000";
					when "01011001001001001" => rgb <= "000000";
					when "01011001001001010" => rgb <= "000000";
					when "01011001001001011" => rgb <= "000000";
					when "01011001001001100" => rgb <= "000000";
					when "01011001001001101" => rgb <= "000000";
					when "01011001001001110" => rgb <= "000000";
					when "01011001001001111" => rgb <= "000000";
					when "01011001001010000" => rgb <= "000000";
					when "01011001001010001" => rgb <= "000000";
					when "01011001001010010" => rgb <= "000000";
					when "01011001001010011" => rgb <= "000000";
					when "01011001001010100" => rgb <= "000000";
					when "01011001001010101" => rgb <= "000000";
					when "01011001001010110" => rgb <= "000000";
					when "01011001001010111" => rgb <= "000000";
					when "01011001001011000" => rgb <= "000000";
					when "01011001001011001" => rgb <= "000000";
					when "01011001001011010" => rgb <= "000000";
					when "01011001001011011" => rgb <= "000000";
					when "01011001001011100" => rgb <= "000000";
					when "01011001001011101" => rgb <= "000000";
					when "01011001001011110" => rgb <= "000000";
					when "01011001001011111" => rgb <= "000000";
					when "01011001001100000" => rgb <= "000000";
					when "01011001001100001" => rgb <= "000000";
					when "01011001001100010" => rgb <= "000000";
					when "01011001001100011" => rgb <= "000000";
					when "01011001001100100" => rgb <= "000000";
					when "01011001001100101" => rgb <= "000000";
					when "01011001001100110" => rgb <= "000000";
					when "01011001001100111" => rgb <= "000000";
					when "01011001001101000" => rgb <= "000000";
					when "01011001001101001" => rgb <= "000000";
					when "01011001001101010" => rgb <= "000000";
					when "01011001001101011" => rgb <= "000000";
					when "01011001001101100" => rgb <= "000000";
					when "01011001001101101" => rgb <= "000000";
					when "01011001001101110" => rgb <= "000000";
					when "01011001001101111" => rgb <= "000000";
					when "01011001001110000" => rgb <= "000000";
					when "01011001001110001" => rgb <= "000000";
					when "01011001001110010" => rgb <= "000000";
					when "01011001001110011" => rgb <= "000000";
					when "01011001001110100" => rgb <= "000000";
					when "01011001001110101" => rgb <= "000000";
					when "01011001001110110" => rgb <= "000000";
					when "01011001001110111" => rgb <= "000000";
					when "01011001001111000" => rgb <= "000000";
					when "01011001001111001" => rgb <= "000000";
					when "01011001001111010" => rgb <= "000000";
					when "01011001001111011" => rgb <= "000000";
					when "01011001001111100" => rgb <= "000000";
					when "01011001001111101" => rgb <= "000000";
					when "01011001001111110" => rgb <= "000000";
					when "01011001001111111" => rgb <= "000000";
					when "01011001010000000" => rgb <= "000000";
					when "01011001010000001" => rgb <= "000000";
					when "01011001010000010" => rgb <= "000000";
					when "01011001010000011" => rgb <= "000000";
					when "01011001010000100" => rgb <= "000000";
					when "01011001010000101" => rgb <= "000000";
					when "01011001010000110" => rgb <= "000000";
					when "01011001010000111" => rgb <= "000000";
					when "01011001010001000" => rgb <= "000000";
					when "01011001010001001" => rgb <= "000000";
					when "01011001010001010" => rgb <= "000000";
					when "01011001010001011" => rgb <= "000000";
					when "01011001010001100" => rgb <= "000000";
					when "01011001010001101" => rgb <= "000000";
					when "01011001010001110" => rgb <= "000000";
					when "01011001010001111" => rgb <= "000000";
					when "01011001010010000" => rgb <= "000000";
					when "01011001010010001" => rgb <= "000000";
					when "01011001010010010" => rgb <= "000000";
					when "01011001010010011" => rgb <= "010100";
					when "01011001010010100" => rgb <= "111000";
					when "01011001010010101" => rgb <= "101000";
					when "01011001010010110" => rgb <= "101000";
					when "01011001010010111" => rgb <= "101000";
					when "01011001010011000" => rgb <= "101000";
					when "01011001010011001" => rgb <= "101000";
					when "01011001010011010" => rgb <= "101000";
					when "01011001010011011" => rgb <= "101000";
					when "01011001010011100" => rgb <= "101000";
					when "01011001010011101" => rgb <= "101000";
					when "01011001010011110" => rgb <= "101000";
					when "01011001010011111" => rgb <= "101000";
					when "01011001010100000" => rgb <= "101000";
					when "01011001010100001" => rgb <= "101000";
					when "01011001010100010" => rgb <= "101000";
					when "01011001010100011" => rgb <= "101000";
					when "01011001010100100" => rgb <= "101000";
					when "01011001010100101" => rgb <= "101000";
					when "01011001010100110" => rgb <= "101000";
					when "01011001010100111" => rgb <= "101000";
					when "01011001010101000" => rgb <= "101000";
					when "01011001010101001" => rgb <= "101000";
					when "01011001010101010" => rgb <= "010000";
					when "01011001010101011" => rgb <= "000000";
					when "01011001010101100" => rgb <= "000000";
					when "01011001010101101" => rgb <= "000000";
					when "01011001010101110" => rgb <= "000000";
					when "01011001010101111" => rgb <= "000000";
					when "01011001010110000" => rgb <= "000000";
					when "01011001010110001" => rgb <= "000000";
					when "01011001010110010" => rgb <= "000000";
					when "01011001010110011" => rgb <= "000000";
					when "01011001010110100" => rgb <= "000000";
					when "01011001010110101" => rgb <= "000000";
					when "01011001010110110" => rgb <= "000000";
					when "01011001010110111" => rgb <= "000000";
					when "01011001010111000" => rgb <= "000000";
					when "01011001010111001" => rgb <= "000000";
					when "01011001010111010" => rgb <= "000000";
					when "01011001010111011" => rgb <= "000000";
					when "01011001010111100" => rgb <= "000000";
					when "01011001010111101" => rgb <= "000000";
					when "01011001010111110" => rgb <= "000000";
					when "01011001010111111" => rgb <= "000000";
					when "01011001011000000" => rgb <= "000000";
					when "01011001011000001" => rgb <= "000000";
					when "01011001011000010" => rgb <= "000000";
					when "01011001011000011" => rgb <= "000000";
					when "01011001011000100" => rgb <= "000000";
					when "01011001011000101" => rgb <= "000000";
					when "01011001011000110" => rgb <= "000000";
					when "01011001011000111" => rgb <= "000000";
					when "01011001011001000" => rgb <= "000000";
					when "01011001011001001" => rgb <= "000000";
					when "01011001011001010" => rgb <= "000000";
					when "01011001011001011" => rgb <= "000000";
					when "01011001011001100" => rgb <= "000000";
					when "01011001011001101" => rgb <= "000000";
					when "01011001011001110" => rgb <= "000000";
					when "01011001011001111" => rgb <= "000000";
					when "01011001011010000" => rgb <= "000000";
					when "01011001011010001" => rgb <= "000000";
					when "01011001011010010" => rgb <= "000000";
					when "01011001011010011" => rgb <= "000000";
					when "01011001011010100" => rgb <= "000000";
					when "01011001011010101" => rgb <= "000000";
					when "01011001011010110" => rgb <= "000000";
					when "01011001011010111" => rgb <= "000000";
					when "01011001011011000" => rgb <= "000000";
					when "01011001011011001" => rgb <= "000000";
					when "01011001011011010" => rgb <= "000000";
					when "01011001011011011" => rgb <= "000000";
					when "01011001011011100" => rgb <= "000000";
					when "01011001011011101" => rgb <= "000000";
					when "01011001011011110" => rgb <= "000000";
					when "01011001011011111" => rgb <= "000000";
					when "01011001011100000" => rgb <= "000000";
					when "01011001011100001" => rgb <= "000000";
					when "01011001011100010" => rgb <= "000000";
					when "01011001011100011" => rgb <= "000000";
					when "01011001011100100" => rgb <= "000000";
					when "01011001011100101" => rgb <= "000000";
					when "01011001011100110" => rgb <= "000000";
					when "01011001011100111" => rgb <= "000000";
					when "01011001011101000" => rgb <= "000000";
					when "01011001011101001" => rgb <= "000000";
					when "01011001011101010" => rgb <= "000000";
					when "01011001011101011" => rgb <= "000000";
					when "01011001011101100" => rgb <= "000000";
					when "01011001011101101" => rgb <= "000000";
					when "01011001011101110" => rgb <= "000000";
					when "01011001011101111" => rgb <= "000000";
					when "01011001011110000" => rgb <= "000000";
					when "01011001011110001" => rgb <= "000000";
					when "01011001011110010" => rgb <= "000000";
					when "01011001011110011" => rgb <= "000000";
					when "01011001011110100" => rgb <= "000000";
					when "01011001011110101" => rgb <= "000000";
					when "01011001011110110" => rgb <= "000000";
					when "01011001011110111" => rgb <= "000000";
					when "01011001011111000" => rgb <= "000000";
					when "01011001011111001" => rgb <= "000000";
					when "01011001011111010" => rgb <= "000000";
					when "01011001011111011" => rgb <= "000000";
					when "01011001011111100" => rgb <= "000000";
					when "01011001011111101" => rgb <= "000000";
					when "01011001011111110" => rgb <= "000000";
					when "01011001011111111" => rgb <= "000000";
					when "01011001100000000" => rgb <= "000000";
					when "01011001100000001" => rgb <= "000000";
					when "01011001100000010" => rgb <= "000000";
					when "01011001100000011" => rgb <= "000000";
					when "01011001100000100" => rgb <= "000000";
					when "01011001100000101" => rgb <= "000000";
					when "01011001100000110" => rgb <= "000000";
					when "01011001100000111" => rgb <= "000000";
					when "01011001100001000" => rgb <= "000000";
					when "01011001100001001" => rgb <= "000000";
					when "01011001100001010" => rgb <= "000000";
					when "01011001100001011" => rgb <= "000000";
					when "01011001100001100" => rgb <= "000000";
					when "01011001100001101" => rgb <= "000000";
					when "01011001100001110" => rgb <= "000000";
					when "01011001100001111" => rgb <= "000000";
					when "01011001100010000" => rgb <= "000000";
					when "01011001100010001" => rgb <= "000000";
					when "01011001100010010" => rgb <= "000000";
					when "01011001100010011" => rgb <= "000000";
					when "01011001100010100" => rgb <= "000000";
					when "01011001100010101" => rgb <= "000000";
					when "01011001100010110" => rgb <= "000000";
					when "01011001100010111" => rgb <= "000000";
					when "01011001100011000" => rgb <= "000000";
					when "01011001100011001" => rgb <= "000000";
					when "01011001100011010" => rgb <= "000000";
					when "01011001100011011" => rgb <= "000000";
					when "01011001100011100" => rgb <= "000000";
					when "01011001100011101" => rgb <= "000000";
					when "01011001100011110" => rgb <= "000000";
					when "01011001100011111" => rgb <= "000000";
					when "01011001100100000" => rgb <= "000000";
					when "01011001100100001" => rgb <= "000000";
					when "01011001100100010" => rgb <= "000000";
					when "01011001100100011" => rgb <= "000000";
					when "01011001100100100" => rgb <= "000000";
					when "01011001100100101" => rgb <= "000000";
					when "01011001100100110" => rgb <= "000000";
					when "01011001100100111" => rgb <= "000000";
					when "01011001100101000" => rgb <= "000000";
					when "01011001100101001" => rgb <= "000000";
					when "01011001100101010" => rgb <= "000000";
					when "01011001100101011" => rgb <= "000000";
					when "01011001100101100" => rgb <= "000000";
					when "01011001100101101" => rgb <= "000000";
					when "01011001100101110" => rgb <= "000000";
					when "01011001100101111" => rgb <= "000000";
					when "01011001100110000" => rgb <= "000000";
					when "01011001100110001" => rgb <= "000000";
					when "01011001100110010" => rgb <= "000000";
					when "01011001100110011" => rgb <= "000000";
					when "01011001100110100" => rgb <= "000000";
					when "01011001100110101" => rgb <= "000000";
					when "01011001100110110" => rgb <= "000000";
					when "01011001100110111" => rgb <= "000000";
					when "01011001100111000" => rgb <= "000000";
					when "01011001100111001" => rgb <= "000000";
					when "01011001100111010" => rgb <= "000000";
					when "01011001100111011" => rgb <= "000000";
					when "01011001100111100" => rgb <= "000000";
					when "01011001100111101" => rgb <= "000000";
					when "01011001100111110" => rgb <= "000000";
					when "01011001100111111" => rgb <= "000000";
					when "01011010000000000" => rgb <= "000000";
					when "01011010000000001" => rgb <= "000000";
					when "01011010000000010" => rgb <= "000000";
					when "01011010000000011" => rgb <= "000000";
					when "01011010000000100" => rgb <= "000000";
					when "01011010000000101" => rgb <= "000000";
					when "01011010000000110" => rgb <= "000000";
					when "01011010000000111" => rgb <= "000000";
					when "01011010000001000" => rgb <= "000000";
					when "01011010000001001" => rgb <= "000000";
					when "01011010000001010" => rgb <= "000000";
					when "01011010000001011" => rgb <= "000000";
					when "01011010000001100" => rgb <= "000000";
					when "01011010000001101" => rgb <= "000000";
					when "01011010000001110" => rgb <= "000000";
					when "01011010000001111" => rgb <= "000000";
					when "01011010000010000" => rgb <= "000000";
					when "01011010000010001" => rgb <= "000000";
					when "01011010000010010" => rgb <= "000000";
					when "01011010000010011" => rgb <= "000000";
					when "01011010000010100" => rgb <= "000000";
					when "01011010000010101" => rgb <= "000000";
					when "01011010000010110" => rgb <= "000000";
					when "01011010000010111" => rgb <= "000000";
					when "01011010000011000" => rgb <= "000000";
					when "01011010000011001" => rgb <= "000000";
					when "01011010000011010" => rgb <= "000000";
					when "01011010000011011" => rgb <= "000000";
					when "01011010000011100" => rgb <= "000000";
					when "01011010000011101" => rgb <= "000000";
					when "01011010000011110" => rgb <= "000000";
					when "01011010000011111" => rgb <= "000000";
					when "01011010000100000" => rgb <= "000000";
					when "01011010000100001" => rgb <= "000000";
					when "01011010000100010" => rgb <= "000000";
					when "01011010000100011" => rgb <= "000000";
					when "01011010000100100" => rgb <= "000000";
					when "01011010000100101" => rgb <= "000000";
					when "01011010000100110" => rgb <= "000000";
					when "01011010000100111" => rgb <= "000000";
					when "01011010000101000" => rgb <= "000000";
					when "01011010000101001" => rgb <= "000000";
					when "01011010000101010" => rgb <= "000000";
					when "01011010000101011" => rgb <= "000000";
					when "01011010000101100" => rgb <= "000000";
					when "01011010000101101" => rgb <= "000000";
					when "01011010000101110" => rgb <= "000000";
					when "01011010000101111" => rgb <= "000000";
					when "01011010000110000" => rgb <= "000000";
					when "01011010000110001" => rgb <= "000000";
					when "01011010000110010" => rgb <= "000000";
					when "01011010000110011" => rgb <= "000000";
					when "01011010000110100" => rgb <= "000000";
					when "01011010000110101" => rgb <= "000000";
					when "01011010000110110" => rgb <= "000000";
					when "01011010000110111" => rgb <= "000000";
					when "01011010000111000" => rgb <= "000000";
					when "01011010000111001" => rgb <= "000000";
					when "01011010000111010" => rgb <= "000000";
					when "01011010000111011" => rgb <= "000000";
					when "01011010000111100" => rgb <= "000000";
					when "01011010000111101" => rgb <= "000000";
					when "01011010000111110" => rgb <= "000000";
					when "01011010000111111" => rgb <= "000000";
					when "01011010001000000" => rgb <= "000000";
					when "01011010001000001" => rgb <= "000000";
					when "01011010001000010" => rgb <= "000000";
					when "01011010001000011" => rgb <= "000000";
					when "01011010001000100" => rgb <= "000000";
					when "01011010001000101" => rgb <= "000000";
					when "01011010001000110" => rgb <= "000000";
					when "01011010001000111" => rgb <= "000000";
					when "01011010001001000" => rgb <= "000000";
					when "01011010001001001" => rgb <= "000000";
					when "01011010001001010" => rgb <= "000000";
					when "01011010001001011" => rgb <= "000000";
					when "01011010001001100" => rgb <= "000000";
					when "01011010001001101" => rgb <= "000000";
					when "01011010001001110" => rgb <= "000000";
					when "01011010001001111" => rgb <= "000000";
					when "01011010001010000" => rgb <= "000000";
					when "01011010001010001" => rgb <= "000000";
					when "01011010001010010" => rgb <= "000000";
					when "01011010001010011" => rgb <= "000000";
					when "01011010001010100" => rgb <= "000000";
					when "01011010001010101" => rgb <= "000000";
					when "01011010001010110" => rgb <= "000000";
					when "01011010001010111" => rgb <= "000000";
					when "01011010001011000" => rgb <= "000000";
					when "01011010001011001" => rgb <= "000000";
					when "01011010001011010" => rgb <= "000000";
					when "01011010001011011" => rgb <= "000000";
					when "01011010001011100" => rgb <= "000000";
					when "01011010001011101" => rgb <= "000000";
					when "01011010001011110" => rgb <= "000000";
					when "01011010001011111" => rgb <= "000000";
					when "01011010001100000" => rgb <= "000000";
					when "01011010001100001" => rgb <= "000000";
					when "01011010001100010" => rgb <= "000000";
					when "01011010001100011" => rgb <= "000000";
					when "01011010001100100" => rgb <= "000000";
					when "01011010001100101" => rgb <= "000000";
					when "01011010001100110" => rgb <= "000000";
					when "01011010001100111" => rgb <= "000000";
					when "01011010001101000" => rgb <= "000000";
					when "01011010001101001" => rgb <= "000000";
					when "01011010001101010" => rgb <= "000000";
					when "01011010001101011" => rgb <= "000000";
					when "01011010001101100" => rgb <= "000000";
					when "01011010001101101" => rgb <= "000000";
					when "01011010001101110" => rgb <= "000000";
					when "01011010001101111" => rgb <= "000000";
					when "01011010001110000" => rgb <= "000000";
					when "01011010001110001" => rgb <= "000000";
					when "01011010001110010" => rgb <= "000000";
					when "01011010001110011" => rgb <= "000000";
					when "01011010001110100" => rgb <= "000000";
					when "01011010001110101" => rgb <= "000000";
					when "01011010001110110" => rgb <= "000000";
					when "01011010001110111" => rgb <= "000000";
					when "01011010001111000" => rgb <= "000000";
					when "01011010001111001" => rgb <= "000000";
					when "01011010001111010" => rgb <= "000000";
					when "01011010001111011" => rgb <= "000000";
					when "01011010001111100" => rgb <= "000000";
					when "01011010001111101" => rgb <= "000000";
					when "01011010001111110" => rgb <= "000000";
					when "01011010001111111" => rgb <= "000000";
					when "01011010010000000" => rgb <= "000000";
					when "01011010010000001" => rgb <= "000000";
					when "01011010010000010" => rgb <= "000000";
					when "01011010010000011" => rgb <= "000000";
					when "01011010010000100" => rgb <= "000000";
					when "01011010010000101" => rgb <= "000000";
					when "01011010010000110" => rgb <= "000000";
					when "01011010010000111" => rgb <= "000000";
					when "01011010010001000" => rgb <= "000000";
					when "01011010010001001" => rgb <= "000000";
					when "01011010010001010" => rgb <= "000000";
					when "01011010010001011" => rgb <= "000000";
					when "01011010010001100" => rgb <= "000000";
					when "01011010010001101" => rgb <= "000000";
					when "01011010010001110" => rgb <= "000000";
					when "01011010010001111" => rgb <= "000000";
					when "01011010010010000" => rgb <= "000000";
					when "01011010010010001" => rgb <= "000000";
					when "01011010010010010" => rgb <= "000000";
					when "01011010010010011" => rgb <= "010100";
					when "01011010010010100" => rgb <= "111000";
					when "01011010010010101" => rgb <= "101000";
					when "01011010010010110" => rgb <= "101000";
					when "01011010010010111" => rgb <= "101000";
					when "01011010010011000" => rgb <= "101000";
					when "01011010010011001" => rgb <= "101000";
					when "01011010010011010" => rgb <= "101000";
					when "01011010010011011" => rgb <= "101000";
					when "01011010010011100" => rgb <= "101000";
					when "01011010010011101" => rgb <= "101000";
					when "01011010010011110" => rgb <= "101000";
					when "01011010010011111" => rgb <= "101000";
					when "01011010010100000" => rgb <= "101000";
					when "01011010010100001" => rgb <= "101000";
					when "01011010010100010" => rgb <= "101000";
					when "01011010010100011" => rgb <= "101000";
					when "01011010010100100" => rgb <= "101000";
					when "01011010010100101" => rgb <= "101000";
					when "01011010010100110" => rgb <= "101000";
					when "01011010010100111" => rgb <= "101000";
					when "01011010010101000" => rgb <= "101000";
					when "01011010010101001" => rgb <= "101000";
					when "01011010010101010" => rgb <= "010000";
					when "01011010010101011" => rgb <= "000000";
					when "01011010010101100" => rgb <= "000000";
					when "01011010010101101" => rgb <= "000000";
					when "01011010010101110" => rgb <= "000000";
					when "01011010010101111" => rgb <= "000000";
					when "01011010010110000" => rgb <= "000000";
					when "01011010010110001" => rgb <= "000000";
					when "01011010010110010" => rgb <= "000000";
					when "01011010010110011" => rgb <= "000000";
					when "01011010010110100" => rgb <= "000000";
					when "01011010010110101" => rgb <= "000000";
					when "01011010010110110" => rgb <= "000000";
					when "01011010010110111" => rgb <= "000000";
					when "01011010010111000" => rgb <= "000000";
					when "01011010010111001" => rgb <= "000000";
					when "01011010010111010" => rgb <= "000000";
					when "01011010010111011" => rgb <= "000000";
					when "01011010010111100" => rgb <= "000000";
					when "01011010010111101" => rgb <= "000000";
					when "01011010010111110" => rgb <= "000000";
					when "01011010010111111" => rgb <= "000000";
					when "01011010011000000" => rgb <= "000000";
					when "01011010011000001" => rgb <= "000000";
					when "01011010011000010" => rgb <= "000000";
					when "01011010011000011" => rgb <= "000000";
					when "01011010011000100" => rgb <= "000000";
					when "01011010011000101" => rgb <= "000000";
					when "01011010011000110" => rgb <= "000000";
					when "01011010011000111" => rgb <= "000000";
					when "01011010011001000" => rgb <= "000000";
					when "01011010011001001" => rgb <= "000000";
					when "01011010011001010" => rgb <= "000000";
					when "01011010011001011" => rgb <= "000000";
					when "01011010011001100" => rgb <= "000000";
					when "01011010011001101" => rgb <= "000000";
					when "01011010011001110" => rgb <= "000000";
					when "01011010011001111" => rgb <= "000000";
					when "01011010011010000" => rgb <= "000000";
					when "01011010011010001" => rgb <= "000000";
					when "01011010011010010" => rgb <= "000000";
					when "01011010011010011" => rgb <= "000000";
					when "01011010011010100" => rgb <= "000000";
					when "01011010011010101" => rgb <= "000000";
					when "01011010011010110" => rgb <= "000000";
					when "01011010011010111" => rgb <= "000000";
					when "01011010011011000" => rgb <= "000000";
					when "01011010011011001" => rgb <= "000000";
					when "01011010011011010" => rgb <= "000000";
					when "01011010011011011" => rgb <= "000000";
					when "01011010011011100" => rgb <= "000000";
					when "01011010011011101" => rgb <= "000000";
					when "01011010011011110" => rgb <= "000000";
					when "01011010011011111" => rgb <= "000000";
					when "01011010011100000" => rgb <= "000000";
					when "01011010011100001" => rgb <= "000000";
					when "01011010011100010" => rgb <= "000000";
					when "01011010011100011" => rgb <= "000000";
					when "01011010011100100" => rgb <= "000000";
					when "01011010011100101" => rgb <= "000000";
					when "01011010011100110" => rgb <= "000000";
					when "01011010011100111" => rgb <= "000000";
					when "01011010011101000" => rgb <= "000000";
					when "01011010011101001" => rgb <= "000000";
					when "01011010011101010" => rgb <= "000000";
					when "01011010011101011" => rgb <= "000000";
					when "01011010011101100" => rgb <= "000000";
					when "01011010011101101" => rgb <= "000000";
					when "01011010011101110" => rgb <= "000000";
					when "01011010011101111" => rgb <= "000000";
					when "01011010011110000" => rgb <= "000000";
					when "01011010011110001" => rgb <= "000000";
					when "01011010011110010" => rgb <= "000000";
					when "01011010011110011" => rgb <= "000000";
					when "01011010011110100" => rgb <= "000000";
					when "01011010011110101" => rgb <= "000000";
					when "01011010011110110" => rgb <= "000000";
					when "01011010011110111" => rgb <= "000000";
					when "01011010011111000" => rgb <= "000000";
					when "01011010011111001" => rgb <= "000000";
					when "01011010011111010" => rgb <= "000000";
					when "01011010011111011" => rgb <= "000000";
					when "01011010011111100" => rgb <= "000000";
					when "01011010011111101" => rgb <= "000000";
					when "01011010011111110" => rgb <= "000000";
					when "01011010011111111" => rgb <= "000000";
					when "01011010100000000" => rgb <= "000000";
					when "01011010100000001" => rgb <= "000000";
					when "01011010100000010" => rgb <= "000000";
					when "01011010100000011" => rgb <= "000000";
					when "01011010100000100" => rgb <= "000000";
					when "01011010100000101" => rgb <= "000000";
					when "01011010100000110" => rgb <= "000000";
					when "01011010100000111" => rgb <= "000000";
					when "01011010100001000" => rgb <= "000000";
					when "01011010100001001" => rgb <= "000000";
					when "01011010100001010" => rgb <= "000000";
					when "01011010100001011" => rgb <= "000000";
					when "01011010100001100" => rgb <= "000000";
					when "01011010100001101" => rgb <= "000000";
					when "01011010100001110" => rgb <= "000000";
					when "01011010100001111" => rgb <= "000000";
					when "01011010100010000" => rgb <= "000000";
					when "01011010100010001" => rgb <= "000000";
					when "01011010100010010" => rgb <= "000000";
					when "01011010100010011" => rgb <= "000000";
					when "01011010100010100" => rgb <= "000000";
					when "01011010100010101" => rgb <= "000000";
					when "01011010100010110" => rgb <= "000000";
					when "01011010100010111" => rgb <= "000000";
					when "01011010100011000" => rgb <= "000000";
					when "01011010100011001" => rgb <= "000000";
					when "01011010100011010" => rgb <= "000000";
					when "01011010100011011" => rgb <= "000000";
					when "01011010100011100" => rgb <= "000000";
					when "01011010100011101" => rgb <= "000000";
					when "01011010100011110" => rgb <= "000000";
					when "01011010100011111" => rgb <= "000000";
					when "01011010100100000" => rgb <= "000000";
					when "01011010100100001" => rgb <= "000000";
					when "01011010100100010" => rgb <= "000000";
					when "01011010100100011" => rgb <= "000000";
					when "01011010100100100" => rgb <= "000000";
					when "01011010100100101" => rgb <= "000000";
					when "01011010100100110" => rgb <= "000000";
					when "01011010100100111" => rgb <= "000000";
					when "01011010100101000" => rgb <= "000000";
					when "01011010100101001" => rgb <= "000000";
					when "01011010100101010" => rgb <= "000000";
					when "01011010100101011" => rgb <= "000000";
					when "01011010100101100" => rgb <= "000000";
					when "01011010100101101" => rgb <= "000000";
					when "01011010100101110" => rgb <= "000000";
					when "01011010100101111" => rgb <= "000000";
					when "01011010100110000" => rgb <= "000000";
					when "01011010100110001" => rgb <= "000000";
					when "01011010100110010" => rgb <= "000000";
					when "01011010100110011" => rgb <= "000000";
					when "01011010100110100" => rgb <= "000000";
					when "01011010100110101" => rgb <= "000000";
					when "01011010100110110" => rgb <= "000000";
					when "01011010100110111" => rgb <= "000000";
					when "01011010100111000" => rgb <= "000000";
					when "01011010100111001" => rgb <= "000000";
					when "01011010100111010" => rgb <= "000000";
					when "01011010100111011" => rgb <= "000000";
					when "01011010100111100" => rgb <= "000000";
					when "01011010100111101" => rgb <= "000000";
					when "01011010100111110" => rgb <= "000000";
					when "01011010100111111" => rgb <= "000000";
					when "01011011000000000" => rgb <= "000000";
					when "01011011000000001" => rgb <= "000000";
					when "01011011000000010" => rgb <= "000000";
					when "01011011000000011" => rgb <= "000000";
					when "01011011000000100" => rgb <= "000000";
					when "01011011000000101" => rgb <= "000000";
					when "01011011000000110" => rgb <= "000000";
					when "01011011000000111" => rgb <= "000000";
					when "01011011000001000" => rgb <= "000000";
					when "01011011000001001" => rgb <= "000000";
					when "01011011000001010" => rgb <= "000000";
					when "01011011000001011" => rgb <= "000000";
					when "01011011000001100" => rgb <= "000000";
					when "01011011000001101" => rgb <= "000000";
					when "01011011000001110" => rgb <= "000000";
					when "01011011000001111" => rgb <= "000000";
					when "01011011000010000" => rgb <= "000000";
					when "01011011000010001" => rgb <= "000000";
					when "01011011000010010" => rgb <= "000000";
					when "01011011000010011" => rgb <= "000000";
					when "01011011000010100" => rgb <= "000000";
					when "01011011000010101" => rgb <= "000000";
					when "01011011000010110" => rgb <= "000000";
					when "01011011000010111" => rgb <= "000000";
					when "01011011000011000" => rgb <= "000000";
					when "01011011000011001" => rgb <= "000000";
					when "01011011000011010" => rgb <= "000000";
					when "01011011000011011" => rgb <= "000000";
					when "01011011000011100" => rgb <= "000000";
					when "01011011000011101" => rgb <= "000000";
					when "01011011000011110" => rgb <= "000000";
					when "01011011000011111" => rgb <= "000000";
					when "01011011000100000" => rgb <= "000000";
					when "01011011000100001" => rgb <= "000000";
					when "01011011000100010" => rgb <= "000000";
					when "01011011000100011" => rgb <= "000000";
					when "01011011000100100" => rgb <= "000000";
					when "01011011000100101" => rgb <= "000000";
					when "01011011000100110" => rgb <= "000000";
					when "01011011000100111" => rgb <= "000000";
					when "01011011000101000" => rgb <= "000000";
					when "01011011000101001" => rgb <= "000000";
					when "01011011000101010" => rgb <= "000000";
					when "01011011000101011" => rgb <= "000000";
					when "01011011000101100" => rgb <= "000000";
					when "01011011000101101" => rgb <= "000000";
					when "01011011000101110" => rgb <= "000000";
					when "01011011000101111" => rgb <= "000000";
					when "01011011000110000" => rgb <= "000000";
					when "01011011000110001" => rgb <= "000000";
					when "01011011000110010" => rgb <= "000000";
					when "01011011000110011" => rgb <= "000000";
					when "01011011000110100" => rgb <= "000000";
					when "01011011000110101" => rgb <= "000000";
					when "01011011000110110" => rgb <= "000000";
					when "01011011000110111" => rgb <= "000000";
					when "01011011000111000" => rgb <= "000000";
					when "01011011000111001" => rgb <= "000000";
					when "01011011000111010" => rgb <= "000000";
					when "01011011000111011" => rgb <= "000000";
					when "01011011000111100" => rgb <= "000000";
					when "01011011000111101" => rgb <= "000000";
					when "01011011000111110" => rgb <= "000000";
					when "01011011000111111" => rgb <= "000000";
					when "01011011001000000" => rgb <= "000000";
					when "01011011001000001" => rgb <= "000000";
					when "01011011001000010" => rgb <= "000000";
					when "01011011001000011" => rgb <= "000000";
					when "01011011001000100" => rgb <= "000000";
					when "01011011001000101" => rgb <= "000000";
					when "01011011001000110" => rgb <= "000000";
					when "01011011001000111" => rgb <= "000000";
					when "01011011001001000" => rgb <= "000000";
					when "01011011001001001" => rgb <= "000000";
					when "01011011001001010" => rgb <= "000000";
					when "01011011001001011" => rgb <= "000000";
					when "01011011001001100" => rgb <= "000000";
					when "01011011001001101" => rgb <= "000000";
					when "01011011001001110" => rgb <= "000000";
					when "01011011001001111" => rgb <= "000000";
					when "01011011001010000" => rgb <= "000000";
					when "01011011001010001" => rgb <= "000000";
					when "01011011001010010" => rgb <= "000000";
					when "01011011001010011" => rgb <= "000000";
					when "01011011001010100" => rgb <= "000000";
					when "01011011001010101" => rgb <= "000000";
					when "01011011001010110" => rgb <= "000000";
					when "01011011001010111" => rgb <= "000000";
					when "01011011001011000" => rgb <= "000000";
					when "01011011001011001" => rgb <= "000000";
					when "01011011001011010" => rgb <= "000000";
					when "01011011001011011" => rgb <= "000000";
					when "01011011001011100" => rgb <= "000000";
					when "01011011001011101" => rgb <= "000000";
					when "01011011001011110" => rgb <= "000000";
					when "01011011001011111" => rgb <= "000000";
					when "01011011001100000" => rgb <= "000000";
					when "01011011001100001" => rgb <= "000000";
					when "01011011001100010" => rgb <= "000000";
					when "01011011001100011" => rgb <= "000000";
					when "01011011001100100" => rgb <= "000000";
					when "01011011001100101" => rgb <= "000000";
					when "01011011001100110" => rgb <= "000000";
					when "01011011001100111" => rgb <= "000000";
					when "01011011001101000" => rgb <= "000000";
					when "01011011001101001" => rgb <= "000000";
					when "01011011001101010" => rgb <= "000000";
					when "01011011001101011" => rgb <= "000000";
					when "01011011001101100" => rgb <= "000000";
					when "01011011001101101" => rgb <= "000000";
					when "01011011001101110" => rgb <= "000000";
					when "01011011001101111" => rgb <= "000000";
					when "01011011001110000" => rgb <= "000000";
					when "01011011001110001" => rgb <= "000000";
					when "01011011001110010" => rgb <= "000000";
					when "01011011001110011" => rgb <= "000000";
					when "01011011001110100" => rgb <= "000000";
					when "01011011001110101" => rgb <= "000000";
					when "01011011001110110" => rgb <= "000000";
					when "01011011001110111" => rgb <= "000000";
					when "01011011001111000" => rgb <= "000000";
					when "01011011001111001" => rgb <= "000000";
					when "01011011001111010" => rgb <= "000000";
					when "01011011001111011" => rgb <= "000000";
					when "01011011001111100" => rgb <= "000000";
					when "01011011001111101" => rgb <= "000000";
					when "01011011001111110" => rgb <= "000000";
					when "01011011001111111" => rgb <= "000000";
					when "01011011010000000" => rgb <= "000000";
					when "01011011010000001" => rgb <= "000000";
					when "01011011010000010" => rgb <= "000000";
					when "01011011010000011" => rgb <= "000000";
					when "01011011010000100" => rgb <= "000000";
					when "01011011010000101" => rgb <= "000000";
					when "01011011010000110" => rgb <= "000000";
					when "01011011010000111" => rgb <= "000000";
					when "01011011010001000" => rgb <= "000000";
					when "01011011010001001" => rgb <= "000000";
					when "01011011010001010" => rgb <= "000000";
					when "01011011010001011" => rgb <= "000000";
					when "01011011010001100" => rgb <= "000000";
					when "01011011010001101" => rgb <= "000000";
					when "01011011010001110" => rgb <= "000000";
					when "01011011010001111" => rgb <= "000000";
					when "01011011010010000" => rgb <= "000000";
					when "01011011010010001" => rgb <= "000000";
					when "01011011010010010" => rgb <= "000000";
					when "01011011010010011" => rgb <= "010100";
					when "01011011010010100" => rgb <= "111000";
					when "01011011010010101" => rgb <= "101000";
					when "01011011010010110" => rgb <= "101000";
					when "01011011010010111" => rgb <= "101000";
					when "01011011010011000" => rgb <= "101000";
					when "01011011010011001" => rgb <= "101000";
					when "01011011010011010" => rgb <= "101000";
					when "01011011010011011" => rgb <= "101000";
					when "01011011010011100" => rgb <= "101000";
					when "01011011010011101" => rgb <= "101000";
					when "01011011010011110" => rgb <= "101000";
					when "01011011010011111" => rgb <= "101000";
					when "01011011010100000" => rgb <= "101000";
					when "01011011010100001" => rgb <= "101000";
					when "01011011010100010" => rgb <= "101000";
					when "01011011010100011" => rgb <= "101000";
					when "01011011010100100" => rgb <= "101000";
					when "01011011010100101" => rgb <= "101000";
					when "01011011010100110" => rgb <= "101000";
					when "01011011010100111" => rgb <= "101000";
					when "01011011010101000" => rgb <= "101000";
					when "01011011010101001" => rgb <= "101000";
					when "01011011010101010" => rgb <= "010000";
					when "01011011010101011" => rgb <= "000000";
					when "01011011010101100" => rgb <= "000000";
					when "01011011010101101" => rgb <= "000000";
					when "01011011010101110" => rgb <= "000000";
					when "01011011010101111" => rgb <= "000000";
					when "01011011010110000" => rgb <= "000000";
					when "01011011010110001" => rgb <= "000000";
					when "01011011010110010" => rgb <= "000000";
					when "01011011010110011" => rgb <= "000000";
					when "01011011010110100" => rgb <= "000000";
					when "01011011010110101" => rgb <= "000000";
					when "01011011010110110" => rgb <= "000000";
					when "01011011010110111" => rgb <= "000000";
					when "01011011010111000" => rgb <= "000000";
					when "01011011010111001" => rgb <= "000000";
					when "01011011010111010" => rgb <= "000000";
					when "01011011010111011" => rgb <= "000000";
					when "01011011010111100" => rgb <= "000000";
					when "01011011010111101" => rgb <= "000000";
					when "01011011010111110" => rgb <= "000000";
					when "01011011010111111" => rgb <= "000000";
					when "01011011011000000" => rgb <= "000000";
					when "01011011011000001" => rgb <= "000000";
					when "01011011011000010" => rgb <= "000000";
					when "01011011011000011" => rgb <= "000000";
					when "01011011011000100" => rgb <= "000000";
					when "01011011011000101" => rgb <= "000000";
					when "01011011011000110" => rgb <= "000000";
					when "01011011011000111" => rgb <= "000000";
					when "01011011011001000" => rgb <= "000000";
					when "01011011011001001" => rgb <= "000000";
					when "01011011011001010" => rgb <= "000000";
					when "01011011011001011" => rgb <= "000000";
					when "01011011011001100" => rgb <= "000000";
					when "01011011011001101" => rgb <= "000000";
					when "01011011011001110" => rgb <= "000000";
					when "01011011011001111" => rgb <= "000000";
					when "01011011011010000" => rgb <= "000000";
					when "01011011011010001" => rgb <= "000000";
					when "01011011011010010" => rgb <= "000000";
					when "01011011011010011" => rgb <= "000000";
					when "01011011011010100" => rgb <= "000000";
					when "01011011011010101" => rgb <= "000000";
					when "01011011011010110" => rgb <= "000000";
					when "01011011011010111" => rgb <= "000000";
					when "01011011011011000" => rgb <= "000000";
					when "01011011011011001" => rgb <= "000000";
					when "01011011011011010" => rgb <= "000000";
					when "01011011011011011" => rgb <= "000000";
					when "01011011011011100" => rgb <= "000000";
					when "01011011011011101" => rgb <= "000000";
					when "01011011011011110" => rgb <= "000000";
					when "01011011011011111" => rgb <= "000000";
					when "01011011011100000" => rgb <= "000000";
					when "01011011011100001" => rgb <= "000000";
					when "01011011011100010" => rgb <= "000000";
					when "01011011011100011" => rgb <= "000000";
					when "01011011011100100" => rgb <= "000000";
					when "01011011011100101" => rgb <= "000000";
					when "01011011011100110" => rgb <= "000000";
					when "01011011011100111" => rgb <= "000000";
					when "01011011011101000" => rgb <= "000000";
					when "01011011011101001" => rgb <= "000000";
					when "01011011011101010" => rgb <= "000000";
					when "01011011011101011" => rgb <= "000000";
					when "01011011011101100" => rgb <= "000000";
					when "01011011011101101" => rgb <= "000000";
					when "01011011011101110" => rgb <= "000000";
					when "01011011011101111" => rgb <= "000000";
					when "01011011011110000" => rgb <= "000000";
					when "01011011011110001" => rgb <= "000000";
					when "01011011011110010" => rgb <= "000000";
					when "01011011011110011" => rgb <= "000000";
					when "01011011011110100" => rgb <= "000000";
					when "01011011011110101" => rgb <= "000000";
					when "01011011011110110" => rgb <= "000000";
					when "01011011011110111" => rgb <= "000000";
					when "01011011011111000" => rgb <= "000000";
					when "01011011011111001" => rgb <= "000000";
					when "01011011011111010" => rgb <= "000000";
					when "01011011011111011" => rgb <= "000000";
					when "01011011011111100" => rgb <= "000000";
					when "01011011011111101" => rgb <= "000000";
					when "01011011011111110" => rgb <= "000000";
					when "01011011011111111" => rgb <= "000000";
					when "01011011100000000" => rgb <= "000000";
					when "01011011100000001" => rgb <= "000000";
					when "01011011100000010" => rgb <= "000000";
					when "01011011100000011" => rgb <= "000000";
					when "01011011100000100" => rgb <= "000000";
					when "01011011100000101" => rgb <= "000000";
					when "01011011100000110" => rgb <= "000000";
					when "01011011100000111" => rgb <= "000000";
					when "01011011100001000" => rgb <= "000000";
					when "01011011100001001" => rgb <= "000000";
					when "01011011100001010" => rgb <= "000000";
					when "01011011100001011" => rgb <= "000000";
					when "01011011100001100" => rgb <= "000000";
					when "01011011100001101" => rgb <= "000000";
					when "01011011100001110" => rgb <= "000000";
					when "01011011100001111" => rgb <= "000000";
					when "01011011100010000" => rgb <= "000000";
					when "01011011100010001" => rgb <= "000000";
					when "01011011100010010" => rgb <= "000000";
					when "01011011100010011" => rgb <= "000000";
					when "01011011100010100" => rgb <= "000000";
					when "01011011100010101" => rgb <= "000000";
					when "01011011100010110" => rgb <= "000000";
					when "01011011100010111" => rgb <= "000000";
					when "01011011100011000" => rgb <= "000000";
					when "01011011100011001" => rgb <= "000000";
					when "01011011100011010" => rgb <= "000000";
					when "01011011100011011" => rgb <= "000000";
					when "01011011100011100" => rgb <= "000000";
					when "01011011100011101" => rgb <= "000000";
					when "01011011100011110" => rgb <= "000000";
					when "01011011100011111" => rgb <= "000000";
					when "01011011100100000" => rgb <= "000000";
					when "01011011100100001" => rgb <= "000000";
					when "01011011100100010" => rgb <= "000000";
					when "01011011100100011" => rgb <= "000000";
					when "01011011100100100" => rgb <= "000000";
					when "01011011100100101" => rgb <= "000000";
					when "01011011100100110" => rgb <= "000000";
					when "01011011100100111" => rgb <= "000000";
					when "01011011100101000" => rgb <= "000000";
					when "01011011100101001" => rgb <= "000000";
					when "01011011100101010" => rgb <= "000000";
					when "01011011100101011" => rgb <= "000000";
					when "01011011100101100" => rgb <= "000000";
					when "01011011100101101" => rgb <= "000000";
					when "01011011100101110" => rgb <= "000000";
					when "01011011100101111" => rgb <= "000000";
					when "01011011100110000" => rgb <= "000000";
					when "01011011100110001" => rgb <= "000000";
					when "01011011100110010" => rgb <= "000000";
					when "01011011100110011" => rgb <= "000000";
					when "01011011100110100" => rgb <= "000000";
					when "01011011100110101" => rgb <= "000000";
					when "01011011100110110" => rgb <= "000000";
					when "01011011100110111" => rgb <= "000000";
					when "01011011100111000" => rgb <= "000000";
					when "01011011100111001" => rgb <= "000000";
					when "01011011100111010" => rgb <= "000000";
					when "01011011100111011" => rgb <= "000000";
					when "01011011100111100" => rgb <= "000000";
					when "01011011100111101" => rgb <= "000000";
					when "01011011100111110" => rgb <= "000000";
					when "01011011100111111" => rgb <= "000000";
					when "01011100000000000" => rgb <= "000000";
					when "01011100000000001" => rgb <= "000000";
					when "01011100000000010" => rgb <= "000000";
					when "01011100000000011" => rgb <= "000000";
					when "01011100000000100" => rgb <= "000000";
					when "01011100000000101" => rgb <= "000000";
					when "01011100000000110" => rgb <= "000000";
					when "01011100000000111" => rgb <= "000000";
					when "01011100000001000" => rgb <= "000000";
					when "01011100000001001" => rgb <= "000000";
					when "01011100000001010" => rgb <= "000000";
					when "01011100000001011" => rgb <= "000000";
					when "01011100000001100" => rgb <= "000000";
					when "01011100000001101" => rgb <= "000000";
					when "01011100000001110" => rgb <= "000000";
					when "01011100000001111" => rgb <= "000000";
					when "01011100000010000" => rgb <= "000000";
					when "01011100000010001" => rgb <= "000000";
					when "01011100000010010" => rgb <= "000000";
					when "01011100000010011" => rgb <= "000000";
					when "01011100000010100" => rgb <= "000000";
					when "01011100000010101" => rgb <= "000000";
					when "01011100000010110" => rgb <= "000000";
					when "01011100000010111" => rgb <= "000000";
					when "01011100000011000" => rgb <= "000000";
					when "01011100000011001" => rgb <= "000000";
					when "01011100000011010" => rgb <= "000000";
					when "01011100000011011" => rgb <= "000000";
					when "01011100000011100" => rgb <= "000000";
					when "01011100000011101" => rgb <= "000000";
					when "01011100000011110" => rgb <= "000000";
					when "01011100000011111" => rgb <= "000000";
					when "01011100000100000" => rgb <= "000000";
					when "01011100000100001" => rgb <= "000000";
					when "01011100000100010" => rgb <= "000000";
					when "01011100000100011" => rgb <= "000000";
					when "01011100000100100" => rgb <= "000000";
					when "01011100000100101" => rgb <= "000000";
					when "01011100000100110" => rgb <= "000000";
					when "01011100000100111" => rgb <= "000000";
					when "01011100000101000" => rgb <= "000000";
					when "01011100000101001" => rgb <= "000000";
					when "01011100000101010" => rgb <= "000000";
					when "01011100000101011" => rgb <= "000000";
					when "01011100000101100" => rgb <= "000000";
					when "01011100000101101" => rgb <= "000000";
					when "01011100000101110" => rgb <= "000000";
					when "01011100000101111" => rgb <= "000000";
					when "01011100000110000" => rgb <= "000000";
					when "01011100000110001" => rgb <= "000000";
					when "01011100000110010" => rgb <= "000000";
					when "01011100000110011" => rgb <= "000000";
					when "01011100000110100" => rgb <= "000000";
					when "01011100000110101" => rgb <= "000000";
					when "01011100000110110" => rgb <= "000000";
					when "01011100000110111" => rgb <= "000000";
					when "01011100000111000" => rgb <= "000000";
					when "01011100000111001" => rgb <= "000000";
					when "01011100000111010" => rgb <= "000000";
					when "01011100000111011" => rgb <= "000000";
					when "01011100000111100" => rgb <= "000000";
					when "01011100000111101" => rgb <= "000000";
					when "01011100000111110" => rgb <= "000000";
					when "01011100000111111" => rgb <= "000000";
					when "01011100001000000" => rgb <= "000000";
					when "01011100001000001" => rgb <= "000000";
					when "01011100001000010" => rgb <= "000000";
					when "01011100001000011" => rgb <= "000000";
					when "01011100001000100" => rgb <= "000000";
					when "01011100001000101" => rgb <= "000000";
					when "01011100001000110" => rgb <= "000000";
					when "01011100001000111" => rgb <= "000000";
					when "01011100001001000" => rgb <= "000000";
					when "01011100001001001" => rgb <= "000000";
					when "01011100001001010" => rgb <= "000000";
					when "01011100001001011" => rgb <= "000000";
					when "01011100001001100" => rgb <= "000000";
					when "01011100001001101" => rgb <= "000000";
					when "01011100001001110" => rgb <= "000000";
					when "01011100001001111" => rgb <= "000000";
					when "01011100001010000" => rgb <= "000000";
					when "01011100001010001" => rgb <= "000000";
					when "01011100001010010" => rgb <= "000000";
					when "01011100001010011" => rgb <= "000000";
					when "01011100001010100" => rgb <= "000000";
					when "01011100001010101" => rgb <= "000000";
					when "01011100001010110" => rgb <= "000000";
					when "01011100001010111" => rgb <= "000000";
					when "01011100001011000" => rgb <= "000000";
					when "01011100001011001" => rgb <= "000000";
					when "01011100001011010" => rgb <= "000000";
					when "01011100001011011" => rgb <= "000000";
					when "01011100001011100" => rgb <= "000000";
					when "01011100001011101" => rgb <= "000000";
					when "01011100001011110" => rgb <= "000000";
					when "01011100001011111" => rgb <= "000000";
					when "01011100001100000" => rgb <= "000000";
					when "01011100001100001" => rgb <= "000000";
					when "01011100001100010" => rgb <= "000000";
					when "01011100001100011" => rgb <= "000000";
					when "01011100001100100" => rgb <= "000000";
					when "01011100001100101" => rgb <= "000000";
					when "01011100001100110" => rgb <= "000000";
					when "01011100001100111" => rgb <= "000000";
					when "01011100001101000" => rgb <= "000000";
					when "01011100001101001" => rgb <= "000000";
					when "01011100001101010" => rgb <= "000000";
					when "01011100001101011" => rgb <= "000000";
					when "01011100001101100" => rgb <= "000000";
					when "01011100001101101" => rgb <= "000000";
					when "01011100001101110" => rgb <= "000000";
					when "01011100001101111" => rgb <= "000000";
					when "01011100001110000" => rgb <= "000000";
					when "01011100001110001" => rgb <= "000000";
					when "01011100001110010" => rgb <= "000000";
					when "01011100001110011" => rgb <= "000000";
					when "01011100001110100" => rgb <= "000000";
					when "01011100001110101" => rgb <= "000000";
					when "01011100001110110" => rgb <= "000000";
					when "01011100001110111" => rgb <= "000000";
					when "01011100001111000" => rgb <= "000000";
					when "01011100001111001" => rgb <= "000000";
					when "01011100001111010" => rgb <= "000000";
					when "01011100001111011" => rgb <= "000000";
					when "01011100001111100" => rgb <= "000000";
					when "01011100001111101" => rgb <= "000000";
					when "01011100001111110" => rgb <= "000000";
					when "01011100001111111" => rgb <= "000000";
					when "01011100010000000" => rgb <= "000000";
					when "01011100010000001" => rgb <= "000000";
					when "01011100010000010" => rgb <= "000000";
					when "01011100010000011" => rgb <= "000000";
					when "01011100010000100" => rgb <= "000000";
					when "01011100010000101" => rgb <= "000000";
					when "01011100010000110" => rgb <= "000000";
					when "01011100010000111" => rgb <= "000000";
					when "01011100010001000" => rgb <= "000000";
					when "01011100010001001" => rgb <= "000000";
					when "01011100010001010" => rgb <= "000000";
					when "01011100010001011" => rgb <= "000000";
					when "01011100010001100" => rgb <= "000000";
					when "01011100010001101" => rgb <= "000000";
					when "01011100010001110" => rgb <= "000000";
					when "01011100010001111" => rgb <= "000000";
					when "01011100010010000" => rgb <= "000000";
					when "01011100010010001" => rgb <= "000000";
					when "01011100010010010" => rgb <= "000000";
					when "01011100010010011" => rgb <= "010100";
					when "01011100010010100" => rgb <= "111000";
					when "01011100010010101" => rgb <= "101000";
					when "01011100010010110" => rgb <= "101000";
					when "01011100010010111" => rgb <= "101000";
					when "01011100010011000" => rgb <= "101000";
					when "01011100010011001" => rgb <= "101000";
					when "01011100010011010" => rgb <= "101000";
					when "01011100010011011" => rgb <= "101000";
					when "01011100010011100" => rgb <= "101000";
					when "01011100010011101" => rgb <= "101000";
					when "01011100010011110" => rgb <= "101000";
					when "01011100010011111" => rgb <= "101000";
					when "01011100010100000" => rgb <= "101000";
					when "01011100010100001" => rgb <= "101000";
					when "01011100010100010" => rgb <= "101000";
					when "01011100010100011" => rgb <= "101000";
					when "01011100010100100" => rgb <= "101000";
					when "01011100010100101" => rgb <= "101000";
					when "01011100010100110" => rgb <= "101000";
					when "01011100010100111" => rgb <= "101000";
					when "01011100010101000" => rgb <= "101000";
					when "01011100010101001" => rgb <= "101000";
					when "01011100010101010" => rgb <= "010000";
					when "01011100010101011" => rgb <= "000000";
					when "01011100010101100" => rgb <= "000000";
					when "01011100010101101" => rgb <= "000000";
					when "01011100010101110" => rgb <= "000000";
					when "01011100010101111" => rgb <= "000000";
					when "01011100010110000" => rgb <= "000000";
					when "01011100010110001" => rgb <= "000000";
					when "01011100010110010" => rgb <= "000000";
					when "01011100010110011" => rgb <= "000000";
					when "01011100010110100" => rgb <= "000000";
					when "01011100010110101" => rgb <= "000000";
					when "01011100010110110" => rgb <= "000000";
					when "01011100010110111" => rgb <= "000000";
					when "01011100010111000" => rgb <= "000000";
					when "01011100010111001" => rgb <= "000000";
					when "01011100010111010" => rgb <= "000000";
					when "01011100010111011" => rgb <= "000000";
					when "01011100010111100" => rgb <= "000000";
					when "01011100010111101" => rgb <= "000000";
					when "01011100010111110" => rgb <= "000000";
					when "01011100010111111" => rgb <= "000000";
					when "01011100011000000" => rgb <= "000000";
					when "01011100011000001" => rgb <= "000000";
					when "01011100011000010" => rgb <= "000000";
					when "01011100011000011" => rgb <= "000000";
					when "01011100011000100" => rgb <= "000000";
					when "01011100011000101" => rgb <= "000000";
					when "01011100011000110" => rgb <= "000000";
					when "01011100011000111" => rgb <= "000000";
					when "01011100011001000" => rgb <= "000000";
					when "01011100011001001" => rgb <= "000000";
					when "01011100011001010" => rgb <= "000000";
					when "01011100011001011" => rgb <= "000000";
					when "01011100011001100" => rgb <= "000000";
					when "01011100011001101" => rgb <= "000000";
					when "01011100011001110" => rgb <= "000000";
					when "01011100011001111" => rgb <= "000000";
					when "01011100011010000" => rgb <= "000000";
					when "01011100011010001" => rgb <= "000000";
					when "01011100011010010" => rgb <= "000000";
					when "01011100011010011" => rgb <= "000000";
					when "01011100011010100" => rgb <= "000000";
					when "01011100011010101" => rgb <= "000000";
					when "01011100011010110" => rgb <= "000000";
					when "01011100011010111" => rgb <= "000000";
					when "01011100011011000" => rgb <= "000000";
					when "01011100011011001" => rgb <= "000000";
					when "01011100011011010" => rgb <= "000000";
					when "01011100011011011" => rgb <= "000000";
					when "01011100011011100" => rgb <= "000000";
					when "01011100011011101" => rgb <= "000000";
					when "01011100011011110" => rgb <= "000000";
					when "01011100011011111" => rgb <= "000000";
					when "01011100011100000" => rgb <= "000000";
					when "01011100011100001" => rgb <= "000000";
					when "01011100011100010" => rgb <= "000000";
					when "01011100011100011" => rgb <= "000000";
					when "01011100011100100" => rgb <= "000000";
					when "01011100011100101" => rgb <= "000000";
					when "01011100011100110" => rgb <= "000000";
					when "01011100011100111" => rgb <= "000000";
					when "01011100011101000" => rgb <= "000000";
					when "01011100011101001" => rgb <= "000000";
					when "01011100011101010" => rgb <= "000000";
					when "01011100011101011" => rgb <= "000000";
					when "01011100011101100" => rgb <= "000000";
					when "01011100011101101" => rgb <= "000000";
					when "01011100011101110" => rgb <= "000000";
					when "01011100011101111" => rgb <= "000000";
					when "01011100011110000" => rgb <= "000000";
					when "01011100011110001" => rgb <= "000000";
					when "01011100011110010" => rgb <= "000000";
					when "01011100011110011" => rgb <= "000000";
					when "01011100011110100" => rgb <= "000000";
					when "01011100011110101" => rgb <= "000000";
					when "01011100011110110" => rgb <= "000000";
					when "01011100011110111" => rgb <= "000000";
					when "01011100011111000" => rgb <= "000000";
					when "01011100011111001" => rgb <= "000000";
					when "01011100011111010" => rgb <= "000000";
					when "01011100011111011" => rgb <= "000000";
					when "01011100011111100" => rgb <= "000000";
					when "01011100011111101" => rgb <= "000000";
					when "01011100011111110" => rgb <= "000000";
					when "01011100011111111" => rgb <= "000000";
					when "01011100100000000" => rgb <= "000000";
					when "01011100100000001" => rgb <= "000000";
					when "01011100100000010" => rgb <= "000000";
					when "01011100100000011" => rgb <= "000000";
					when "01011100100000100" => rgb <= "000000";
					when "01011100100000101" => rgb <= "000000";
					when "01011100100000110" => rgb <= "000000";
					when "01011100100000111" => rgb <= "000000";
					when "01011100100001000" => rgb <= "000000";
					when "01011100100001001" => rgb <= "000000";
					when "01011100100001010" => rgb <= "000000";
					when "01011100100001011" => rgb <= "000000";
					when "01011100100001100" => rgb <= "000000";
					when "01011100100001101" => rgb <= "000000";
					when "01011100100001110" => rgb <= "000000";
					when "01011100100001111" => rgb <= "000000";
					when "01011100100010000" => rgb <= "000000";
					when "01011100100010001" => rgb <= "000000";
					when "01011100100010010" => rgb <= "000000";
					when "01011100100010011" => rgb <= "000000";
					when "01011100100010100" => rgb <= "000000";
					when "01011100100010101" => rgb <= "000000";
					when "01011100100010110" => rgb <= "000000";
					when "01011100100010111" => rgb <= "000000";
					when "01011100100011000" => rgb <= "000000";
					when "01011100100011001" => rgb <= "000000";
					when "01011100100011010" => rgb <= "000000";
					when "01011100100011011" => rgb <= "000000";
					when "01011100100011100" => rgb <= "000000";
					when "01011100100011101" => rgb <= "000000";
					when "01011100100011110" => rgb <= "000000";
					when "01011100100011111" => rgb <= "000000";
					when "01011100100100000" => rgb <= "000000";
					when "01011100100100001" => rgb <= "000000";
					when "01011100100100010" => rgb <= "000000";
					when "01011100100100011" => rgb <= "000000";
					when "01011100100100100" => rgb <= "000000";
					when "01011100100100101" => rgb <= "000000";
					when "01011100100100110" => rgb <= "000000";
					when "01011100100100111" => rgb <= "000000";
					when "01011100100101000" => rgb <= "000000";
					when "01011100100101001" => rgb <= "000000";
					when "01011100100101010" => rgb <= "000000";
					when "01011100100101011" => rgb <= "000000";
					when "01011100100101100" => rgb <= "000000";
					when "01011100100101101" => rgb <= "000000";
					when "01011100100101110" => rgb <= "000000";
					when "01011100100101111" => rgb <= "000000";
					when "01011100100110000" => rgb <= "000000";
					when "01011100100110001" => rgb <= "000000";
					when "01011100100110010" => rgb <= "000000";
					when "01011100100110011" => rgb <= "000000";
					when "01011100100110100" => rgb <= "000000";
					when "01011100100110101" => rgb <= "000000";
					when "01011100100110110" => rgb <= "000000";
					when "01011100100110111" => rgb <= "000000";
					when "01011100100111000" => rgb <= "000000";
					when "01011100100111001" => rgb <= "000000";
					when "01011100100111010" => rgb <= "000000";
					when "01011100100111011" => rgb <= "000000";
					when "01011100100111100" => rgb <= "000000";
					when "01011100100111101" => rgb <= "000000";
					when "01011100100111110" => rgb <= "000000";
					when "01011100100111111" => rgb <= "000000";
					when "01011101000000000" => rgb <= "000000";
					when "01011101000000001" => rgb <= "000000";
					when "01011101000000010" => rgb <= "000000";
					when "01011101000000011" => rgb <= "000000";
					when "01011101000000100" => rgb <= "000000";
					when "01011101000000101" => rgb <= "000000";
					when "01011101000000110" => rgb <= "000000";
					when "01011101000000111" => rgb <= "000000";
					when "01011101000001000" => rgb <= "000000";
					when "01011101000001001" => rgb <= "000000";
					when "01011101000001010" => rgb <= "000000";
					when "01011101000001011" => rgb <= "000000";
					when "01011101000001100" => rgb <= "000000";
					when "01011101000001101" => rgb <= "000000";
					when "01011101000001110" => rgb <= "000000";
					when "01011101000001111" => rgb <= "000000";
					when "01011101000010000" => rgb <= "000000";
					when "01011101000010001" => rgb <= "000000";
					when "01011101000010010" => rgb <= "000000";
					when "01011101000010011" => rgb <= "000000";
					when "01011101000010100" => rgb <= "000000";
					when "01011101000010101" => rgb <= "000000";
					when "01011101000010110" => rgb <= "000000";
					when "01011101000010111" => rgb <= "000000";
					when "01011101000011000" => rgb <= "000000";
					when "01011101000011001" => rgb <= "000000";
					when "01011101000011010" => rgb <= "000000";
					when "01011101000011011" => rgb <= "000000";
					when "01011101000011100" => rgb <= "000000";
					when "01011101000011101" => rgb <= "000000";
					when "01011101000011110" => rgb <= "000000";
					when "01011101000011111" => rgb <= "000000";
					when "01011101000100000" => rgb <= "000000";
					when "01011101000100001" => rgb <= "000000";
					when "01011101000100010" => rgb <= "000000";
					when "01011101000100011" => rgb <= "000000";
					when "01011101000100100" => rgb <= "000000";
					when "01011101000100101" => rgb <= "000000";
					when "01011101000100110" => rgb <= "000000";
					when "01011101000100111" => rgb <= "000000";
					when "01011101000101000" => rgb <= "000000";
					when "01011101000101001" => rgb <= "000000";
					when "01011101000101010" => rgb <= "000000";
					when "01011101000101011" => rgb <= "000000";
					when "01011101000101100" => rgb <= "000000";
					when "01011101000101101" => rgb <= "000000";
					when "01011101000101110" => rgb <= "000000";
					when "01011101000101111" => rgb <= "000000";
					when "01011101000110000" => rgb <= "000000";
					when "01011101000110001" => rgb <= "000000";
					when "01011101000110010" => rgb <= "000000";
					when "01011101000110011" => rgb <= "000000";
					when "01011101000110100" => rgb <= "000000";
					when "01011101000110101" => rgb <= "000000";
					when "01011101000110110" => rgb <= "000000";
					when "01011101000110111" => rgb <= "000000";
					when "01011101000111000" => rgb <= "000000";
					when "01011101000111001" => rgb <= "000000";
					when "01011101000111010" => rgb <= "000000";
					when "01011101000111011" => rgb <= "000000";
					when "01011101000111100" => rgb <= "000000";
					when "01011101000111101" => rgb <= "000000";
					when "01011101000111110" => rgb <= "000000";
					when "01011101000111111" => rgb <= "000000";
					when "01011101001000000" => rgb <= "000000";
					when "01011101001000001" => rgb <= "000000";
					when "01011101001000010" => rgb <= "000000";
					when "01011101001000011" => rgb <= "000000";
					when "01011101001000100" => rgb <= "000000";
					when "01011101001000101" => rgb <= "000000";
					when "01011101001000110" => rgb <= "000000";
					when "01011101001000111" => rgb <= "000000";
					when "01011101001001000" => rgb <= "000000";
					when "01011101001001001" => rgb <= "000000";
					when "01011101001001010" => rgb <= "000000";
					when "01011101001001011" => rgb <= "000000";
					when "01011101001001100" => rgb <= "000000";
					when "01011101001001101" => rgb <= "000000";
					when "01011101001001110" => rgb <= "000000";
					when "01011101001001111" => rgb <= "000000";
					when "01011101001010000" => rgb <= "000000";
					when "01011101001010001" => rgb <= "000000";
					when "01011101001010010" => rgb <= "000000";
					when "01011101001010011" => rgb <= "000000";
					when "01011101001010100" => rgb <= "000000";
					when "01011101001010101" => rgb <= "000000";
					when "01011101001010110" => rgb <= "000000";
					when "01011101001010111" => rgb <= "000000";
					when "01011101001011000" => rgb <= "000000";
					when "01011101001011001" => rgb <= "000000";
					when "01011101001011010" => rgb <= "000000";
					when "01011101001011011" => rgb <= "000000";
					when "01011101001011100" => rgb <= "000000";
					when "01011101001011101" => rgb <= "000000";
					when "01011101001011110" => rgb <= "000000";
					when "01011101001011111" => rgb <= "000000";
					when "01011101001100000" => rgb <= "000000";
					when "01011101001100001" => rgb <= "000000";
					when "01011101001100010" => rgb <= "000000";
					when "01011101001100011" => rgb <= "000000";
					when "01011101001100100" => rgb <= "000000";
					when "01011101001100101" => rgb <= "000000";
					when "01011101001100110" => rgb <= "000000";
					when "01011101001100111" => rgb <= "000000";
					when "01011101001101000" => rgb <= "000000";
					when "01011101001101001" => rgb <= "000000";
					when "01011101001101010" => rgb <= "000000";
					when "01011101001101011" => rgb <= "000000";
					when "01011101001101100" => rgb <= "000000";
					when "01011101001101101" => rgb <= "000000";
					when "01011101001101110" => rgb <= "000000";
					when "01011101001101111" => rgb <= "000000";
					when "01011101001110000" => rgb <= "000000";
					when "01011101001110001" => rgb <= "000000";
					when "01011101001110010" => rgb <= "000000";
					when "01011101001110011" => rgb <= "000000";
					when "01011101001110100" => rgb <= "000000";
					when "01011101001110101" => rgb <= "000000";
					when "01011101001110110" => rgb <= "000000";
					when "01011101001110111" => rgb <= "000000";
					when "01011101001111000" => rgb <= "000000";
					when "01011101001111001" => rgb <= "000000";
					when "01011101001111010" => rgb <= "000000";
					when "01011101001111011" => rgb <= "000000";
					when "01011101001111100" => rgb <= "000000";
					when "01011101001111101" => rgb <= "000000";
					when "01011101001111110" => rgb <= "000000";
					when "01011101001111111" => rgb <= "000000";
					when "01011101010000000" => rgb <= "000000";
					when "01011101010000001" => rgb <= "000000";
					when "01011101010000010" => rgb <= "000000";
					when "01011101010000011" => rgb <= "000000";
					when "01011101010000100" => rgb <= "000000";
					when "01011101010000101" => rgb <= "000000";
					when "01011101010000110" => rgb <= "000000";
					when "01011101010000111" => rgb <= "000000";
					when "01011101010001000" => rgb <= "000000";
					when "01011101010001001" => rgb <= "000000";
					when "01011101010001010" => rgb <= "000000";
					when "01011101010001011" => rgb <= "000000";
					when "01011101010001100" => rgb <= "000000";
					when "01011101010001101" => rgb <= "000000";
					when "01011101010001110" => rgb <= "000000";
					when "01011101010001111" => rgb <= "000000";
					when "01011101010010000" => rgb <= "000000";
					when "01011101010010001" => rgb <= "000000";
					when "01011101010010010" => rgb <= "000000";
					when "01011101010010011" => rgb <= "010100";
					when "01011101010010100" => rgb <= "111000";
					when "01011101010010101" => rgb <= "101000";
					when "01011101010010110" => rgb <= "101000";
					when "01011101010010111" => rgb <= "101000";
					when "01011101010011000" => rgb <= "101000";
					when "01011101010011001" => rgb <= "101000";
					when "01011101010011010" => rgb <= "101000";
					when "01011101010011011" => rgb <= "101000";
					when "01011101010011100" => rgb <= "101000";
					when "01011101010011101" => rgb <= "101000";
					when "01011101010011110" => rgb <= "101000";
					when "01011101010011111" => rgb <= "101000";
					when "01011101010100000" => rgb <= "101000";
					when "01011101010100001" => rgb <= "101000";
					when "01011101010100010" => rgb <= "101000";
					when "01011101010100011" => rgb <= "101000";
					when "01011101010100100" => rgb <= "101000";
					when "01011101010100101" => rgb <= "101000";
					when "01011101010100110" => rgb <= "101000";
					when "01011101010100111" => rgb <= "101000";
					when "01011101010101000" => rgb <= "101000";
					when "01011101010101001" => rgb <= "101000";
					when "01011101010101010" => rgb <= "010000";
					when "01011101010101011" => rgb <= "000000";
					when "01011101010101100" => rgb <= "000000";
					when "01011101010101101" => rgb <= "000000";
					when "01011101010101110" => rgb <= "000000";
					when "01011101010101111" => rgb <= "000000";
					when "01011101010110000" => rgb <= "000000";
					when "01011101010110001" => rgb <= "000000";
					when "01011101010110010" => rgb <= "000000";
					when "01011101010110011" => rgb <= "000000";
					when "01011101010110100" => rgb <= "000000";
					when "01011101010110101" => rgb <= "000000";
					when "01011101010110110" => rgb <= "000000";
					when "01011101010110111" => rgb <= "000000";
					when "01011101010111000" => rgb <= "000000";
					when "01011101010111001" => rgb <= "000000";
					when "01011101010111010" => rgb <= "000000";
					when "01011101010111011" => rgb <= "000000";
					when "01011101010111100" => rgb <= "000000";
					when "01011101010111101" => rgb <= "000000";
					when "01011101010111110" => rgb <= "000000";
					when "01011101010111111" => rgb <= "000000";
					when "01011101011000000" => rgb <= "000000";
					when "01011101011000001" => rgb <= "000000";
					when "01011101011000010" => rgb <= "000000";
					when "01011101011000011" => rgb <= "000000";
					when "01011101011000100" => rgb <= "000000";
					when "01011101011000101" => rgb <= "000000";
					when "01011101011000110" => rgb <= "000000";
					when "01011101011000111" => rgb <= "000000";
					when "01011101011001000" => rgb <= "000000";
					when "01011101011001001" => rgb <= "000000";
					when "01011101011001010" => rgb <= "000000";
					when "01011101011001011" => rgb <= "000000";
					when "01011101011001100" => rgb <= "000000";
					when "01011101011001101" => rgb <= "000000";
					when "01011101011001110" => rgb <= "000000";
					when "01011101011001111" => rgb <= "000000";
					when "01011101011010000" => rgb <= "000000";
					when "01011101011010001" => rgb <= "000000";
					when "01011101011010010" => rgb <= "000000";
					when "01011101011010011" => rgb <= "000000";
					when "01011101011010100" => rgb <= "000000";
					when "01011101011010101" => rgb <= "000000";
					when "01011101011010110" => rgb <= "000000";
					when "01011101011010111" => rgb <= "000000";
					when "01011101011011000" => rgb <= "000000";
					when "01011101011011001" => rgb <= "000000";
					when "01011101011011010" => rgb <= "000000";
					when "01011101011011011" => rgb <= "000000";
					when "01011101011011100" => rgb <= "000000";
					when "01011101011011101" => rgb <= "000000";
					when "01011101011011110" => rgb <= "000000";
					when "01011101011011111" => rgb <= "000000";
					when "01011101011100000" => rgb <= "000000";
					when "01011101011100001" => rgb <= "000000";
					when "01011101011100010" => rgb <= "000000";
					when "01011101011100011" => rgb <= "000000";
					when "01011101011100100" => rgb <= "000000";
					when "01011101011100101" => rgb <= "000000";
					when "01011101011100110" => rgb <= "000000";
					when "01011101011100111" => rgb <= "000000";
					when "01011101011101000" => rgb <= "000000";
					when "01011101011101001" => rgb <= "000000";
					when "01011101011101010" => rgb <= "000000";
					when "01011101011101011" => rgb <= "000000";
					when "01011101011101100" => rgb <= "000000";
					when "01011101011101101" => rgb <= "000000";
					when "01011101011101110" => rgb <= "000000";
					when "01011101011101111" => rgb <= "000000";
					when "01011101011110000" => rgb <= "000000";
					when "01011101011110001" => rgb <= "000000";
					when "01011101011110010" => rgb <= "000000";
					when "01011101011110011" => rgb <= "000000";
					when "01011101011110100" => rgb <= "000000";
					when "01011101011110101" => rgb <= "000000";
					when "01011101011110110" => rgb <= "000000";
					when "01011101011110111" => rgb <= "000000";
					when "01011101011111000" => rgb <= "000000";
					when "01011101011111001" => rgb <= "000000";
					when "01011101011111010" => rgb <= "000000";
					when "01011101011111011" => rgb <= "000000";
					when "01011101011111100" => rgb <= "000000";
					when "01011101011111101" => rgb <= "000000";
					when "01011101011111110" => rgb <= "000000";
					when "01011101011111111" => rgb <= "000000";
					when "01011101100000000" => rgb <= "000000";
					when "01011101100000001" => rgb <= "000000";
					when "01011101100000010" => rgb <= "000000";
					when "01011101100000011" => rgb <= "000000";
					when "01011101100000100" => rgb <= "000000";
					when "01011101100000101" => rgb <= "000000";
					when "01011101100000110" => rgb <= "000000";
					when "01011101100000111" => rgb <= "000000";
					when "01011101100001000" => rgb <= "000000";
					when "01011101100001001" => rgb <= "000000";
					when "01011101100001010" => rgb <= "000000";
					when "01011101100001011" => rgb <= "000000";
					when "01011101100001100" => rgb <= "000000";
					when "01011101100001101" => rgb <= "000000";
					when "01011101100001110" => rgb <= "000000";
					when "01011101100001111" => rgb <= "000000";
					when "01011101100010000" => rgb <= "000000";
					when "01011101100010001" => rgb <= "000000";
					when "01011101100010010" => rgb <= "000000";
					when "01011101100010011" => rgb <= "000000";
					when "01011101100010100" => rgb <= "000000";
					when "01011101100010101" => rgb <= "000000";
					when "01011101100010110" => rgb <= "000000";
					when "01011101100010111" => rgb <= "000000";
					when "01011101100011000" => rgb <= "000000";
					when "01011101100011001" => rgb <= "000000";
					when "01011101100011010" => rgb <= "000000";
					when "01011101100011011" => rgb <= "000000";
					when "01011101100011100" => rgb <= "000000";
					when "01011101100011101" => rgb <= "000000";
					when "01011101100011110" => rgb <= "000000";
					when "01011101100011111" => rgb <= "000000";
					when "01011101100100000" => rgb <= "000000";
					when "01011101100100001" => rgb <= "000000";
					when "01011101100100010" => rgb <= "000000";
					when "01011101100100011" => rgb <= "000000";
					when "01011101100100100" => rgb <= "000000";
					when "01011101100100101" => rgb <= "000000";
					when "01011101100100110" => rgb <= "000000";
					when "01011101100100111" => rgb <= "000000";
					when "01011101100101000" => rgb <= "000000";
					when "01011101100101001" => rgb <= "000000";
					when "01011101100101010" => rgb <= "000000";
					when "01011101100101011" => rgb <= "000000";
					when "01011101100101100" => rgb <= "000000";
					when "01011101100101101" => rgb <= "000000";
					when "01011101100101110" => rgb <= "000000";
					when "01011101100101111" => rgb <= "000000";
					when "01011101100110000" => rgb <= "000000";
					when "01011101100110001" => rgb <= "000000";
					when "01011101100110010" => rgb <= "000000";
					when "01011101100110011" => rgb <= "000000";
					when "01011101100110100" => rgb <= "000000";
					when "01011101100110101" => rgb <= "000000";
					when "01011101100110110" => rgb <= "000000";
					when "01011101100110111" => rgb <= "000000";
					when "01011101100111000" => rgb <= "000000";
					when "01011101100111001" => rgb <= "000000";
					when "01011101100111010" => rgb <= "000000";
					when "01011101100111011" => rgb <= "000000";
					when "01011101100111100" => rgb <= "000000";
					when "01011101100111101" => rgb <= "000000";
					when "01011101100111110" => rgb <= "000000";
					when "01011101100111111" => rgb <= "000000";
					when "01011110000000000" => rgb <= "000000";
					when "01011110000000001" => rgb <= "000000";
					when "01011110000000010" => rgb <= "000000";
					when "01011110000000011" => rgb <= "000000";
					when "01011110000000100" => rgb <= "000000";
					when "01011110000000101" => rgb <= "000000";
					when "01011110000000110" => rgb <= "000000";
					when "01011110000000111" => rgb <= "000000";
					when "01011110000001000" => rgb <= "000000";
					when "01011110000001001" => rgb <= "000000";
					when "01011110000001010" => rgb <= "000000";
					when "01011110000001011" => rgb <= "000000";
					when "01011110000001100" => rgb <= "000000";
					when "01011110000001101" => rgb <= "000000";
					when "01011110000001110" => rgb <= "000000";
					when "01011110000001111" => rgb <= "000000";
					when "01011110000010000" => rgb <= "000000";
					when "01011110000010001" => rgb <= "000000";
					when "01011110000010010" => rgb <= "000000";
					when "01011110000010011" => rgb <= "000000";
					when "01011110000010100" => rgb <= "000000";
					when "01011110000010101" => rgb <= "000000";
					when "01011110000010110" => rgb <= "000000";
					when "01011110000010111" => rgb <= "000000";
					when "01011110000011000" => rgb <= "000000";
					when "01011110000011001" => rgb <= "000000";
					when "01011110000011010" => rgb <= "000000";
					when "01011110000011011" => rgb <= "000000";
					when "01011110000011100" => rgb <= "000000";
					when "01011110000011101" => rgb <= "000000";
					when "01011110000011110" => rgb <= "000000";
					when "01011110000011111" => rgb <= "000000";
					when "01011110000100000" => rgb <= "000000";
					when "01011110000100001" => rgb <= "000000";
					when "01011110000100010" => rgb <= "000000";
					when "01011110000100011" => rgb <= "000000";
					when "01011110000100100" => rgb <= "000000";
					when "01011110000100101" => rgb <= "000000";
					when "01011110000100110" => rgb <= "000000";
					when "01011110000100111" => rgb <= "000000";
					when "01011110000101000" => rgb <= "000000";
					when "01011110000101001" => rgb <= "000000";
					when "01011110000101010" => rgb <= "000000";
					when "01011110000101011" => rgb <= "000000";
					when "01011110000101100" => rgb <= "000000";
					when "01011110000101101" => rgb <= "000000";
					when "01011110000101110" => rgb <= "000000";
					when "01011110000101111" => rgb <= "000000";
					when "01011110000110000" => rgb <= "000000";
					when "01011110000110001" => rgb <= "000000";
					when "01011110000110010" => rgb <= "000000";
					when "01011110000110011" => rgb <= "000000";
					when "01011110000110100" => rgb <= "000000";
					when "01011110000110101" => rgb <= "000000";
					when "01011110000110110" => rgb <= "000000";
					when "01011110000110111" => rgb <= "000000";
					when "01011110000111000" => rgb <= "000000";
					when "01011110000111001" => rgb <= "000000";
					when "01011110000111010" => rgb <= "000000";
					when "01011110000111011" => rgb <= "000000";
					when "01011110000111100" => rgb <= "000000";
					when "01011110000111101" => rgb <= "000000";
					when "01011110000111110" => rgb <= "000000";
					when "01011110000111111" => rgb <= "000000";
					when "01011110001000000" => rgb <= "000000";
					when "01011110001000001" => rgb <= "000000";
					when "01011110001000010" => rgb <= "000000";
					when "01011110001000011" => rgb <= "000000";
					when "01011110001000100" => rgb <= "000000";
					when "01011110001000101" => rgb <= "000000";
					when "01011110001000110" => rgb <= "000000";
					when "01011110001000111" => rgb <= "000000";
					when "01011110001001000" => rgb <= "000000";
					when "01011110001001001" => rgb <= "000000";
					when "01011110001001010" => rgb <= "000000";
					when "01011110001001011" => rgb <= "000000";
					when "01011110001001100" => rgb <= "000000";
					when "01011110001001101" => rgb <= "000000";
					when "01011110001001110" => rgb <= "000000";
					when "01011110001001111" => rgb <= "000000";
					when "01011110001010000" => rgb <= "000000";
					when "01011110001010001" => rgb <= "000000";
					when "01011110001010010" => rgb <= "000000";
					when "01011110001010011" => rgb <= "000000";
					when "01011110001010100" => rgb <= "000000";
					when "01011110001010101" => rgb <= "000000";
					when "01011110001010110" => rgb <= "000000";
					when "01011110001010111" => rgb <= "000000";
					when "01011110001011000" => rgb <= "000000";
					when "01011110001011001" => rgb <= "000000";
					when "01011110001011010" => rgb <= "000000";
					when "01011110001011011" => rgb <= "000000";
					when "01011110001011100" => rgb <= "000000";
					when "01011110001011101" => rgb <= "000000";
					when "01011110001011110" => rgb <= "000000";
					when "01011110001011111" => rgb <= "000000";
					when "01011110001100000" => rgb <= "000000";
					when "01011110001100001" => rgb <= "000000";
					when "01011110001100010" => rgb <= "000000";
					when "01011110001100011" => rgb <= "000000";
					when "01011110001100100" => rgb <= "000000";
					when "01011110001100101" => rgb <= "000000";
					when "01011110001100110" => rgb <= "000000";
					when "01011110001100111" => rgb <= "000000";
					when "01011110001101000" => rgb <= "000000";
					when "01011110001101001" => rgb <= "000000";
					when "01011110001101010" => rgb <= "000000";
					when "01011110001101011" => rgb <= "000000";
					when "01011110001101100" => rgb <= "000000";
					when "01011110001101101" => rgb <= "000000";
					when "01011110001101110" => rgb <= "000000";
					when "01011110001101111" => rgb <= "000000";
					when "01011110001110000" => rgb <= "000000";
					when "01011110001110001" => rgb <= "000000";
					when "01011110001110010" => rgb <= "000000";
					when "01011110001110011" => rgb <= "000000";
					when "01011110001110100" => rgb <= "000000";
					when "01011110001110101" => rgb <= "000000";
					when "01011110001110110" => rgb <= "000000";
					when "01011110001110111" => rgb <= "000000";
					when "01011110001111000" => rgb <= "000000";
					when "01011110001111001" => rgb <= "000000";
					when "01011110001111010" => rgb <= "000000";
					when "01011110001111011" => rgb <= "000000";
					when "01011110001111100" => rgb <= "000000";
					when "01011110001111101" => rgb <= "000000";
					when "01011110001111110" => rgb <= "000000";
					when "01011110001111111" => rgb <= "000000";
					when "01011110010000000" => rgb <= "000000";
					when "01011110010000001" => rgb <= "000000";
					when "01011110010000010" => rgb <= "000000";
					when "01011110010000011" => rgb <= "000000";
					when "01011110010000100" => rgb <= "000000";
					when "01011110010000101" => rgb <= "000000";
					when "01011110010000110" => rgb <= "000000";
					when "01011110010000111" => rgb <= "000000";
					when "01011110010001000" => rgb <= "000000";
					when "01011110010001001" => rgb <= "000000";
					when "01011110010001010" => rgb <= "000000";
					when "01011110010001011" => rgb <= "000000";
					when "01011110010001100" => rgb <= "000000";
					when "01011110010001101" => rgb <= "000000";
					when "01011110010001110" => rgb <= "000000";
					when "01011110010001111" => rgb <= "000000";
					when "01011110010010000" => rgb <= "000000";
					when "01011110010010001" => rgb <= "000000";
					when "01011110010010010" => rgb <= "000000";
					when "01011110010010011" => rgb <= "010100";
					when "01011110010010100" => rgb <= "111000";
					when "01011110010010101" => rgb <= "101000";
					when "01011110010010110" => rgb <= "101000";
					when "01011110010010111" => rgb <= "101000";
					when "01011110010011000" => rgb <= "101000";
					when "01011110010011001" => rgb <= "101000";
					when "01011110010011010" => rgb <= "101000";
					when "01011110010011011" => rgb <= "101000";
					when "01011110010011100" => rgb <= "101000";
					when "01011110010011101" => rgb <= "101000";
					when "01011110010011110" => rgb <= "101000";
					when "01011110010011111" => rgb <= "101000";
					when "01011110010100000" => rgb <= "101000";
					when "01011110010100001" => rgb <= "101000";
					when "01011110010100010" => rgb <= "101000";
					when "01011110010100011" => rgb <= "101000";
					when "01011110010100100" => rgb <= "101000";
					when "01011110010100101" => rgb <= "101000";
					when "01011110010100110" => rgb <= "101000";
					when "01011110010100111" => rgb <= "101000";
					when "01011110010101000" => rgb <= "101000";
					when "01011110010101001" => rgb <= "101000";
					when "01011110010101010" => rgb <= "010000";
					when "01011110010101011" => rgb <= "000000";
					when "01011110010101100" => rgb <= "000000";
					when "01011110010101101" => rgb <= "000000";
					when "01011110010101110" => rgb <= "000000";
					when "01011110010101111" => rgb <= "000000";
					when "01011110010110000" => rgb <= "000000";
					when "01011110010110001" => rgb <= "000000";
					when "01011110010110010" => rgb <= "000000";
					when "01011110010110011" => rgb <= "000000";
					when "01011110010110100" => rgb <= "000000";
					when "01011110010110101" => rgb <= "000000";
					when "01011110010110110" => rgb <= "000000";
					when "01011110010110111" => rgb <= "000000";
					when "01011110010111000" => rgb <= "000000";
					when "01011110010111001" => rgb <= "000000";
					when "01011110010111010" => rgb <= "000000";
					when "01011110010111011" => rgb <= "000000";
					when "01011110010111100" => rgb <= "000000";
					when "01011110010111101" => rgb <= "000000";
					when "01011110010111110" => rgb <= "000000";
					when "01011110010111111" => rgb <= "000000";
					when "01011110011000000" => rgb <= "000000";
					when "01011110011000001" => rgb <= "000000";
					when "01011110011000010" => rgb <= "000000";
					when "01011110011000011" => rgb <= "000000";
					when "01011110011000100" => rgb <= "000000";
					when "01011110011000101" => rgb <= "000000";
					when "01011110011000110" => rgb <= "000000";
					when "01011110011000111" => rgb <= "000000";
					when "01011110011001000" => rgb <= "000000";
					when "01011110011001001" => rgb <= "000000";
					when "01011110011001010" => rgb <= "000000";
					when "01011110011001011" => rgb <= "000000";
					when "01011110011001100" => rgb <= "000000";
					when "01011110011001101" => rgb <= "000000";
					when "01011110011001110" => rgb <= "000000";
					when "01011110011001111" => rgb <= "000000";
					when "01011110011010000" => rgb <= "000000";
					when "01011110011010001" => rgb <= "000000";
					when "01011110011010010" => rgb <= "000000";
					when "01011110011010011" => rgb <= "000000";
					when "01011110011010100" => rgb <= "000000";
					when "01011110011010101" => rgb <= "000000";
					when "01011110011010110" => rgb <= "000000";
					when "01011110011010111" => rgb <= "000000";
					when "01011110011011000" => rgb <= "000000";
					when "01011110011011001" => rgb <= "000000";
					when "01011110011011010" => rgb <= "000000";
					when "01011110011011011" => rgb <= "000000";
					when "01011110011011100" => rgb <= "000000";
					when "01011110011011101" => rgb <= "000000";
					when "01011110011011110" => rgb <= "000000";
					when "01011110011011111" => rgb <= "000000";
					when "01011110011100000" => rgb <= "000000";
					when "01011110011100001" => rgb <= "000000";
					when "01011110011100010" => rgb <= "000000";
					when "01011110011100011" => rgb <= "000000";
					when "01011110011100100" => rgb <= "000000";
					when "01011110011100101" => rgb <= "000000";
					when "01011110011100110" => rgb <= "000000";
					when "01011110011100111" => rgb <= "000000";
					when "01011110011101000" => rgb <= "000000";
					when "01011110011101001" => rgb <= "000000";
					when "01011110011101010" => rgb <= "000000";
					when "01011110011101011" => rgb <= "000000";
					when "01011110011101100" => rgb <= "000000";
					when "01011110011101101" => rgb <= "000000";
					when "01011110011101110" => rgb <= "000000";
					when "01011110011101111" => rgb <= "000000";
					when "01011110011110000" => rgb <= "000000";
					when "01011110011110001" => rgb <= "000000";
					when "01011110011110010" => rgb <= "000000";
					when "01011110011110011" => rgb <= "000000";
					when "01011110011110100" => rgb <= "000000";
					when "01011110011110101" => rgb <= "000000";
					when "01011110011110110" => rgb <= "000000";
					when "01011110011110111" => rgb <= "000000";
					when "01011110011111000" => rgb <= "000000";
					when "01011110011111001" => rgb <= "000000";
					when "01011110011111010" => rgb <= "000000";
					when "01011110011111011" => rgb <= "000000";
					when "01011110011111100" => rgb <= "000000";
					when "01011110011111101" => rgb <= "000000";
					when "01011110011111110" => rgb <= "000000";
					when "01011110011111111" => rgb <= "000000";
					when "01011110100000000" => rgb <= "000000";
					when "01011110100000001" => rgb <= "000000";
					when "01011110100000010" => rgb <= "000000";
					when "01011110100000011" => rgb <= "000000";
					when "01011110100000100" => rgb <= "000000";
					when "01011110100000101" => rgb <= "000000";
					when "01011110100000110" => rgb <= "000000";
					when "01011110100000111" => rgb <= "000000";
					when "01011110100001000" => rgb <= "000000";
					when "01011110100001001" => rgb <= "000000";
					when "01011110100001010" => rgb <= "000000";
					when "01011110100001011" => rgb <= "000000";
					when "01011110100001100" => rgb <= "000000";
					when "01011110100001101" => rgb <= "000000";
					when "01011110100001110" => rgb <= "000000";
					when "01011110100001111" => rgb <= "000000";
					when "01011110100010000" => rgb <= "000000";
					when "01011110100010001" => rgb <= "000000";
					when "01011110100010010" => rgb <= "000000";
					when "01011110100010011" => rgb <= "000000";
					when "01011110100010100" => rgb <= "000000";
					when "01011110100010101" => rgb <= "000000";
					when "01011110100010110" => rgb <= "000000";
					when "01011110100010111" => rgb <= "000000";
					when "01011110100011000" => rgb <= "000000";
					when "01011110100011001" => rgb <= "000000";
					when "01011110100011010" => rgb <= "000000";
					when "01011110100011011" => rgb <= "000000";
					when "01011110100011100" => rgb <= "000000";
					when "01011110100011101" => rgb <= "000000";
					when "01011110100011110" => rgb <= "000000";
					when "01011110100011111" => rgb <= "000000";
					when "01011110100100000" => rgb <= "000000";
					when "01011110100100001" => rgb <= "000000";
					when "01011110100100010" => rgb <= "000000";
					when "01011110100100011" => rgb <= "000000";
					when "01011110100100100" => rgb <= "000000";
					when "01011110100100101" => rgb <= "000000";
					when "01011110100100110" => rgb <= "000000";
					when "01011110100100111" => rgb <= "000000";
					when "01011110100101000" => rgb <= "000000";
					when "01011110100101001" => rgb <= "000000";
					when "01011110100101010" => rgb <= "000000";
					when "01011110100101011" => rgb <= "000000";
					when "01011110100101100" => rgb <= "000000";
					when "01011110100101101" => rgb <= "000000";
					when "01011110100101110" => rgb <= "000000";
					when "01011110100101111" => rgb <= "000000";
					when "01011110100110000" => rgb <= "000000";
					when "01011110100110001" => rgb <= "000000";
					when "01011110100110010" => rgb <= "000000";
					when "01011110100110011" => rgb <= "000000";
					when "01011110100110100" => rgb <= "000000";
					when "01011110100110101" => rgb <= "000000";
					when "01011110100110110" => rgb <= "000000";
					when "01011110100110111" => rgb <= "000000";
					when "01011110100111000" => rgb <= "000000";
					when "01011110100111001" => rgb <= "000000";
					when "01011110100111010" => rgb <= "000000";
					when "01011110100111011" => rgb <= "000000";
					when "01011110100111100" => rgb <= "000000";
					when "01011110100111101" => rgb <= "000000";
					when "01011110100111110" => rgb <= "000000";
					when "01011110100111111" => rgb <= "000000";
					when "01011111000000000" => rgb <= "000000";
					when "01011111000000001" => rgb <= "000000";
					when "01011111000000010" => rgb <= "000000";
					when "01011111000000011" => rgb <= "000000";
					when "01011111000000100" => rgb <= "000000";
					when "01011111000000101" => rgb <= "000000";
					when "01011111000000110" => rgb <= "000000";
					when "01011111000000111" => rgb <= "000000";
					when "01011111000001000" => rgb <= "000000";
					when "01011111000001001" => rgb <= "000000";
					when "01011111000001010" => rgb <= "000000";
					when "01011111000001011" => rgb <= "000000";
					when "01011111000001100" => rgb <= "000000";
					when "01011111000001101" => rgb <= "000000";
					when "01011111000001110" => rgb <= "000000";
					when "01011111000001111" => rgb <= "000000";
					when "01011111000010000" => rgb <= "000000";
					when "01011111000010001" => rgb <= "000000";
					when "01011111000010010" => rgb <= "000000";
					when "01011111000010011" => rgb <= "000000";
					when "01011111000010100" => rgb <= "000000";
					when "01011111000010101" => rgb <= "000000";
					when "01011111000010110" => rgb <= "000000";
					when "01011111000010111" => rgb <= "000000";
					when "01011111000011000" => rgb <= "000000";
					when "01011111000011001" => rgb <= "000000";
					when "01011111000011010" => rgb <= "000000";
					when "01011111000011011" => rgb <= "000000";
					when "01011111000011100" => rgb <= "000000";
					when "01011111000011101" => rgb <= "000000";
					when "01011111000011110" => rgb <= "000000";
					when "01011111000011111" => rgb <= "000000";
					when "01011111000100000" => rgb <= "000000";
					when "01011111000100001" => rgb <= "000000";
					when "01011111000100010" => rgb <= "000000";
					when "01011111000100011" => rgb <= "000000";
					when "01011111000100100" => rgb <= "000000";
					when "01011111000100101" => rgb <= "000000";
					when "01011111000100110" => rgb <= "000000";
					when "01011111000100111" => rgb <= "000000";
					when "01011111000101000" => rgb <= "000000";
					when "01011111000101001" => rgb <= "000000";
					when "01011111000101010" => rgb <= "000000";
					when "01011111000101011" => rgb <= "000000";
					when "01011111000101100" => rgb <= "000000";
					when "01011111000101101" => rgb <= "000000";
					when "01011111000101110" => rgb <= "000000";
					when "01011111000101111" => rgb <= "000000";
					when "01011111000110000" => rgb <= "000000";
					when "01011111000110001" => rgb <= "000000";
					when "01011111000110010" => rgb <= "000000";
					when "01011111000110011" => rgb <= "000000";
					when "01011111000110100" => rgb <= "000000";
					when "01011111000110101" => rgb <= "000000";
					when "01011111000110110" => rgb <= "000000";
					when "01011111000110111" => rgb <= "000000";
					when "01011111000111000" => rgb <= "000000";
					when "01011111000111001" => rgb <= "000000";
					when "01011111000111010" => rgb <= "000000";
					when "01011111000111011" => rgb <= "000000";
					when "01011111000111100" => rgb <= "000000";
					when "01011111000111101" => rgb <= "000000";
					when "01011111000111110" => rgb <= "000000";
					when "01011111000111111" => rgb <= "000000";
					when "01011111001000000" => rgb <= "000000";
					when "01011111001000001" => rgb <= "000000";
					when "01011111001000010" => rgb <= "000000";
					when "01011111001000011" => rgb <= "000000";
					when "01011111001000100" => rgb <= "000000";
					when "01011111001000101" => rgb <= "000000";
					when "01011111001000110" => rgb <= "000000";
					when "01011111001000111" => rgb <= "000000";
					when "01011111001001000" => rgb <= "000000";
					when "01011111001001001" => rgb <= "000000";
					when "01011111001001010" => rgb <= "000000";
					when "01011111001001011" => rgb <= "000000";
					when "01011111001001100" => rgb <= "000000";
					when "01011111001001101" => rgb <= "000000";
					when "01011111001001110" => rgb <= "000000";
					when "01011111001001111" => rgb <= "000000";
					when "01011111001010000" => rgb <= "000000";
					when "01011111001010001" => rgb <= "000000";
					when "01011111001010010" => rgb <= "000000";
					when "01011111001010011" => rgb <= "000000";
					when "01011111001010100" => rgb <= "000000";
					when "01011111001010101" => rgb <= "000000";
					when "01011111001010110" => rgb <= "000000";
					when "01011111001010111" => rgb <= "000000";
					when "01011111001011000" => rgb <= "000000";
					when "01011111001011001" => rgb <= "000000";
					when "01011111001011010" => rgb <= "000000";
					when "01011111001011011" => rgb <= "000000";
					when "01011111001011100" => rgb <= "000000";
					when "01011111001011101" => rgb <= "000000";
					when "01011111001011110" => rgb <= "000000";
					when "01011111001011111" => rgb <= "000000";
					when "01011111001100000" => rgb <= "000000";
					when "01011111001100001" => rgb <= "000000";
					when "01011111001100010" => rgb <= "000000";
					when "01011111001100011" => rgb <= "000000";
					when "01011111001100100" => rgb <= "000000";
					when "01011111001100101" => rgb <= "000000";
					when "01011111001100110" => rgb <= "000000";
					when "01011111001100111" => rgb <= "000000";
					when "01011111001101000" => rgb <= "000000";
					when "01011111001101001" => rgb <= "000000";
					when "01011111001101010" => rgb <= "000000";
					when "01011111001101011" => rgb <= "000000";
					when "01011111001101100" => rgb <= "000000";
					when "01011111001101101" => rgb <= "000000";
					when "01011111001101110" => rgb <= "000000";
					when "01011111001101111" => rgb <= "000000";
					when "01011111001110000" => rgb <= "000000";
					when "01011111001110001" => rgb <= "000000";
					when "01011111001110010" => rgb <= "000000";
					when "01011111001110011" => rgb <= "000000";
					when "01011111001110100" => rgb <= "000000";
					when "01011111001110101" => rgb <= "000000";
					when "01011111001110110" => rgb <= "000000";
					when "01011111001110111" => rgb <= "000000";
					when "01011111001111000" => rgb <= "000000";
					when "01011111001111001" => rgb <= "000000";
					when "01011111001111010" => rgb <= "000000";
					when "01011111001111011" => rgb <= "000000";
					when "01011111001111100" => rgb <= "000000";
					when "01011111001111101" => rgb <= "000000";
					when "01011111001111110" => rgb <= "000000";
					when "01011111001111111" => rgb <= "000000";
					when "01011111010000000" => rgb <= "000000";
					when "01011111010000001" => rgb <= "000000";
					when "01011111010000010" => rgb <= "000000";
					when "01011111010000011" => rgb <= "000000";
					when "01011111010000100" => rgb <= "000000";
					when "01011111010000101" => rgb <= "000000";
					when "01011111010000110" => rgb <= "000000";
					when "01011111010000111" => rgb <= "000000";
					when "01011111010001000" => rgb <= "000000";
					when "01011111010001001" => rgb <= "000000";
					when "01011111010001010" => rgb <= "000000";
					when "01011111010001011" => rgb <= "000000";
					when "01011111010001100" => rgb <= "000000";
					when "01011111010001101" => rgb <= "000000";
					when "01011111010001110" => rgb <= "000000";
					when "01011111010001111" => rgb <= "000000";
					when "01011111010010000" => rgb <= "000000";
					when "01011111010010001" => rgb <= "000000";
					when "01011111010010010" => rgb <= "000000";
					when "01011111010010011" => rgb <= "010100";
					when "01011111010010100" => rgb <= "111000";
					when "01011111010010101" => rgb <= "101000";
					when "01011111010010110" => rgb <= "101000";
					when "01011111010010111" => rgb <= "101000";
					when "01011111010011000" => rgb <= "101000";
					when "01011111010011001" => rgb <= "101000";
					when "01011111010011010" => rgb <= "101000";
					when "01011111010011011" => rgb <= "101000";
					when "01011111010011100" => rgb <= "101000";
					when "01011111010011101" => rgb <= "101000";
					when "01011111010011110" => rgb <= "101000";
					when "01011111010011111" => rgb <= "101000";
					when "01011111010100000" => rgb <= "101000";
					when "01011111010100001" => rgb <= "101000";
					when "01011111010100010" => rgb <= "101000";
					when "01011111010100011" => rgb <= "101000";
					when "01011111010100100" => rgb <= "101000";
					when "01011111010100101" => rgb <= "101000";
					when "01011111010100110" => rgb <= "101000";
					when "01011111010100111" => rgb <= "101000";
					when "01011111010101000" => rgb <= "101000";
					when "01011111010101001" => rgb <= "101000";
					when "01011111010101010" => rgb <= "010000";
					when "01011111010101011" => rgb <= "000000";
					when "01011111010101100" => rgb <= "000000";
					when "01011111010101101" => rgb <= "000000";
					when "01011111010101110" => rgb <= "000000";
					when "01011111010101111" => rgb <= "000000";
					when "01011111010110000" => rgb <= "000000";
					when "01011111010110001" => rgb <= "000000";
					when "01011111010110010" => rgb <= "000000";
					when "01011111010110011" => rgb <= "000000";
					when "01011111010110100" => rgb <= "000000";
					when "01011111010110101" => rgb <= "000000";
					when "01011111010110110" => rgb <= "000000";
					when "01011111010110111" => rgb <= "000000";
					when "01011111010111000" => rgb <= "000000";
					when "01011111010111001" => rgb <= "000000";
					when "01011111010111010" => rgb <= "000000";
					when "01011111010111011" => rgb <= "000000";
					when "01011111010111100" => rgb <= "000000";
					when "01011111010111101" => rgb <= "000000";
					when "01011111010111110" => rgb <= "000000";
					when "01011111010111111" => rgb <= "000000";
					when "01011111011000000" => rgb <= "000000";
					when "01011111011000001" => rgb <= "000000";
					when "01011111011000010" => rgb <= "000000";
					when "01011111011000011" => rgb <= "000000";
					when "01011111011000100" => rgb <= "000000";
					when "01011111011000101" => rgb <= "000000";
					when "01011111011000110" => rgb <= "000000";
					when "01011111011000111" => rgb <= "000000";
					when "01011111011001000" => rgb <= "000000";
					when "01011111011001001" => rgb <= "000000";
					when "01011111011001010" => rgb <= "000000";
					when "01011111011001011" => rgb <= "000000";
					when "01011111011001100" => rgb <= "000000";
					when "01011111011001101" => rgb <= "000000";
					when "01011111011001110" => rgb <= "000000";
					when "01011111011001111" => rgb <= "000000";
					when "01011111011010000" => rgb <= "000000";
					when "01011111011010001" => rgb <= "000000";
					when "01011111011010010" => rgb <= "000000";
					when "01011111011010011" => rgb <= "000000";
					when "01011111011010100" => rgb <= "000000";
					when "01011111011010101" => rgb <= "000000";
					when "01011111011010110" => rgb <= "000000";
					when "01011111011010111" => rgb <= "000000";
					when "01011111011011000" => rgb <= "000000";
					when "01011111011011001" => rgb <= "000000";
					when "01011111011011010" => rgb <= "000000";
					when "01011111011011011" => rgb <= "000000";
					when "01011111011011100" => rgb <= "000000";
					when "01011111011011101" => rgb <= "000000";
					when "01011111011011110" => rgb <= "000000";
					when "01011111011011111" => rgb <= "000000";
					when "01011111011100000" => rgb <= "000000";
					when "01011111011100001" => rgb <= "000000";
					when "01011111011100010" => rgb <= "000000";
					when "01011111011100011" => rgb <= "000000";
					when "01011111011100100" => rgb <= "000000";
					when "01011111011100101" => rgb <= "000000";
					when "01011111011100110" => rgb <= "000000";
					when "01011111011100111" => rgb <= "000000";
					when "01011111011101000" => rgb <= "000000";
					when "01011111011101001" => rgb <= "000000";
					when "01011111011101010" => rgb <= "000000";
					when "01011111011101011" => rgb <= "000000";
					when "01011111011101100" => rgb <= "000000";
					when "01011111011101101" => rgb <= "000000";
					when "01011111011101110" => rgb <= "000000";
					when "01011111011101111" => rgb <= "000000";
					when "01011111011110000" => rgb <= "000000";
					when "01011111011110001" => rgb <= "000000";
					when "01011111011110010" => rgb <= "000000";
					when "01011111011110011" => rgb <= "000000";
					when "01011111011110100" => rgb <= "000000";
					when "01011111011110101" => rgb <= "000000";
					when "01011111011110110" => rgb <= "000000";
					when "01011111011110111" => rgb <= "000000";
					when "01011111011111000" => rgb <= "000000";
					when "01011111011111001" => rgb <= "000000";
					when "01011111011111010" => rgb <= "000000";
					when "01011111011111011" => rgb <= "000000";
					when "01011111011111100" => rgb <= "000000";
					when "01011111011111101" => rgb <= "000000";
					when "01011111011111110" => rgb <= "000000";
					when "01011111011111111" => rgb <= "000000";
					when "01011111100000000" => rgb <= "000000";
					when "01011111100000001" => rgb <= "000000";
					when "01011111100000010" => rgb <= "000000";
					when "01011111100000011" => rgb <= "000000";
					when "01011111100000100" => rgb <= "000000";
					when "01011111100000101" => rgb <= "000000";
					when "01011111100000110" => rgb <= "000000";
					when "01011111100000111" => rgb <= "000000";
					when "01011111100001000" => rgb <= "000000";
					when "01011111100001001" => rgb <= "000000";
					when "01011111100001010" => rgb <= "000000";
					when "01011111100001011" => rgb <= "000000";
					when "01011111100001100" => rgb <= "000000";
					when "01011111100001101" => rgb <= "000000";
					when "01011111100001110" => rgb <= "000000";
					when "01011111100001111" => rgb <= "000000";
					when "01011111100010000" => rgb <= "000000";
					when "01011111100010001" => rgb <= "000000";
					when "01011111100010010" => rgb <= "000000";
					when "01011111100010011" => rgb <= "000000";
					when "01011111100010100" => rgb <= "000000";
					when "01011111100010101" => rgb <= "000000";
					when "01011111100010110" => rgb <= "000000";
					when "01011111100010111" => rgb <= "000000";
					when "01011111100011000" => rgb <= "000000";
					when "01011111100011001" => rgb <= "000000";
					when "01011111100011010" => rgb <= "000000";
					when "01011111100011011" => rgb <= "000000";
					when "01011111100011100" => rgb <= "000000";
					when "01011111100011101" => rgb <= "000000";
					when "01011111100011110" => rgb <= "000000";
					when "01011111100011111" => rgb <= "000000";
					when "01011111100100000" => rgb <= "000000";
					when "01011111100100001" => rgb <= "000000";
					when "01011111100100010" => rgb <= "000000";
					when "01011111100100011" => rgb <= "000000";
					when "01011111100100100" => rgb <= "000000";
					when "01011111100100101" => rgb <= "000000";
					when "01011111100100110" => rgb <= "000000";
					when "01011111100100111" => rgb <= "000000";
					when "01011111100101000" => rgb <= "000000";
					when "01011111100101001" => rgb <= "000000";
					when "01011111100101010" => rgb <= "000000";
					when "01011111100101011" => rgb <= "000000";
					when "01011111100101100" => rgb <= "000000";
					when "01011111100101101" => rgb <= "000000";
					when "01011111100101110" => rgb <= "000000";
					when "01011111100101111" => rgb <= "000000";
					when "01011111100110000" => rgb <= "000000";
					when "01011111100110001" => rgb <= "000000";
					when "01011111100110010" => rgb <= "000000";
					when "01011111100110011" => rgb <= "000000";
					when "01011111100110100" => rgb <= "000000";
					when "01011111100110101" => rgb <= "000000";
					when "01011111100110110" => rgb <= "000000";
					when "01011111100110111" => rgb <= "000000";
					when "01011111100111000" => rgb <= "000000";
					when "01011111100111001" => rgb <= "000000";
					when "01011111100111010" => rgb <= "000000";
					when "01011111100111011" => rgb <= "000000";
					when "01011111100111100" => rgb <= "000000";
					when "01011111100111101" => rgb <= "000000";
					when "01011111100111110" => rgb <= "000000";
					when "01011111100111111" => rgb <= "000000";
					when "01100000000000000" => rgb <= "000000";
					when "01100000000000001" => rgb <= "000000";
					when "01100000000000010" => rgb <= "000000";
					when "01100000000000011" => rgb <= "000000";
					when "01100000000000100" => rgb <= "000000";
					when "01100000000000101" => rgb <= "000000";
					when "01100000000000110" => rgb <= "000000";
					when "01100000000000111" => rgb <= "000000";
					when "01100000000001000" => rgb <= "000000";
					when "01100000000001001" => rgb <= "000000";
					when "01100000000001010" => rgb <= "000000";
					when "01100000000001011" => rgb <= "000000";
					when "01100000000001100" => rgb <= "000000";
					when "01100000000001101" => rgb <= "000000";
					when "01100000000001110" => rgb <= "000000";
					when "01100000000001111" => rgb <= "000000";
					when "01100000000010000" => rgb <= "000000";
					when "01100000000010001" => rgb <= "000000";
					when "01100000000010010" => rgb <= "000000";
					when "01100000000010011" => rgb <= "000000";
					when "01100000000010100" => rgb <= "000000";
					when "01100000000010101" => rgb <= "000000";
					when "01100000000010110" => rgb <= "000000";
					when "01100000000010111" => rgb <= "000000";
					when "01100000000011000" => rgb <= "000000";
					when "01100000000011001" => rgb <= "000000";
					when "01100000000011010" => rgb <= "000000";
					when "01100000000011011" => rgb <= "000000";
					when "01100000000011100" => rgb <= "000000";
					when "01100000000011101" => rgb <= "000000";
					when "01100000000011110" => rgb <= "000000";
					when "01100000000011111" => rgb <= "000000";
					when "01100000000100000" => rgb <= "000000";
					when "01100000000100001" => rgb <= "000000";
					when "01100000000100010" => rgb <= "000000";
					when "01100000000100011" => rgb <= "000000";
					when "01100000000100100" => rgb <= "000000";
					when "01100000000100101" => rgb <= "000000";
					when "01100000000100110" => rgb <= "000000";
					when "01100000000100111" => rgb <= "000000";
					when "01100000000101000" => rgb <= "000000";
					when "01100000000101001" => rgb <= "000000";
					when "01100000000101010" => rgb <= "000000";
					when "01100000000101011" => rgb <= "000000";
					when "01100000000101100" => rgb <= "000000";
					when "01100000000101101" => rgb <= "000000";
					when "01100000000101110" => rgb <= "000000";
					when "01100000000101111" => rgb <= "000000";
					when "01100000000110000" => rgb <= "000000";
					when "01100000000110001" => rgb <= "000000";
					when "01100000000110010" => rgb <= "000000";
					when "01100000000110011" => rgb <= "000000";
					when "01100000000110100" => rgb <= "000000";
					when "01100000000110101" => rgb <= "000000";
					when "01100000000110110" => rgb <= "000000";
					when "01100000000110111" => rgb <= "000000";
					when "01100000000111000" => rgb <= "000000";
					when "01100000000111001" => rgb <= "000000";
					when "01100000000111010" => rgb <= "000000";
					when "01100000000111011" => rgb <= "000000";
					when "01100000000111100" => rgb <= "000000";
					when "01100000000111101" => rgb <= "000000";
					when "01100000000111110" => rgb <= "000000";
					when "01100000000111111" => rgb <= "000000";
					when "01100000001000000" => rgb <= "000000";
					when "01100000001000001" => rgb <= "000000";
					when "01100000001000010" => rgb <= "000000";
					when "01100000001000011" => rgb <= "000000";
					when "01100000001000100" => rgb <= "000000";
					when "01100000001000101" => rgb <= "000000";
					when "01100000001000110" => rgb <= "000000";
					when "01100000001000111" => rgb <= "000000";
					when "01100000001001000" => rgb <= "000000";
					when "01100000001001001" => rgb <= "000000";
					when "01100000001001010" => rgb <= "000000";
					when "01100000001001011" => rgb <= "000000";
					when "01100000001001100" => rgb <= "000000";
					when "01100000001001101" => rgb <= "000000";
					when "01100000001001110" => rgb <= "000000";
					when "01100000001001111" => rgb <= "000000";
					when "01100000001010000" => rgb <= "000000";
					when "01100000001010001" => rgb <= "000000";
					when "01100000001010010" => rgb <= "000000";
					when "01100000001010011" => rgb <= "000000";
					when "01100000001010100" => rgb <= "000000";
					when "01100000001010101" => rgb <= "000000";
					when "01100000001010110" => rgb <= "000000";
					when "01100000001010111" => rgb <= "000000";
					when "01100000001011000" => rgb <= "000000";
					when "01100000001011001" => rgb <= "000000";
					when "01100000001011010" => rgb <= "000000";
					when "01100000001011011" => rgb <= "000000";
					when "01100000001011100" => rgb <= "000000";
					when "01100000001011101" => rgb <= "000000";
					when "01100000001011110" => rgb <= "000000";
					when "01100000001011111" => rgb <= "000000";
					when "01100000001100000" => rgb <= "000000";
					when "01100000001100001" => rgb <= "000000";
					when "01100000001100010" => rgb <= "000000";
					when "01100000001100011" => rgb <= "000000";
					when "01100000001100100" => rgb <= "000000";
					when "01100000001100101" => rgb <= "000000";
					when "01100000001100110" => rgb <= "000000";
					when "01100000001100111" => rgb <= "000000";
					when "01100000001101000" => rgb <= "000000";
					when "01100000001101001" => rgb <= "000000";
					when "01100000001101010" => rgb <= "000000";
					when "01100000001101011" => rgb <= "000000";
					when "01100000001101100" => rgb <= "000000";
					when "01100000001101101" => rgb <= "000000";
					when "01100000001101110" => rgb <= "000000";
					when "01100000001101111" => rgb <= "000000";
					when "01100000001110000" => rgb <= "000000";
					when "01100000001110001" => rgb <= "000000";
					when "01100000001110010" => rgb <= "000000";
					when "01100000001110011" => rgb <= "000000";
					when "01100000001110100" => rgb <= "000000";
					when "01100000001110101" => rgb <= "000000";
					when "01100000001110110" => rgb <= "000000";
					when "01100000001110111" => rgb <= "000000";
					when "01100000001111000" => rgb <= "000000";
					when "01100000001111001" => rgb <= "000000";
					when "01100000001111010" => rgb <= "000000";
					when "01100000001111011" => rgb <= "000000";
					when "01100000001111100" => rgb <= "000000";
					when "01100000001111101" => rgb <= "000000";
					when "01100000001111110" => rgb <= "000000";
					when "01100000001111111" => rgb <= "000000";
					when "01100000010000000" => rgb <= "000000";
					when "01100000010000001" => rgb <= "000000";
					when "01100000010000010" => rgb <= "000000";
					when "01100000010000011" => rgb <= "000000";
					when "01100000010000100" => rgb <= "000000";
					when "01100000010000101" => rgb <= "000000";
					when "01100000010000110" => rgb <= "000000";
					when "01100000010000111" => rgb <= "000000";
					when "01100000010001000" => rgb <= "000000";
					when "01100000010001001" => rgb <= "000000";
					when "01100000010001010" => rgb <= "000000";
					when "01100000010001011" => rgb <= "000000";
					when "01100000010001100" => rgb <= "000000";
					when "01100000010001101" => rgb <= "000000";
					when "01100000010001110" => rgb <= "000000";
					when "01100000010001111" => rgb <= "000000";
					when "01100000010010000" => rgb <= "000000";
					when "01100000010010001" => rgb <= "000000";
					when "01100000010010010" => rgb <= "000000";
					when "01100000010010011" => rgb <= "010000";
					when "01100000010010100" => rgb <= "101000";
					when "01100000010010101" => rgb <= "101000";
					when "01100000010010110" => rgb <= "101000";
					when "01100000010010111" => rgb <= "101000";
					when "01100000010011000" => rgb <= "101000";
					when "01100000010011001" => rgb <= "101000";
					when "01100000010011010" => rgb <= "101000";
					when "01100000010011011" => rgb <= "101000";
					when "01100000010011100" => rgb <= "101000";
					when "01100000010011101" => rgb <= "101000";
					when "01100000010011110" => rgb <= "101000";
					when "01100000010011111" => rgb <= "101000";
					when "01100000010100000" => rgb <= "101000";
					when "01100000010100001" => rgb <= "101000";
					when "01100000010100010" => rgb <= "101000";
					when "01100000010100011" => rgb <= "101000";
					when "01100000010100100" => rgb <= "101000";
					when "01100000010100101" => rgb <= "101000";
					when "01100000010100110" => rgb <= "101000";
					when "01100000010100111" => rgb <= "101000";
					when "01100000010101000" => rgb <= "101000";
					when "01100000010101001" => rgb <= "101000";
					when "01100000010101010" => rgb <= "010000";
					when "01100000010101011" => rgb <= "000000";
					when "01100000010101100" => rgb <= "000000";
					when "01100000010101101" => rgb <= "000000";
					when "01100000010101110" => rgb <= "000000";
					when "01100000010101111" => rgb <= "000000";
					when "01100000010110000" => rgb <= "000000";
					when "01100000010110001" => rgb <= "000000";
					when "01100000010110010" => rgb <= "000000";
					when "01100000010110011" => rgb <= "000000";
					when "01100000010110100" => rgb <= "000000";
					when "01100000010110101" => rgb <= "000000";
					when "01100000010110110" => rgb <= "000000";
					when "01100000010110111" => rgb <= "000000";
					when "01100000010111000" => rgb <= "000000";
					when "01100000010111001" => rgb <= "000000";
					when "01100000010111010" => rgb <= "000000";
					when "01100000010111011" => rgb <= "000000";
					when "01100000010111100" => rgb <= "000000";
					when "01100000010111101" => rgb <= "000000";
					when "01100000010111110" => rgb <= "000000";
					when "01100000010111111" => rgb <= "000000";
					when "01100000011000000" => rgb <= "000000";
					when "01100000011000001" => rgb <= "000000";
					when "01100000011000010" => rgb <= "000000";
					when "01100000011000011" => rgb <= "000000";
					when "01100000011000100" => rgb <= "000000";
					when "01100000011000101" => rgb <= "000000";
					when "01100000011000110" => rgb <= "000000";
					when "01100000011000111" => rgb <= "000000";
					when "01100000011001000" => rgb <= "000000";
					when "01100000011001001" => rgb <= "000000";
					when "01100000011001010" => rgb <= "000000";
					when "01100000011001011" => rgb <= "000000";
					when "01100000011001100" => rgb <= "000000";
					when "01100000011001101" => rgb <= "000000";
					when "01100000011001110" => rgb <= "000000";
					when "01100000011001111" => rgb <= "000000";
					when "01100000011010000" => rgb <= "000000";
					when "01100000011010001" => rgb <= "000000";
					when "01100000011010010" => rgb <= "000000";
					when "01100000011010011" => rgb <= "000000";
					when "01100000011010100" => rgb <= "000000";
					when "01100000011010101" => rgb <= "000000";
					when "01100000011010110" => rgb <= "000000";
					when "01100000011010111" => rgb <= "000000";
					when "01100000011011000" => rgb <= "000000";
					when "01100000011011001" => rgb <= "000000";
					when "01100000011011010" => rgb <= "000000";
					when "01100000011011011" => rgb <= "000000";
					when "01100000011011100" => rgb <= "000000";
					when "01100000011011101" => rgb <= "000000";
					when "01100000011011110" => rgb <= "000000";
					when "01100000011011111" => rgb <= "000000";
					when "01100000011100000" => rgb <= "000000";
					when "01100000011100001" => rgb <= "000000";
					when "01100000011100010" => rgb <= "000000";
					when "01100000011100011" => rgb <= "000000";
					when "01100000011100100" => rgb <= "000000";
					when "01100000011100101" => rgb <= "000000";
					when "01100000011100110" => rgb <= "000000";
					when "01100000011100111" => rgb <= "000000";
					when "01100000011101000" => rgb <= "000000";
					when "01100000011101001" => rgb <= "000000";
					when "01100000011101010" => rgb <= "000000";
					when "01100000011101011" => rgb <= "000000";
					when "01100000011101100" => rgb <= "000000";
					when "01100000011101101" => rgb <= "000000";
					when "01100000011101110" => rgb <= "000000";
					when "01100000011101111" => rgb <= "000000";
					when "01100000011110000" => rgb <= "000000";
					when "01100000011110001" => rgb <= "000000";
					when "01100000011110010" => rgb <= "000000";
					when "01100000011110011" => rgb <= "000000";
					when "01100000011110100" => rgb <= "000000";
					when "01100000011110101" => rgb <= "000000";
					when "01100000011110110" => rgb <= "000000";
					when "01100000011110111" => rgb <= "000000";
					when "01100000011111000" => rgb <= "000000";
					when "01100000011111001" => rgb <= "000000";
					when "01100000011111010" => rgb <= "000000";
					when "01100000011111011" => rgb <= "000000";
					when "01100000011111100" => rgb <= "000000";
					when "01100000011111101" => rgb <= "000000";
					when "01100000011111110" => rgb <= "000000";
					when "01100000011111111" => rgb <= "000000";
					when "01100000100000000" => rgb <= "000000";
					when "01100000100000001" => rgb <= "000000";
					when "01100000100000010" => rgb <= "000000";
					when "01100000100000011" => rgb <= "000000";
					when "01100000100000100" => rgb <= "000000";
					when "01100000100000101" => rgb <= "000000";
					when "01100000100000110" => rgb <= "000000";
					when "01100000100000111" => rgb <= "000000";
					when "01100000100001000" => rgb <= "000000";
					when "01100000100001001" => rgb <= "000000";
					when "01100000100001010" => rgb <= "000000";
					when "01100000100001011" => rgb <= "000000";
					when "01100000100001100" => rgb <= "000000";
					when "01100000100001101" => rgb <= "000000";
					when "01100000100001110" => rgb <= "000000";
					when "01100000100001111" => rgb <= "000000";
					when "01100000100010000" => rgb <= "000000";
					when "01100000100010001" => rgb <= "000000";
					when "01100000100010010" => rgb <= "000000";
					when "01100000100010011" => rgb <= "000000";
					when "01100000100010100" => rgb <= "000000";
					when "01100000100010101" => rgb <= "000000";
					when "01100000100010110" => rgb <= "000000";
					when "01100000100010111" => rgb <= "000000";
					when "01100000100011000" => rgb <= "000000";
					when "01100000100011001" => rgb <= "000000";
					when "01100000100011010" => rgb <= "000000";
					when "01100000100011011" => rgb <= "000000";
					when "01100000100011100" => rgb <= "000000";
					when "01100000100011101" => rgb <= "000000";
					when "01100000100011110" => rgb <= "000000";
					when "01100000100011111" => rgb <= "000000";
					when "01100000100100000" => rgb <= "000000";
					when "01100000100100001" => rgb <= "000000";
					when "01100000100100010" => rgb <= "000000";
					when "01100000100100011" => rgb <= "000000";
					when "01100000100100100" => rgb <= "000000";
					when "01100000100100101" => rgb <= "000000";
					when "01100000100100110" => rgb <= "000000";
					when "01100000100100111" => rgb <= "000000";
					when "01100000100101000" => rgb <= "000000";
					when "01100000100101001" => rgb <= "000000";
					when "01100000100101010" => rgb <= "000000";
					when "01100000100101011" => rgb <= "000000";
					when "01100000100101100" => rgb <= "000000";
					when "01100000100101101" => rgb <= "000000";
					when "01100000100101110" => rgb <= "000000";
					when "01100000100101111" => rgb <= "000000";
					when "01100000100110000" => rgb <= "000000";
					when "01100000100110001" => rgb <= "000000";
					when "01100000100110010" => rgb <= "000000";
					when "01100000100110011" => rgb <= "000000";
					when "01100000100110100" => rgb <= "000000";
					when "01100000100110101" => rgb <= "000000";
					when "01100000100110110" => rgb <= "000000";
					when "01100000100110111" => rgb <= "000000";
					when "01100000100111000" => rgb <= "000000";
					when "01100000100111001" => rgb <= "000000";
					when "01100000100111010" => rgb <= "000000";
					when "01100000100111011" => rgb <= "000000";
					when "01100000100111100" => rgb <= "000000";
					when "01100000100111101" => rgb <= "000000";
					when "01100000100111110" => rgb <= "000000";
					when "01100000100111111" => rgb <= "000000";
					when "01100001000000000" => rgb <= "000000";
					when "01100001000000001" => rgb <= "000000";
					when "01100001000000010" => rgb <= "000000";
					when "01100001000000011" => rgb <= "000000";
					when "01100001000000100" => rgb <= "000000";
					when "01100001000000101" => rgb <= "000000";
					when "01100001000000110" => rgb <= "000000";
					when "01100001000000111" => rgb <= "000000";
					when "01100001000001000" => rgb <= "000000";
					when "01100001000001001" => rgb <= "000000";
					when "01100001000001010" => rgb <= "000000";
					when "01100001000001011" => rgb <= "000000";
					when "01100001000001100" => rgb <= "000000";
					when "01100001000001101" => rgb <= "000000";
					when "01100001000001110" => rgb <= "000000";
					when "01100001000001111" => rgb <= "000000";
					when "01100001000010000" => rgb <= "000000";
					when "01100001000010001" => rgb <= "000000";
					when "01100001000010010" => rgb <= "000000";
					when "01100001000010011" => rgb <= "000000";
					when "01100001000010100" => rgb <= "000000";
					when "01100001000010101" => rgb <= "000000";
					when "01100001000010110" => rgb <= "000000";
					when "01100001000010111" => rgb <= "000000";
					when "01100001000011000" => rgb <= "000000";
					when "01100001000011001" => rgb <= "000000";
					when "01100001000011010" => rgb <= "000000";
					when "01100001000011011" => rgb <= "000000";
					when "01100001000011100" => rgb <= "000000";
					when "01100001000011101" => rgb <= "000000";
					when "01100001000011110" => rgb <= "000000";
					when "01100001000011111" => rgb <= "000000";
					when "01100001000100000" => rgb <= "000000";
					when "01100001000100001" => rgb <= "000000";
					when "01100001000100010" => rgb <= "000000";
					when "01100001000100011" => rgb <= "000000";
					when "01100001000100100" => rgb <= "000000";
					when "01100001000100101" => rgb <= "000000";
					when "01100001000100110" => rgb <= "000000";
					when "01100001000100111" => rgb <= "000000";
					when "01100001000101000" => rgb <= "000000";
					when "01100001000101001" => rgb <= "000000";
					when "01100001000101010" => rgb <= "000000";
					when "01100001000101011" => rgb <= "000000";
					when "01100001000101100" => rgb <= "000000";
					when "01100001000101101" => rgb <= "000000";
					when "01100001000101110" => rgb <= "000000";
					when "01100001000101111" => rgb <= "000000";
					when "01100001000110000" => rgb <= "000000";
					when "01100001000110001" => rgb <= "000000";
					when "01100001000110010" => rgb <= "000000";
					when "01100001000110011" => rgb <= "000000";
					when "01100001000110100" => rgb <= "000000";
					when "01100001000110101" => rgb <= "000000";
					when "01100001000110110" => rgb <= "000000";
					when "01100001000110111" => rgb <= "000000";
					when "01100001000111000" => rgb <= "000000";
					when "01100001000111001" => rgb <= "000000";
					when "01100001000111010" => rgb <= "000000";
					when "01100001000111011" => rgb <= "000000";
					when "01100001000111100" => rgb <= "000000";
					when "01100001000111101" => rgb <= "000000";
					when "01100001000111110" => rgb <= "000000";
					when "01100001000111111" => rgb <= "000000";
					when "01100001001000000" => rgb <= "000000";
					when "01100001001000001" => rgb <= "000000";
					when "01100001001000010" => rgb <= "000000";
					when "01100001001000011" => rgb <= "000000";
					when "01100001001000100" => rgb <= "000000";
					when "01100001001000101" => rgb <= "000000";
					when "01100001001000110" => rgb <= "000000";
					when "01100001001000111" => rgb <= "000000";
					when "01100001001001000" => rgb <= "000000";
					when "01100001001001001" => rgb <= "000000";
					when "01100001001001010" => rgb <= "000000";
					when "01100001001001011" => rgb <= "000000";
					when "01100001001001100" => rgb <= "000000";
					when "01100001001001101" => rgb <= "000000";
					when "01100001001001110" => rgb <= "000000";
					when "01100001001001111" => rgb <= "000000";
					when "01100001001010000" => rgb <= "000000";
					when "01100001001010001" => rgb <= "000000";
					when "01100001001010010" => rgb <= "000000";
					when "01100001001010011" => rgb <= "000000";
					when "01100001001010100" => rgb <= "000000";
					when "01100001001010101" => rgb <= "000000";
					when "01100001001010110" => rgb <= "000000";
					when "01100001001010111" => rgb <= "000000";
					when "01100001001011000" => rgb <= "000000";
					when "01100001001011001" => rgb <= "000000";
					when "01100001001011010" => rgb <= "000000";
					when "01100001001011011" => rgb <= "000000";
					when "01100001001011100" => rgb <= "000000";
					when "01100001001011101" => rgb <= "000000";
					when "01100001001011110" => rgb <= "000000";
					when "01100001001011111" => rgb <= "000000";
					when "01100001001100000" => rgb <= "000000";
					when "01100001001100001" => rgb <= "000000";
					when "01100001001100010" => rgb <= "000000";
					when "01100001001100011" => rgb <= "000000";
					when "01100001001100100" => rgb <= "000000";
					when "01100001001100101" => rgb <= "000000";
					when "01100001001100110" => rgb <= "000000";
					when "01100001001100111" => rgb <= "000000";
					when "01100001001101000" => rgb <= "000000";
					when "01100001001101001" => rgb <= "000000";
					when "01100001001101010" => rgb <= "000000";
					when "01100001001101011" => rgb <= "000000";
					when "01100001001101100" => rgb <= "000000";
					when "01100001001101101" => rgb <= "000000";
					when "01100001001101110" => rgb <= "000000";
					when "01100001001101111" => rgb <= "000000";
					when "01100001001110000" => rgb <= "000000";
					when "01100001001110001" => rgb <= "000000";
					when "01100001001110010" => rgb <= "000000";
					when "01100001001110011" => rgb <= "000000";
					when "01100001001110100" => rgb <= "000000";
					when "01100001001110101" => rgb <= "000000";
					when "01100001001110110" => rgb <= "000000";
					when "01100001001110111" => rgb <= "000000";
					when "01100001001111000" => rgb <= "000000";
					when "01100001001111001" => rgb <= "000000";
					when "01100001001111010" => rgb <= "000000";
					when "01100001001111011" => rgb <= "000000";
					when "01100001001111100" => rgb <= "000000";
					when "01100001001111101" => rgb <= "000000";
					when "01100001001111110" => rgb <= "000000";
					when "01100001001111111" => rgb <= "000000";
					when "01100001010000000" => rgb <= "000000";
					when "01100001010000001" => rgb <= "000000";
					when "01100001010000010" => rgb <= "000000";
					when "01100001010000011" => rgb <= "000000";
					when "01100001010000100" => rgb <= "000000";
					when "01100001010000101" => rgb <= "000000";
					when "01100001010000110" => rgb <= "000000";
					when "01100001010000111" => rgb <= "000000";
					when "01100001010001000" => rgb <= "000000";
					when "01100001010001001" => rgb <= "000000";
					when "01100001010001010" => rgb <= "000000";
					when "01100001010001011" => rgb <= "000000";
					when "01100001010001100" => rgb <= "000000";
					when "01100001010001101" => rgb <= "000000";
					when "01100001010001110" => rgb <= "000000";
					when "01100001010001111" => rgb <= "000000";
					when "01100001010010000" => rgb <= "000000";
					when "01100001010010001" => rgb <= "000000";
					when "01100001010010010" => rgb <= "000000";
					when "01100001010010011" => rgb <= "010000";
					when "01100001010010100" => rgb <= "101000";
					when "01100001010010101" => rgb <= "101000";
					when "01100001010010110" => rgb <= "101000";
					when "01100001010010111" => rgb <= "101000";
					when "01100001010011000" => rgb <= "101000";
					when "01100001010011001" => rgb <= "101000";
					when "01100001010011010" => rgb <= "101000";
					when "01100001010011011" => rgb <= "101000";
					when "01100001010011100" => rgb <= "101000";
					when "01100001010011101" => rgb <= "101000";
					when "01100001010011110" => rgb <= "101000";
					when "01100001010011111" => rgb <= "101000";
					when "01100001010100000" => rgb <= "101000";
					when "01100001010100001" => rgb <= "101000";
					when "01100001010100010" => rgb <= "101000";
					when "01100001010100011" => rgb <= "101000";
					when "01100001010100100" => rgb <= "101000";
					when "01100001010100101" => rgb <= "101000";
					when "01100001010100110" => rgb <= "101000";
					when "01100001010100111" => rgb <= "101000";
					when "01100001010101000" => rgb <= "101000";
					when "01100001010101001" => rgb <= "101000";
					when "01100001010101010" => rgb <= "010000";
					when "01100001010101011" => rgb <= "000000";
					when "01100001010101100" => rgb <= "000000";
					when "01100001010101101" => rgb <= "000000";
					when "01100001010101110" => rgb <= "000000";
					when "01100001010101111" => rgb <= "000000";
					when "01100001010110000" => rgb <= "000000";
					when "01100001010110001" => rgb <= "000000";
					when "01100001010110010" => rgb <= "000000";
					when "01100001010110011" => rgb <= "000000";
					when "01100001010110100" => rgb <= "000000";
					when "01100001010110101" => rgb <= "000000";
					when "01100001010110110" => rgb <= "000000";
					when "01100001010110111" => rgb <= "000000";
					when "01100001010111000" => rgb <= "000000";
					when "01100001010111001" => rgb <= "000000";
					when "01100001010111010" => rgb <= "000000";
					when "01100001010111011" => rgb <= "000000";
					when "01100001010111100" => rgb <= "000000";
					when "01100001010111101" => rgb <= "000000";
					when "01100001010111110" => rgb <= "000000";
					when "01100001010111111" => rgb <= "000000";
					when "01100001011000000" => rgb <= "000000";
					when "01100001011000001" => rgb <= "000000";
					when "01100001011000010" => rgb <= "000000";
					when "01100001011000011" => rgb <= "000000";
					when "01100001011000100" => rgb <= "000000";
					when "01100001011000101" => rgb <= "000000";
					when "01100001011000110" => rgb <= "000000";
					when "01100001011000111" => rgb <= "000000";
					when "01100001011001000" => rgb <= "000000";
					when "01100001011001001" => rgb <= "000000";
					when "01100001011001010" => rgb <= "000000";
					when "01100001011001011" => rgb <= "000000";
					when "01100001011001100" => rgb <= "000000";
					when "01100001011001101" => rgb <= "000000";
					when "01100001011001110" => rgb <= "000000";
					when "01100001011001111" => rgb <= "000000";
					when "01100001011010000" => rgb <= "000000";
					when "01100001011010001" => rgb <= "000000";
					when "01100001011010010" => rgb <= "000000";
					when "01100001011010011" => rgb <= "000000";
					when "01100001011010100" => rgb <= "000000";
					when "01100001011010101" => rgb <= "000000";
					when "01100001011010110" => rgb <= "000000";
					when "01100001011010111" => rgb <= "000000";
					when "01100001011011000" => rgb <= "000000";
					when "01100001011011001" => rgb <= "000000";
					when "01100001011011010" => rgb <= "000000";
					when "01100001011011011" => rgb <= "000000";
					when "01100001011011100" => rgb <= "000000";
					when "01100001011011101" => rgb <= "000000";
					when "01100001011011110" => rgb <= "000000";
					when "01100001011011111" => rgb <= "000000";
					when "01100001011100000" => rgb <= "000000";
					when "01100001011100001" => rgb <= "000000";
					when "01100001011100010" => rgb <= "000000";
					when "01100001011100011" => rgb <= "000000";
					when "01100001011100100" => rgb <= "000000";
					when "01100001011100101" => rgb <= "000000";
					when "01100001011100110" => rgb <= "000000";
					when "01100001011100111" => rgb <= "000000";
					when "01100001011101000" => rgb <= "000000";
					when "01100001011101001" => rgb <= "000000";
					when "01100001011101010" => rgb <= "000000";
					when "01100001011101011" => rgb <= "000000";
					when "01100001011101100" => rgb <= "000000";
					when "01100001011101101" => rgb <= "000000";
					when "01100001011101110" => rgb <= "000000";
					when "01100001011101111" => rgb <= "000000";
					when "01100001011110000" => rgb <= "000000";
					when "01100001011110001" => rgb <= "000000";
					when "01100001011110010" => rgb <= "000000";
					when "01100001011110011" => rgb <= "000000";
					when "01100001011110100" => rgb <= "000000";
					when "01100001011110101" => rgb <= "000000";
					when "01100001011110110" => rgb <= "000000";
					when "01100001011110111" => rgb <= "000000";
					when "01100001011111000" => rgb <= "000000";
					when "01100001011111001" => rgb <= "000000";
					when "01100001011111010" => rgb <= "000000";
					when "01100001011111011" => rgb <= "000000";
					when "01100001011111100" => rgb <= "000000";
					when "01100001011111101" => rgb <= "000000";
					when "01100001011111110" => rgb <= "000000";
					when "01100001011111111" => rgb <= "000000";
					when "01100001100000000" => rgb <= "000000";
					when "01100001100000001" => rgb <= "000000";
					when "01100001100000010" => rgb <= "000000";
					when "01100001100000011" => rgb <= "000000";
					when "01100001100000100" => rgb <= "000000";
					when "01100001100000101" => rgb <= "000000";
					when "01100001100000110" => rgb <= "000000";
					when "01100001100000111" => rgb <= "000000";
					when "01100001100001000" => rgb <= "000000";
					when "01100001100001001" => rgb <= "000000";
					when "01100001100001010" => rgb <= "000000";
					when "01100001100001011" => rgb <= "000000";
					when "01100001100001100" => rgb <= "000000";
					when "01100001100001101" => rgb <= "000000";
					when "01100001100001110" => rgb <= "000000";
					when "01100001100001111" => rgb <= "000000";
					when "01100001100010000" => rgb <= "000000";
					when "01100001100010001" => rgb <= "000000";
					when "01100001100010010" => rgb <= "000000";
					when "01100001100010011" => rgb <= "000000";
					when "01100001100010100" => rgb <= "000000";
					when "01100001100010101" => rgb <= "000000";
					when "01100001100010110" => rgb <= "000000";
					when "01100001100010111" => rgb <= "000000";
					when "01100001100011000" => rgb <= "000000";
					when "01100001100011001" => rgb <= "000000";
					when "01100001100011010" => rgb <= "000000";
					when "01100001100011011" => rgb <= "000000";
					when "01100001100011100" => rgb <= "000000";
					when "01100001100011101" => rgb <= "000000";
					when "01100001100011110" => rgb <= "000000";
					when "01100001100011111" => rgb <= "000000";
					when "01100001100100000" => rgb <= "000000";
					when "01100001100100001" => rgb <= "000000";
					when "01100001100100010" => rgb <= "000000";
					when "01100001100100011" => rgb <= "000000";
					when "01100001100100100" => rgb <= "000000";
					when "01100001100100101" => rgb <= "000000";
					when "01100001100100110" => rgb <= "000000";
					when "01100001100100111" => rgb <= "000000";
					when "01100001100101000" => rgb <= "000000";
					when "01100001100101001" => rgb <= "000000";
					when "01100001100101010" => rgb <= "000000";
					when "01100001100101011" => rgb <= "000000";
					when "01100001100101100" => rgb <= "000000";
					when "01100001100101101" => rgb <= "000000";
					when "01100001100101110" => rgb <= "000000";
					when "01100001100101111" => rgb <= "000000";
					when "01100001100110000" => rgb <= "000000";
					when "01100001100110001" => rgb <= "000000";
					when "01100001100110010" => rgb <= "000000";
					when "01100001100110011" => rgb <= "000000";
					when "01100001100110100" => rgb <= "000000";
					when "01100001100110101" => rgb <= "000000";
					when "01100001100110110" => rgb <= "000000";
					when "01100001100110111" => rgb <= "000000";
					when "01100001100111000" => rgb <= "000000";
					when "01100001100111001" => rgb <= "000000";
					when "01100001100111010" => rgb <= "000000";
					when "01100001100111011" => rgb <= "000000";
					when "01100001100111100" => rgb <= "000000";
					when "01100001100111101" => rgb <= "000000";
					when "01100001100111110" => rgb <= "000000";
					when "01100001100111111" => rgb <= "000000";
					when "01100010000000000" => rgb <= "000000";
					when "01100010000000001" => rgb <= "000000";
					when "01100010000000010" => rgb <= "000000";
					when "01100010000000011" => rgb <= "000000";
					when "01100010000000100" => rgb <= "000000";
					when "01100010000000101" => rgb <= "000000";
					when "01100010000000110" => rgb <= "000000";
					when "01100010000000111" => rgb <= "000000";
					when "01100010000001000" => rgb <= "000000";
					when "01100010000001001" => rgb <= "000000";
					when "01100010000001010" => rgb <= "000000";
					when "01100010000001011" => rgb <= "000000";
					when "01100010000001100" => rgb <= "000000";
					when "01100010000001101" => rgb <= "000000";
					when "01100010000001110" => rgb <= "000000";
					when "01100010000001111" => rgb <= "000000";
					when "01100010000010000" => rgb <= "000000";
					when "01100010000010001" => rgb <= "000000";
					when "01100010000010010" => rgb <= "000000";
					when "01100010000010011" => rgb <= "000000";
					when "01100010000010100" => rgb <= "000000";
					when "01100010000010101" => rgb <= "000000";
					when "01100010000010110" => rgb <= "000000";
					when "01100010000010111" => rgb <= "000000";
					when "01100010000011000" => rgb <= "000000";
					when "01100010000011001" => rgb <= "000000";
					when "01100010000011010" => rgb <= "000000";
					when "01100010000011011" => rgb <= "000000";
					when "01100010000011100" => rgb <= "000000";
					when "01100010000011101" => rgb <= "000000";
					when "01100010000011110" => rgb <= "000000";
					when "01100010000011111" => rgb <= "000000";
					when "01100010000100000" => rgb <= "000000";
					when "01100010000100001" => rgb <= "000000";
					when "01100010000100010" => rgb <= "000000";
					when "01100010000100011" => rgb <= "000000";
					when "01100010000100100" => rgb <= "000000";
					when "01100010000100101" => rgb <= "000000";
					when "01100010000100110" => rgb <= "000000";
					when "01100010000100111" => rgb <= "000000";
					when "01100010000101000" => rgb <= "000000";
					when "01100010000101001" => rgb <= "000000";
					when "01100010000101010" => rgb <= "000000";
					when "01100010000101011" => rgb <= "000000";
					when "01100010000101100" => rgb <= "000000";
					when "01100010000101101" => rgb <= "000000";
					when "01100010000101110" => rgb <= "000000";
					when "01100010000101111" => rgb <= "000000";
					when "01100010000110000" => rgb <= "000000";
					when "01100010000110001" => rgb <= "000000";
					when "01100010000110010" => rgb <= "000000";
					when "01100010000110011" => rgb <= "000000";
					when "01100010000110100" => rgb <= "000000";
					when "01100010000110101" => rgb <= "000000";
					when "01100010000110110" => rgb <= "000000";
					when "01100010000110111" => rgb <= "000000";
					when "01100010000111000" => rgb <= "000000";
					when "01100010000111001" => rgb <= "000000";
					when "01100010000111010" => rgb <= "000000";
					when "01100010000111011" => rgb <= "000000";
					when "01100010000111100" => rgb <= "000000";
					when "01100010000111101" => rgb <= "000000";
					when "01100010000111110" => rgb <= "000000";
					when "01100010000111111" => rgb <= "000000";
					when "01100010001000000" => rgb <= "000000";
					when "01100010001000001" => rgb <= "000000";
					when "01100010001000010" => rgb <= "000000";
					when "01100010001000011" => rgb <= "000000";
					when "01100010001000100" => rgb <= "000000";
					when "01100010001000101" => rgb <= "000000";
					when "01100010001000110" => rgb <= "000000";
					when "01100010001000111" => rgb <= "000000";
					when "01100010001001000" => rgb <= "000000";
					when "01100010001001001" => rgb <= "000000";
					when "01100010001001010" => rgb <= "000000";
					when "01100010001001011" => rgb <= "000000";
					when "01100010001001100" => rgb <= "000000";
					when "01100010001001101" => rgb <= "000000";
					when "01100010001001110" => rgb <= "000000";
					when "01100010001001111" => rgb <= "000000";
					when "01100010001010000" => rgb <= "000000";
					when "01100010001010001" => rgb <= "000000";
					when "01100010001010010" => rgb <= "000000";
					when "01100010001010011" => rgb <= "000000";
					when "01100010001010100" => rgb <= "000000";
					when "01100010001010101" => rgb <= "000000";
					when "01100010001010110" => rgb <= "000000";
					when "01100010001010111" => rgb <= "000000";
					when "01100010001011000" => rgb <= "000000";
					when "01100010001011001" => rgb <= "000000";
					when "01100010001011010" => rgb <= "000000";
					when "01100010001011011" => rgb <= "000000";
					when "01100010001011100" => rgb <= "000000";
					when "01100010001011101" => rgb <= "000000";
					when "01100010001011110" => rgb <= "000000";
					when "01100010001011111" => rgb <= "000000";
					when "01100010001100000" => rgb <= "000000";
					when "01100010001100001" => rgb <= "000000";
					when "01100010001100010" => rgb <= "000000";
					when "01100010001100011" => rgb <= "000000";
					when "01100010001100100" => rgb <= "000000";
					when "01100010001100101" => rgb <= "000000";
					when "01100010001100110" => rgb <= "000000";
					when "01100010001100111" => rgb <= "000000";
					when "01100010001101000" => rgb <= "000000";
					when "01100010001101001" => rgb <= "000000";
					when "01100010001101010" => rgb <= "000000";
					when "01100010001101011" => rgb <= "000000";
					when "01100010001101100" => rgb <= "000000";
					when "01100010001101101" => rgb <= "000000";
					when "01100010001101110" => rgb <= "000000";
					when "01100010001101111" => rgb <= "000000";
					when "01100010001110000" => rgb <= "000000";
					when "01100010001110001" => rgb <= "000000";
					when "01100010001110010" => rgb <= "000000";
					when "01100010001110011" => rgb <= "000000";
					when "01100010001110100" => rgb <= "000000";
					when "01100010001110101" => rgb <= "000000";
					when "01100010001110110" => rgb <= "000000";
					when "01100010001110111" => rgb <= "000000";
					when "01100010001111000" => rgb <= "000000";
					when "01100010001111001" => rgb <= "000000";
					when "01100010001111010" => rgb <= "000000";
					when "01100010001111011" => rgb <= "000000";
					when "01100010001111100" => rgb <= "000000";
					when "01100010001111101" => rgb <= "000000";
					when "01100010001111110" => rgb <= "000000";
					when "01100010001111111" => rgb <= "000000";
					when "01100010010000000" => rgb <= "000000";
					when "01100010010000001" => rgb <= "000000";
					when "01100010010000010" => rgb <= "000000";
					when "01100010010000011" => rgb <= "000000";
					when "01100010010000100" => rgb <= "000000";
					when "01100010010000101" => rgb <= "000000";
					when "01100010010000110" => rgb <= "000000";
					when "01100010010000111" => rgb <= "000000";
					when "01100010010001000" => rgb <= "000000";
					when "01100010010001001" => rgb <= "000000";
					when "01100010010001010" => rgb <= "000000";
					when "01100010010001011" => rgb <= "000000";
					when "01100010010001100" => rgb <= "000000";
					when "01100010010001101" => rgb <= "000000";
					when "01100010010001110" => rgb <= "000000";
					when "01100010010001111" => rgb <= "000000";
					when "01100010010010000" => rgb <= "000000";
					when "01100010010010001" => rgb <= "000000";
					when "01100010010010010" => rgb <= "000000";
					when "01100010010010011" => rgb <= "010000";
					when "01100010010010100" => rgb <= "101000";
					when "01100010010010101" => rgb <= "101000";
					when "01100010010010110" => rgb <= "101000";
					when "01100010010010111" => rgb <= "101000";
					when "01100010010011000" => rgb <= "101000";
					when "01100010010011001" => rgb <= "101000";
					when "01100010010011010" => rgb <= "101000";
					when "01100010010011011" => rgb <= "101000";
					when "01100010010011100" => rgb <= "101000";
					when "01100010010011101" => rgb <= "101000";
					when "01100010010011110" => rgb <= "101000";
					when "01100010010011111" => rgb <= "101000";
					when "01100010010100000" => rgb <= "101000";
					when "01100010010100001" => rgb <= "101000";
					when "01100010010100010" => rgb <= "101000";
					when "01100010010100011" => rgb <= "101000";
					when "01100010010100100" => rgb <= "101000";
					when "01100010010100101" => rgb <= "101000";
					when "01100010010100110" => rgb <= "101000";
					when "01100010010100111" => rgb <= "101000";
					when "01100010010101000" => rgb <= "101000";
					when "01100010010101001" => rgb <= "101000";
					when "01100010010101010" => rgb <= "010000";
					when "01100010010101011" => rgb <= "000000";
					when "01100010010101100" => rgb <= "000000";
					when "01100010010101101" => rgb <= "000000";
					when "01100010010101110" => rgb <= "000000";
					when "01100010010101111" => rgb <= "000000";
					when "01100010010110000" => rgb <= "000000";
					when "01100010010110001" => rgb <= "000000";
					when "01100010010110010" => rgb <= "000000";
					when "01100010010110011" => rgb <= "000000";
					when "01100010010110100" => rgb <= "000000";
					when "01100010010110101" => rgb <= "000000";
					when "01100010010110110" => rgb <= "000000";
					when "01100010010110111" => rgb <= "000000";
					when "01100010010111000" => rgb <= "000000";
					when "01100010010111001" => rgb <= "000000";
					when "01100010010111010" => rgb <= "000000";
					when "01100010010111011" => rgb <= "000000";
					when "01100010010111100" => rgb <= "000000";
					when "01100010010111101" => rgb <= "000000";
					when "01100010010111110" => rgb <= "000000";
					when "01100010010111111" => rgb <= "000000";
					when "01100010011000000" => rgb <= "000000";
					when "01100010011000001" => rgb <= "000000";
					when "01100010011000010" => rgb <= "000000";
					when "01100010011000011" => rgb <= "000000";
					when "01100010011000100" => rgb <= "000000";
					when "01100010011000101" => rgb <= "000000";
					when "01100010011000110" => rgb <= "000000";
					when "01100010011000111" => rgb <= "000000";
					when "01100010011001000" => rgb <= "000000";
					when "01100010011001001" => rgb <= "000000";
					when "01100010011001010" => rgb <= "000000";
					when "01100010011001011" => rgb <= "000000";
					when "01100010011001100" => rgb <= "000000";
					when "01100010011001101" => rgb <= "000000";
					when "01100010011001110" => rgb <= "000000";
					when "01100010011001111" => rgb <= "000000";
					when "01100010011010000" => rgb <= "000000";
					when "01100010011010001" => rgb <= "000000";
					when "01100010011010010" => rgb <= "000000";
					when "01100010011010011" => rgb <= "000000";
					when "01100010011010100" => rgb <= "000000";
					when "01100010011010101" => rgb <= "000000";
					when "01100010011010110" => rgb <= "000000";
					when "01100010011010111" => rgb <= "000000";
					when "01100010011011000" => rgb <= "000000";
					when "01100010011011001" => rgb <= "000000";
					when "01100010011011010" => rgb <= "000000";
					when "01100010011011011" => rgb <= "000000";
					when "01100010011011100" => rgb <= "000000";
					when "01100010011011101" => rgb <= "000000";
					when "01100010011011110" => rgb <= "000000";
					when "01100010011011111" => rgb <= "000000";
					when "01100010011100000" => rgb <= "000000";
					when "01100010011100001" => rgb <= "000000";
					when "01100010011100010" => rgb <= "000000";
					when "01100010011100011" => rgb <= "000000";
					when "01100010011100100" => rgb <= "000000";
					when "01100010011100101" => rgb <= "000000";
					when "01100010011100110" => rgb <= "000000";
					when "01100010011100111" => rgb <= "000000";
					when "01100010011101000" => rgb <= "000000";
					when "01100010011101001" => rgb <= "000000";
					when "01100010011101010" => rgb <= "000000";
					when "01100010011101011" => rgb <= "000000";
					when "01100010011101100" => rgb <= "000000";
					when "01100010011101101" => rgb <= "000000";
					when "01100010011101110" => rgb <= "000000";
					when "01100010011101111" => rgb <= "000000";
					when "01100010011110000" => rgb <= "000000";
					when "01100010011110001" => rgb <= "000000";
					when "01100010011110010" => rgb <= "000000";
					when "01100010011110011" => rgb <= "000000";
					when "01100010011110100" => rgb <= "000000";
					when "01100010011110101" => rgb <= "000000";
					when "01100010011110110" => rgb <= "000000";
					when "01100010011110111" => rgb <= "000000";
					when "01100010011111000" => rgb <= "000000";
					when "01100010011111001" => rgb <= "000000";
					when "01100010011111010" => rgb <= "000000";
					when "01100010011111011" => rgb <= "000000";
					when "01100010011111100" => rgb <= "000000";
					when "01100010011111101" => rgb <= "000000";
					when "01100010011111110" => rgb <= "000000";
					when "01100010011111111" => rgb <= "000000";
					when "01100010100000000" => rgb <= "000000";
					when "01100010100000001" => rgb <= "000000";
					when "01100010100000010" => rgb <= "000000";
					when "01100010100000011" => rgb <= "000000";
					when "01100010100000100" => rgb <= "000000";
					when "01100010100000101" => rgb <= "000000";
					when "01100010100000110" => rgb <= "000000";
					when "01100010100000111" => rgb <= "000000";
					when "01100010100001000" => rgb <= "000000";
					when "01100010100001001" => rgb <= "000000";
					when "01100010100001010" => rgb <= "000000";
					when "01100010100001011" => rgb <= "000000";
					when "01100010100001100" => rgb <= "000000";
					when "01100010100001101" => rgb <= "000000";
					when "01100010100001110" => rgb <= "000000";
					when "01100010100001111" => rgb <= "000000";
					when "01100010100010000" => rgb <= "000000";
					when "01100010100010001" => rgb <= "000000";
					when "01100010100010010" => rgb <= "000000";
					when "01100010100010011" => rgb <= "000000";
					when "01100010100010100" => rgb <= "000000";
					when "01100010100010101" => rgb <= "000000";
					when "01100010100010110" => rgb <= "000000";
					when "01100010100010111" => rgb <= "000000";
					when "01100010100011000" => rgb <= "000000";
					when "01100010100011001" => rgb <= "000000";
					when "01100010100011010" => rgb <= "000000";
					when "01100010100011011" => rgb <= "000000";
					when "01100010100011100" => rgb <= "000000";
					when "01100010100011101" => rgb <= "000000";
					when "01100010100011110" => rgb <= "000000";
					when "01100010100011111" => rgb <= "000000";
					when "01100010100100000" => rgb <= "000000";
					when "01100010100100001" => rgb <= "000000";
					when "01100010100100010" => rgb <= "000000";
					when "01100010100100011" => rgb <= "000000";
					when "01100010100100100" => rgb <= "000000";
					when "01100010100100101" => rgb <= "000000";
					when "01100010100100110" => rgb <= "000000";
					when "01100010100100111" => rgb <= "000000";
					when "01100010100101000" => rgb <= "000000";
					when "01100010100101001" => rgb <= "000000";
					when "01100010100101010" => rgb <= "000000";
					when "01100010100101011" => rgb <= "000000";
					when "01100010100101100" => rgb <= "000000";
					when "01100010100101101" => rgb <= "000000";
					when "01100010100101110" => rgb <= "000000";
					when "01100010100101111" => rgb <= "000000";
					when "01100010100110000" => rgb <= "000000";
					when "01100010100110001" => rgb <= "000000";
					when "01100010100110010" => rgb <= "000000";
					when "01100010100110011" => rgb <= "000000";
					when "01100010100110100" => rgb <= "000000";
					when "01100010100110101" => rgb <= "000000";
					when "01100010100110110" => rgb <= "000000";
					when "01100010100110111" => rgb <= "000000";
					when "01100010100111000" => rgb <= "000000";
					when "01100010100111001" => rgb <= "000000";
					when "01100010100111010" => rgb <= "000000";
					when "01100010100111011" => rgb <= "000000";
					when "01100010100111100" => rgb <= "000000";
					when "01100010100111101" => rgb <= "000000";
					when "01100010100111110" => rgb <= "000000";
					when "01100010100111111" => rgb <= "000000";
					when "01100011000000000" => rgb <= "000000";
					when "01100011000000001" => rgb <= "000000";
					when "01100011000000010" => rgb <= "000000";
					when "01100011000000011" => rgb <= "000000";
					when "01100011000000100" => rgb <= "000000";
					when "01100011000000101" => rgb <= "000000";
					when "01100011000000110" => rgb <= "000000";
					when "01100011000000111" => rgb <= "000000";
					when "01100011000001000" => rgb <= "000000";
					when "01100011000001001" => rgb <= "000000";
					when "01100011000001010" => rgb <= "000000";
					when "01100011000001011" => rgb <= "000000";
					when "01100011000001100" => rgb <= "000000";
					when "01100011000001101" => rgb <= "000000";
					when "01100011000001110" => rgb <= "000000";
					when "01100011000001111" => rgb <= "000000";
					when "01100011000010000" => rgb <= "000000";
					when "01100011000010001" => rgb <= "000000";
					when "01100011000010010" => rgb <= "000000";
					when "01100011000010011" => rgb <= "000000";
					when "01100011000010100" => rgb <= "000000";
					when "01100011000010101" => rgb <= "000000";
					when "01100011000010110" => rgb <= "000000";
					when "01100011000010111" => rgb <= "000000";
					when "01100011000011000" => rgb <= "000000";
					when "01100011000011001" => rgb <= "000000";
					when "01100011000011010" => rgb <= "000000";
					when "01100011000011011" => rgb <= "000000";
					when "01100011000011100" => rgb <= "000000";
					when "01100011000011101" => rgb <= "000000";
					when "01100011000011110" => rgb <= "000000";
					when "01100011000011111" => rgb <= "000000";
					when "01100011000100000" => rgb <= "000000";
					when "01100011000100001" => rgb <= "000000";
					when "01100011000100010" => rgb <= "000000";
					when "01100011000100011" => rgb <= "000000";
					when "01100011000100100" => rgb <= "000000";
					when "01100011000100101" => rgb <= "000000";
					when "01100011000100110" => rgb <= "000000";
					when "01100011000100111" => rgb <= "000000";
					when "01100011000101000" => rgb <= "000000";
					when "01100011000101001" => rgb <= "000000";
					when "01100011000101010" => rgb <= "000000";
					when "01100011000101011" => rgb <= "000000";
					when "01100011000101100" => rgb <= "000000";
					when "01100011000101101" => rgb <= "000000";
					when "01100011000101110" => rgb <= "000000";
					when "01100011000101111" => rgb <= "000000";
					when "01100011000110000" => rgb <= "000000";
					when "01100011000110001" => rgb <= "000000";
					when "01100011000110010" => rgb <= "000000";
					when "01100011000110011" => rgb <= "000000";
					when "01100011000110100" => rgb <= "000000";
					when "01100011000110101" => rgb <= "000000";
					when "01100011000110110" => rgb <= "000000";
					when "01100011000110111" => rgb <= "000000";
					when "01100011000111000" => rgb <= "000000";
					when "01100011000111001" => rgb <= "000000";
					when "01100011000111010" => rgb <= "000000";
					when "01100011000111011" => rgb <= "000000";
					when "01100011000111100" => rgb <= "000000";
					when "01100011000111101" => rgb <= "000000";
					when "01100011000111110" => rgb <= "000000";
					when "01100011000111111" => rgb <= "000000";
					when "01100011001000000" => rgb <= "000000";
					when "01100011001000001" => rgb <= "000000";
					when "01100011001000010" => rgb <= "000000";
					when "01100011001000011" => rgb <= "000000";
					when "01100011001000100" => rgb <= "000000";
					when "01100011001000101" => rgb <= "000000";
					when "01100011001000110" => rgb <= "000000";
					when "01100011001000111" => rgb <= "000000";
					when "01100011001001000" => rgb <= "000000";
					when "01100011001001001" => rgb <= "000000";
					when "01100011001001010" => rgb <= "000000";
					when "01100011001001011" => rgb <= "000000";
					when "01100011001001100" => rgb <= "000000";
					when "01100011001001101" => rgb <= "000000";
					when "01100011001001110" => rgb <= "000000";
					when "01100011001001111" => rgb <= "000000";
					when "01100011001010000" => rgb <= "000000";
					when "01100011001010001" => rgb <= "000000";
					when "01100011001010010" => rgb <= "000000";
					when "01100011001010011" => rgb <= "000000";
					when "01100011001010100" => rgb <= "000000";
					when "01100011001010101" => rgb <= "000000";
					when "01100011001010110" => rgb <= "000000";
					when "01100011001010111" => rgb <= "000000";
					when "01100011001011000" => rgb <= "000000";
					when "01100011001011001" => rgb <= "000000";
					when "01100011001011010" => rgb <= "000000";
					when "01100011001011011" => rgb <= "000000";
					when "01100011001011100" => rgb <= "000000";
					when "01100011001011101" => rgb <= "000000";
					when "01100011001011110" => rgb <= "000000";
					when "01100011001011111" => rgb <= "000000";
					when "01100011001100000" => rgb <= "000000";
					when "01100011001100001" => rgb <= "000000";
					when "01100011001100010" => rgb <= "000000";
					when "01100011001100011" => rgb <= "000000";
					when "01100011001100100" => rgb <= "000000";
					when "01100011001100101" => rgb <= "000000";
					when "01100011001100110" => rgb <= "000000";
					when "01100011001100111" => rgb <= "000000";
					when "01100011001101000" => rgb <= "000000";
					when "01100011001101001" => rgb <= "000000";
					when "01100011001101010" => rgb <= "000000";
					when "01100011001101011" => rgb <= "000000";
					when "01100011001101100" => rgb <= "000000";
					when "01100011001101101" => rgb <= "000000";
					when "01100011001101110" => rgb <= "000000";
					when "01100011001101111" => rgb <= "000000";
					when "01100011001110000" => rgb <= "000000";
					when "01100011001110001" => rgb <= "000000";
					when "01100011001110010" => rgb <= "000000";
					when "01100011001110011" => rgb <= "000000";
					when "01100011001110100" => rgb <= "000000";
					when "01100011001110101" => rgb <= "000000";
					when "01100011001110110" => rgb <= "000000";
					when "01100011001110111" => rgb <= "000000";
					when "01100011001111000" => rgb <= "000000";
					when "01100011001111001" => rgb <= "000000";
					when "01100011001111010" => rgb <= "000000";
					when "01100011001111011" => rgb <= "000000";
					when "01100011001111100" => rgb <= "000000";
					when "01100011001111101" => rgb <= "000000";
					when "01100011001111110" => rgb <= "000000";
					when "01100011001111111" => rgb <= "000000";
					when "01100011010000000" => rgb <= "000000";
					when "01100011010000001" => rgb <= "000000";
					when "01100011010000010" => rgb <= "000000";
					when "01100011010000011" => rgb <= "000000";
					when "01100011010000100" => rgb <= "000000";
					when "01100011010000101" => rgb <= "000000";
					when "01100011010000110" => rgb <= "000000";
					when "01100011010000111" => rgb <= "000000";
					when "01100011010001000" => rgb <= "000000";
					when "01100011010001001" => rgb <= "000000";
					when "01100011010001010" => rgb <= "000000";
					when "01100011010001011" => rgb <= "000000";
					when "01100011010001100" => rgb <= "000000";
					when "01100011010001101" => rgb <= "000000";
					when "01100011010001110" => rgb <= "000000";
					when "01100011010001111" => rgb <= "000000";
					when "01100011010010000" => rgb <= "000000";
					when "01100011010010001" => rgb <= "000000";
					when "01100011010010010" => rgb <= "000000";
					when "01100011010010011" => rgb <= "010000";
					when "01100011010010100" => rgb <= "101000";
					when "01100011010010101" => rgb <= "101000";
					when "01100011010010110" => rgb <= "101000";
					when "01100011010010111" => rgb <= "101000";
					when "01100011010011000" => rgb <= "101000";
					when "01100011010011001" => rgb <= "101000";
					when "01100011010011010" => rgb <= "101000";
					when "01100011010011011" => rgb <= "101000";
					when "01100011010011100" => rgb <= "101000";
					when "01100011010011101" => rgb <= "101000";
					when "01100011010011110" => rgb <= "101000";
					when "01100011010011111" => rgb <= "101000";
					when "01100011010100000" => rgb <= "101000";
					when "01100011010100001" => rgb <= "101000";
					when "01100011010100010" => rgb <= "101000";
					when "01100011010100011" => rgb <= "101000";
					when "01100011010100100" => rgb <= "101000";
					when "01100011010100101" => rgb <= "101000";
					when "01100011010100110" => rgb <= "101000";
					when "01100011010100111" => rgb <= "101000";
					when "01100011010101000" => rgb <= "101000";
					when "01100011010101001" => rgb <= "101000";
					when "01100011010101010" => rgb <= "010000";
					when "01100011010101011" => rgb <= "000000";
					when "01100011010101100" => rgb <= "000000";
					when "01100011010101101" => rgb <= "000000";
					when "01100011010101110" => rgb <= "000000";
					when "01100011010101111" => rgb <= "000000";
					when "01100011010110000" => rgb <= "000000";
					when "01100011010110001" => rgb <= "000000";
					when "01100011010110010" => rgb <= "000000";
					when "01100011010110011" => rgb <= "000000";
					when "01100011010110100" => rgb <= "000000";
					when "01100011010110101" => rgb <= "000000";
					when "01100011010110110" => rgb <= "000000";
					when "01100011010110111" => rgb <= "000000";
					when "01100011010111000" => rgb <= "000000";
					when "01100011010111001" => rgb <= "000000";
					when "01100011010111010" => rgb <= "000000";
					when "01100011010111011" => rgb <= "000000";
					when "01100011010111100" => rgb <= "000000";
					when "01100011010111101" => rgb <= "000000";
					when "01100011010111110" => rgb <= "000000";
					when "01100011010111111" => rgb <= "000000";
					when "01100011011000000" => rgb <= "000000";
					when "01100011011000001" => rgb <= "000000";
					when "01100011011000010" => rgb <= "000000";
					when "01100011011000011" => rgb <= "000000";
					when "01100011011000100" => rgb <= "000000";
					when "01100011011000101" => rgb <= "000000";
					when "01100011011000110" => rgb <= "000000";
					when "01100011011000111" => rgb <= "000000";
					when "01100011011001000" => rgb <= "000000";
					when "01100011011001001" => rgb <= "000000";
					when "01100011011001010" => rgb <= "000000";
					when "01100011011001011" => rgb <= "000000";
					when "01100011011001100" => rgb <= "000000";
					when "01100011011001101" => rgb <= "000000";
					when "01100011011001110" => rgb <= "000000";
					when "01100011011001111" => rgb <= "000000";
					when "01100011011010000" => rgb <= "000000";
					when "01100011011010001" => rgb <= "000000";
					when "01100011011010010" => rgb <= "000000";
					when "01100011011010011" => rgb <= "000000";
					when "01100011011010100" => rgb <= "000000";
					when "01100011011010101" => rgb <= "000000";
					when "01100011011010110" => rgb <= "000000";
					when "01100011011010111" => rgb <= "000000";
					when "01100011011011000" => rgb <= "000000";
					when "01100011011011001" => rgb <= "000000";
					when "01100011011011010" => rgb <= "000000";
					when "01100011011011011" => rgb <= "000000";
					when "01100011011011100" => rgb <= "000000";
					when "01100011011011101" => rgb <= "000000";
					when "01100011011011110" => rgb <= "000000";
					when "01100011011011111" => rgb <= "000000";
					when "01100011011100000" => rgb <= "000000";
					when "01100011011100001" => rgb <= "000000";
					when "01100011011100010" => rgb <= "000000";
					when "01100011011100011" => rgb <= "000000";
					when "01100011011100100" => rgb <= "000000";
					when "01100011011100101" => rgb <= "000000";
					when "01100011011100110" => rgb <= "000000";
					when "01100011011100111" => rgb <= "000000";
					when "01100011011101000" => rgb <= "000000";
					when "01100011011101001" => rgb <= "000000";
					when "01100011011101010" => rgb <= "000000";
					when "01100011011101011" => rgb <= "000000";
					when "01100011011101100" => rgb <= "000000";
					when "01100011011101101" => rgb <= "000000";
					when "01100011011101110" => rgb <= "000000";
					when "01100011011101111" => rgb <= "000000";
					when "01100011011110000" => rgb <= "000000";
					when "01100011011110001" => rgb <= "000000";
					when "01100011011110010" => rgb <= "000000";
					when "01100011011110011" => rgb <= "000000";
					when "01100011011110100" => rgb <= "000000";
					when "01100011011110101" => rgb <= "000000";
					when "01100011011110110" => rgb <= "000000";
					when "01100011011110111" => rgb <= "000000";
					when "01100011011111000" => rgb <= "000000";
					when "01100011011111001" => rgb <= "000000";
					when "01100011011111010" => rgb <= "000000";
					when "01100011011111011" => rgb <= "000000";
					when "01100011011111100" => rgb <= "000000";
					when "01100011011111101" => rgb <= "000000";
					when "01100011011111110" => rgb <= "000000";
					when "01100011011111111" => rgb <= "000000";
					when "01100011100000000" => rgb <= "000000";
					when "01100011100000001" => rgb <= "000000";
					when "01100011100000010" => rgb <= "000000";
					when "01100011100000011" => rgb <= "000000";
					when "01100011100000100" => rgb <= "000000";
					when "01100011100000101" => rgb <= "000000";
					when "01100011100000110" => rgb <= "000000";
					when "01100011100000111" => rgb <= "000000";
					when "01100011100001000" => rgb <= "000000";
					when "01100011100001001" => rgb <= "000000";
					when "01100011100001010" => rgb <= "000000";
					when "01100011100001011" => rgb <= "000000";
					when "01100011100001100" => rgb <= "000000";
					when "01100011100001101" => rgb <= "000000";
					when "01100011100001110" => rgb <= "000000";
					when "01100011100001111" => rgb <= "000000";
					when "01100011100010000" => rgb <= "000000";
					when "01100011100010001" => rgb <= "000000";
					when "01100011100010010" => rgb <= "000000";
					when "01100011100010011" => rgb <= "000000";
					when "01100011100010100" => rgb <= "000000";
					when "01100011100010101" => rgb <= "000000";
					when "01100011100010110" => rgb <= "000000";
					when "01100011100010111" => rgb <= "000000";
					when "01100011100011000" => rgb <= "000000";
					when "01100011100011001" => rgb <= "000000";
					when "01100011100011010" => rgb <= "000000";
					when "01100011100011011" => rgb <= "000000";
					when "01100011100011100" => rgb <= "000000";
					when "01100011100011101" => rgb <= "000000";
					when "01100011100011110" => rgb <= "000000";
					when "01100011100011111" => rgb <= "000000";
					when "01100011100100000" => rgb <= "000000";
					when "01100011100100001" => rgb <= "000000";
					when "01100011100100010" => rgb <= "000000";
					when "01100011100100011" => rgb <= "000000";
					when "01100011100100100" => rgb <= "000000";
					when "01100011100100101" => rgb <= "000000";
					when "01100011100100110" => rgb <= "000000";
					when "01100011100100111" => rgb <= "000000";
					when "01100011100101000" => rgb <= "000000";
					when "01100011100101001" => rgb <= "000000";
					when "01100011100101010" => rgb <= "000000";
					when "01100011100101011" => rgb <= "000000";
					when "01100011100101100" => rgb <= "000000";
					when "01100011100101101" => rgb <= "000000";
					when "01100011100101110" => rgb <= "000000";
					when "01100011100101111" => rgb <= "000000";
					when "01100011100110000" => rgb <= "000000";
					when "01100011100110001" => rgb <= "000000";
					when "01100011100110010" => rgb <= "000000";
					when "01100011100110011" => rgb <= "000000";
					when "01100011100110100" => rgb <= "000000";
					when "01100011100110101" => rgb <= "000000";
					when "01100011100110110" => rgb <= "000000";
					when "01100011100110111" => rgb <= "000000";
					when "01100011100111000" => rgb <= "000000";
					when "01100011100111001" => rgb <= "000000";
					when "01100011100111010" => rgb <= "000000";
					when "01100011100111011" => rgb <= "000000";
					when "01100011100111100" => rgb <= "000000";
					when "01100011100111101" => rgb <= "000000";
					when "01100011100111110" => rgb <= "000000";
					when "01100011100111111" => rgb <= "000000";
					when "01100100000000000" => rgb <= "000000";
					when "01100100000000001" => rgb <= "000000";
					when "01100100000000010" => rgb <= "000000";
					when "01100100000000011" => rgb <= "000000";
					when "01100100000000100" => rgb <= "000000";
					when "01100100000000101" => rgb <= "000000";
					when "01100100000000110" => rgb <= "000000";
					when "01100100000000111" => rgb <= "000000";
					when "01100100000001000" => rgb <= "000000";
					when "01100100000001001" => rgb <= "000000";
					when "01100100000001010" => rgb <= "000000";
					when "01100100000001011" => rgb <= "000000";
					when "01100100000001100" => rgb <= "000000";
					when "01100100000001101" => rgb <= "000000";
					when "01100100000001110" => rgb <= "000000";
					when "01100100000001111" => rgb <= "000000";
					when "01100100000010000" => rgb <= "000000";
					when "01100100000010001" => rgb <= "000000";
					when "01100100000010010" => rgb <= "000000";
					when "01100100000010011" => rgb <= "000000";
					when "01100100000010100" => rgb <= "000000";
					when "01100100000010101" => rgb <= "000000";
					when "01100100000010110" => rgb <= "000000";
					when "01100100000010111" => rgb <= "000000";
					when "01100100000011000" => rgb <= "000000";
					when "01100100000011001" => rgb <= "000000";
					when "01100100000011010" => rgb <= "000000";
					when "01100100000011011" => rgb <= "000000";
					when "01100100000011100" => rgb <= "000000";
					when "01100100000011101" => rgb <= "000000";
					when "01100100000011110" => rgb <= "000000";
					when "01100100000011111" => rgb <= "000000";
					when "01100100000100000" => rgb <= "000000";
					when "01100100000100001" => rgb <= "000000";
					when "01100100000100010" => rgb <= "000000";
					when "01100100000100011" => rgb <= "000000";
					when "01100100000100100" => rgb <= "000000";
					when "01100100000100101" => rgb <= "000000";
					when "01100100000100110" => rgb <= "000000";
					when "01100100000100111" => rgb <= "000000";
					when "01100100000101000" => rgb <= "000000";
					when "01100100000101001" => rgb <= "000000";
					when "01100100000101010" => rgb <= "000000";
					when "01100100000101011" => rgb <= "000000";
					when "01100100000101100" => rgb <= "000000";
					when "01100100000101101" => rgb <= "000000";
					when "01100100000101110" => rgb <= "000000";
					when "01100100000101111" => rgb <= "000000";
					when "01100100000110000" => rgb <= "000000";
					when "01100100000110001" => rgb <= "000000";
					when "01100100000110010" => rgb <= "000000";
					when "01100100000110011" => rgb <= "000000";
					when "01100100000110100" => rgb <= "000000";
					when "01100100000110101" => rgb <= "000000";
					when "01100100000110110" => rgb <= "000000";
					when "01100100000110111" => rgb <= "000000";
					when "01100100000111000" => rgb <= "000000";
					when "01100100000111001" => rgb <= "000000";
					when "01100100000111010" => rgb <= "000000";
					when "01100100000111011" => rgb <= "000000";
					when "01100100000111100" => rgb <= "000000";
					when "01100100000111101" => rgb <= "000000";
					when "01100100000111110" => rgb <= "000000";
					when "01100100000111111" => rgb <= "000000";
					when "01100100001000000" => rgb <= "000000";
					when "01100100001000001" => rgb <= "000000";
					when "01100100001000010" => rgb <= "000000";
					when "01100100001000011" => rgb <= "000000";
					when "01100100001000100" => rgb <= "000000";
					when "01100100001000101" => rgb <= "000000";
					when "01100100001000110" => rgb <= "000000";
					when "01100100001000111" => rgb <= "000000";
					when "01100100001001000" => rgb <= "000000";
					when "01100100001001001" => rgb <= "000000";
					when "01100100001001010" => rgb <= "000000";
					when "01100100001001011" => rgb <= "000000";
					when "01100100001001100" => rgb <= "000000";
					when "01100100001001101" => rgb <= "000000";
					when "01100100001001110" => rgb <= "000000";
					when "01100100001001111" => rgb <= "000000";
					when "01100100001010000" => rgb <= "000000";
					when "01100100001010001" => rgb <= "000000";
					when "01100100001010010" => rgb <= "000000";
					when "01100100001010011" => rgb <= "000000";
					when "01100100001010100" => rgb <= "000000";
					when "01100100001010101" => rgb <= "000000";
					when "01100100001010110" => rgb <= "000000";
					when "01100100001010111" => rgb <= "000000";
					when "01100100001011000" => rgb <= "000000";
					when "01100100001011001" => rgb <= "000000";
					when "01100100001011010" => rgb <= "000000";
					when "01100100001011011" => rgb <= "000000";
					when "01100100001011100" => rgb <= "000000";
					when "01100100001011101" => rgb <= "000000";
					when "01100100001011110" => rgb <= "000000";
					when "01100100001011111" => rgb <= "000000";
					when "01100100001100000" => rgb <= "000000";
					when "01100100001100001" => rgb <= "000000";
					when "01100100001100010" => rgb <= "000000";
					when "01100100001100011" => rgb <= "000000";
					when "01100100001100100" => rgb <= "000000";
					when "01100100001100101" => rgb <= "000000";
					when "01100100001100110" => rgb <= "000000";
					when "01100100001100111" => rgb <= "000000";
					when "01100100001101000" => rgb <= "000000";
					when "01100100001101001" => rgb <= "000000";
					when "01100100001101010" => rgb <= "000000";
					when "01100100001101011" => rgb <= "000000";
					when "01100100001101100" => rgb <= "000000";
					when "01100100001101101" => rgb <= "000000";
					when "01100100001101110" => rgb <= "000000";
					when "01100100001101111" => rgb <= "000000";
					when "01100100001110000" => rgb <= "000000";
					when "01100100001110001" => rgb <= "000000";
					when "01100100001110010" => rgb <= "000000";
					when "01100100001110011" => rgb <= "000000";
					when "01100100001110100" => rgb <= "000000";
					when "01100100001110101" => rgb <= "000000";
					when "01100100001110110" => rgb <= "000000";
					when "01100100001110111" => rgb <= "000000";
					when "01100100001111000" => rgb <= "000000";
					when "01100100001111001" => rgb <= "000000";
					when "01100100001111010" => rgb <= "000000";
					when "01100100001111011" => rgb <= "000000";
					when "01100100001111100" => rgb <= "000000";
					when "01100100001111101" => rgb <= "000000";
					when "01100100001111110" => rgb <= "000000";
					when "01100100001111111" => rgb <= "000000";
					when "01100100010000000" => rgb <= "000000";
					when "01100100010000001" => rgb <= "000000";
					when "01100100010000010" => rgb <= "000000";
					when "01100100010000011" => rgb <= "000000";
					when "01100100010000100" => rgb <= "000000";
					when "01100100010000101" => rgb <= "000000";
					when "01100100010000110" => rgb <= "000000";
					when "01100100010000111" => rgb <= "000000";
					when "01100100010001000" => rgb <= "000000";
					when "01100100010001001" => rgb <= "000000";
					when "01100100010001010" => rgb <= "000000";
					when "01100100010001011" => rgb <= "000000";
					when "01100100010001100" => rgb <= "000000";
					when "01100100010001101" => rgb <= "000000";
					when "01100100010001110" => rgb <= "000000";
					when "01100100010001111" => rgb <= "000000";
					when "01100100010010000" => rgb <= "000000";
					when "01100100010010001" => rgb <= "000000";
					when "01100100010010010" => rgb <= "000000";
					when "01100100010010011" => rgb <= "010000";
					when "01100100010010100" => rgb <= "101000";
					when "01100100010010101" => rgb <= "101000";
					when "01100100010010110" => rgb <= "101000";
					when "01100100010010111" => rgb <= "101000";
					when "01100100010011000" => rgb <= "101000";
					when "01100100010011001" => rgb <= "101000";
					when "01100100010011010" => rgb <= "101000";
					when "01100100010011011" => rgb <= "101000";
					when "01100100010011100" => rgb <= "101000";
					when "01100100010011101" => rgb <= "101000";
					when "01100100010011110" => rgb <= "101000";
					when "01100100010011111" => rgb <= "101000";
					when "01100100010100000" => rgb <= "101000";
					when "01100100010100001" => rgb <= "101000";
					when "01100100010100010" => rgb <= "101000";
					when "01100100010100011" => rgb <= "101000";
					when "01100100010100100" => rgb <= "101000";
					when "01100100010100101" => rgb <= "101000";
					when "01100100010100110" => rgb <= "101000";
					when "01100100010100111" => rgb <= "101000";
					when "01100100010101000" => rgb <= "101000";
					when "01100100010101001" => rgb <= "101000";
					when "01100100010101010" => rgb <= "010000";
					when "01100100010101011" => rgb <= "000000";
					when "01100100010101100" => rgb <= "000000";
					when "01100100010101101" => rgb <= "000000";
					when "01100100010101110" => rgb <= "000000";
					when "01100100010101111" => rgb <= "000000";
					when "01100100010110000" => rgb <= "000000";
					when "01100100010110001" => rgb <= "000000";
					when "01100100010110010" => rgb <= "000000";
					when "01100100010110011" => rgb <= "000000";
					when "01100100010110100" => rgb <= "000000";
					when "01100100010110101" => rgb <= "000000";
					when "01100100010110110" => rgb <= "000000";
					when "01100100010110111" => rgb <= "000000";
					when "01100100010111000" => rgb <= "000000";
					when "01100100010111001" => rgb <= "000000";
					when "01100100010111010" => rgb <= "000000";
					when "01100100010111011" => rgb <= "000000";
					when "01100100010111100" => rgb <= "000000";
					when "01100100010111101" => rgb <= "000000";
					when "01100100010111110" => rgb <= "000000";
					when "01100100010111111" => rgb <= "000000";
					when "01100100011000000" => rgb <= "000000";
					when "01100100011000001" => rgb <= "000000";
					when "01100100011000010" => rgb <= "000000";
					when "01100100011000011" => rgb <= "000000";
					when "01100100011000100" => rgb <= "000000";
					when "01100100011000101" => rgb <= "000000";
					when "01100100011000110" => rgb <= "000000";
					when "01100100011000111" => rgb <= "000000";
					when "01100100011001000" => rgb <= "000000";
					when "01100100011001001" => rgb <= "000000";
					when "01100100011001010" => rgb <= "000000";
					when "01100100011001011" => rgb <= "000000";
					when "01100100011001100" => rgb <= "000000";
					when "01100100011001101" => rgb <= "000000";
					when "01100100011001110" => rgb <= "000000";
					when "01100100011001111" => rgb <= "000000";
					when "01100100011010000" => rgb <= "000000";
					when "01100100011010001" => rgb <= "000000";
					when "01100100011010010" => rgb <= "000000";
					when "01100100011010011" => rgb <= "000000";
					when "01100100011010100" => rgb <= "000000";
					when "01100100011010101" => rgb <= "000000";
					when "01100100011010110" => rgb <= "000000";
					when "01100100011010111" => rgb <= "000000";
					when "01100100011011000" => rgb <= "000000";
					when "01100100011011001" => rgb <= "000000";
					when "01100100011011010" => rgb <= "000000";
					when "01100100011011011" => rgb <= "000000";
					when "01100100011011100" => rgb <= "000000";
					when "01100100011011101" => rgb <= "000000";
					when "01100100011011110" => rgb <= "000000";
					when "01100100011011111" => rgb <= "000000";
					when "01100100011100000" => rgb <= "000000";
					when "01100100011100001" => rgb <= "000000";
					when "01100100011100010" => rgb <= "000000";
					when "01100100011100011" => rgb <= "000000";
					when "01100100011100100" => rgb <= "000000";
					when "01100100011100101" => rgb <= "000000";
					when "01100100011100110" => rgb <= "000000";
					when "01100100011100111" => rgb <= "000000";
					when "01100100011101000" => rgb <= "000000";
					when "01100100011101001" => rgb <= "000000";
					when "01100100011101010" => rgb <= "000000";
					when "01100100011101011" => rgb <= "000000";
					when "01100100011101100" => rgb <= "000000";
					when "01100100011101101" => rgb <= "000000";
					when "01100100011101110" => rgb <= "000000";
					when "01100100011101111" => rgb <= "000000";
					when "01100100011110000" => rgb <= "000000";
					when "01100100011110001" => rgb <= "000000";
					when "01100100011110010" => rgb <= "000000";
					when "01100100011110011" => rgb <= "000000";
					when "01100100011110100" => rgb <= "000000";
					when "01100100011110101" => rgb <= "000000";
					when "01100100011110110" => rgb <= "000000";
					when "01100100011110111" => rgb <= "000000";
					when "01100100011111000" => rgb <= "000000";
					when "01100100011111001" => rgb <= "000000";
					when "01100100011111010" => rgb <= "000000";
					when "01100100011111011" => rgb <= "000000";
					when "01100100011111100" => rgb <= "000000";
					when "01100100011111101" => rgb <= "000000";
					when "01100100011111110" => rgb <= "000000";
					when "01100100011111111" => rgb <= "000000";
					when "01100100100000000" => rgb <= "000000";
					when "01100100100000001" => rgb <= "000000";
					when "01100100100000010" => rgb <= "000000";
					when "01100100100000011" => rgb <= "000000";
					when "01100100100000100" => rgb <= "000000";
					when "01100100100000101" => rgb <= "000000";
					when "01100100100000110" => rgb <= "000000";
					when "01100100100000111" => rgb <= "000000";
					when "01100100100001000" => rgb <= "000000";
					when "01100100100001001" => rgb <= "000000";
					when "01100100100001010" => rgb <= "000000";
					when "01100100100001011" => rgb <= "000000";
					when "01100100100001100" => rgb <= "000000";
					when "01100100100001101" => rgb <= "000000";
					when "01100100100001110" => rgb <= "000000";
					when "01100100100001111" => rgb <= "000000";
					when "01100100100010000" => rgb <= "000000";
					when "01100100100010001" => rgb <= "000000";
					when "01100100100010010" => rgb <= "000000";
					when "01100100100010011" => rgb <= "000000";
					when "01100100100010100" => rgb <= "000000";
					when "01100100100010101" => rgb <= "000000";
					when "01100100100010110" => rgb <= "000000";
					when "01100100100010111" => rgb <= "000000";
					when "01100100100011000" => rgb <= "000000";
					when "01100100100011001" => rgb <= "000000";
					when "01100100100011010" => rgb <= "000000";
					when "01100100100011011" => rgb <= "000000";
					when "01100100100011100" => rgb <= "000000";
					when "01100100100011101" => rgb <= "000000";
					when "01100100100011110" => rgb <= "000000";
					when "01100100100011111" => rgb <= "000000";
					when "01100100100100000" => rgb <= "000000";
					when "01100100100100001" => rgb <= "000000";
					when "01100100100100010" => rgb <= "000000";
					when "01100100100100011" => rgb <= "000000";
					when "01100100100100100" => rgb <= "000000";
					when "01100100100100101" => rgb <= "000000";
					when "01100100100100110" => rgb <= "000000";
					when "01100100100100111" => rgb <= "000000";
					when "01100100100101000" => rgb <= "000000";
					when "01100100100101001" => rgb <= "000000";
					when "01100100100101010" => rgb <= "000000";
					when "01100100100101011" => rgb <= "000000";
					when "01100100100101100" => rgb <= "000000";
					when "01100100100101101" => rgb <= "000000";
					when "01100100100101110" => rgb <= "000000";
					when "01100100100101111" => rgb <= "000000";
					when "01100100100110000" => rgb <= "000000";
					when "01100100100110001" => rgb <= "000000";
					when "01100100100110010" => rgb <= "000000";
					when "01100100100110011" => rgb <= "000000";
					when "01100100100110100" => rgb <= "000000";
					when "01100100100110101" => rgb <= "000000";
					when "01100100100110110" => rgb <= "000000";
					when "01100100100110111" => rgb <= "000000";
					when "01100100100111000" => rgb <= "000000";
					when "01100100100111001" => rgb <= "000000";
					when "01100100100111010" => rgb <= "000000";
					when "01100100100111011" => rgb <= "000000";
					when "01100100100111100" => rgb <= "000000";
					when "01100100100111101" => rgb <= "000000";
					when "01100100100111110" => rgb <= "000000";
					when "01100100100111111" => rgb <= "000000";
					when "01100101000000000" => rgb <= "000000";
					when "01100101000000001" => rgb <= "000000";
					when "01100101000000010" => rgb <= "000000";
					when "01100101000000011" => rgb <= "000000";
					when "01100101000000100" => rgb <= "000000";
					when "01100101000000101" => rgb <= "000000";
					when "01100101000000110" => rgb <= "000000";
					when "01100101000000111" => rgb <= "000000";
					when "01100101000001000" => rgb <= "000000";
					when "01100101000001001" => rgb <= "000000";
					when "01100101000001010" => rgb <= "000000";
					when "01100101000001011" => rgb <= "000000";
					when "01100101000001100" => rgb <= "000000";
					when "01100101000001101" => rgb <= "000000";
					when "01100101000001110" => rgb <= "000000";
					when "01100101000001111" => rgb <= "000000";
					when "01100101000010000" => rgb <= "000000";
					when "01100101000010001" => rgb <= "000000";
					when "01100101000010010" => rgb <= "000000";
					when "01100101000010011" => rgb <= "000000";
					when "01100101000010100" => rgb <= "000000";
					when "01100101000010101" => rgb <= "000000";
					when "01100101000010110" => rgb <= "000000";
					when "01100101000010111" => rgb <= "000000";
					when "01100101000011000" => rgb <= "000000";
					when "01100101000011001" => rgb <= "000000";
					when "01100101000011010" => rgb <= "000000";
					when "01100101000011011" => rgb <= "000000";
					when "01100101000011100" => rgb <= "000000";
					when "01100101000011101" => rgb <= "000000";
					when "01100101000011110" => rgb <= "000000";
					when "01100101000011111" => rgb <= "000000";
					when "01100101000100000" => rgb <= "000000";
					when "01100101000100001" => rgb <= "000000";
					when "01100101000100010" => rgb <= "000000";
					when "01100101000100011" => rgb <= "000000";
					when "01100101000100100" => rgb <= "000000";
					when "01100101000100101" => rgb <= "000000";
					when "01100101000100110" => rgb <= "000000";
					when "01100101000100111" => rgb <= "000000";
					when "01100101000101000" => rgb <= "000000";
					when "01100101000101001" => rgb <= "000000";
					when "01100101000101010" => rgb <= "000000";
					when "01100101000101011" => rgb <= "000000";
					when "01100101000101100" => rgb <= "000000";
					when "01100101000101101" => rgb <= "000000";
					when "01100101000101110" => rgb <= "000000";
					when "01100101000101111" => rgb <= "000000";
					when "01100101000110000" => rgb <= "000000";
					when "01100101000110001" => rgb <= "000000";
					when "01100101000110010" => rgb <= "000000";
					when "01100101000110011" => rgb <= "000000";
					when "01100101000110100" => rgb <= "000000";
					when "01100101000110101" => rgb <= "000000";
					when "01100101000110110" => rgb <= "000000";
					when "01100101000110111" => rgb <= "000000";
					when "01100101000111000" => rgb <= "000000";
					when "01100101000111001" => rgb <= "000000";
					when "01100101000111010" => rgb <= "000000";
					when "01100101000111011" => rgb <= "000000";
					when "01100101000111100" => rgb <= "000000";
					when "01100101000111101" => rgb <= "000000";
					when "01100101000111110" => rgb <= "000000";
					when "01100101000111111" => rgb <= "000000";
					when "01100101001000000" => rgb <= "000000";
					when "01100101001000001" => rgb <= "000000";
					when "01100101001000010" => rgb <= "000000";
					when "01100101001000011" => rgb <= "000000";
					when "01100101001000100" => rgb <= "000000";
					when "01100101001000101" => rgb <= "000000";
					when "01100101001000110" => rgb <= "000000";
					when "01100101001000111" => rgb <= "000000";
					when "01100101001001000" => rgb <= "000000";
					when "01100101001001001" => rgb <= "000000";
					when "01100101001001010" => rgb <= "000000";
					when "01100101001001011" => rgb <= "000000";
					when "01100101001001100" => rgb <= "000000";
					when "01100101001001101" => rgb <= "000000";
					when "01100101001001110" => rgb <= "000000";
					when "01100101001001111" => rgb <= "000000";
					when "01100101001010000" => rgb <= "000000";
					when "01100101001010001" => rgb <= "000000";
					when "01100101001010010" => rgb <= "000000";
					when "01100101001010011" => rgb <= "000000";
					when "01100101001010100" => rgb <= "000000";
					when "01100101001010101" => rgb <= "000000";
					when "01100101001010110" => rgb <= "000000";
					when "01100101001010111" => rgb <= "000000";
					when "01100101001011000" => rgb <= "000000";
					when "01100101001011001" => rgb <= "000000";
					when "01100101001011010" => rgb <= "000000";
					when "01100101001011011" => rgb <= "000000";
					when "01100101001011100" => rgb <= "000000";
					when "01100101001011101" => rgb <= "000000";
					when "01100101001011110" => rgb <= "000000";
					when "01100101001011111" => rgb <= "000000";
					when "01100101001100000" => rgb <= "000000";
					when "01100101001100001" => rgb <= "000000";
					when "01100101001100010" => rgb <= "000000";
					when "01100101001100011" => rgb <= "000000";
					when "01100101001100100" => rgb <= "000000";
					when "01100101001100101" => rgb <= "000000";
					when "01100101001100110" => rgb <= "000000";
					when "01100101001100111" => rgb <= "000000";
					when "01100101001101000" => rgb <= "000000";
					when "01100101001101001" => rgb <= "000000";
					when "01100101001101010" => rgb <= "000000";
					when "01100101001101011" => rgb <= "000000";
					when "01100101001101100" => rgb <= "000000";
					when "01100101001101101" => rgb <= "000000";
					when "01100101001101110" => rgb <= "000000";
					when "01100101001101111" => rgb <= "000000";
					when "01100101001110000" => rgb <= "000000";
					when "01100101001110001" => rgb <= "000000";
					when "01100101001110010" => rgb <= "000000";
					when "01100101001110011" => rgb <= "000000";
					when "01100101001110100" => rgb <= "000000";
					when "01100101001110101" => rgb <= "000000";
					when "01100101001110110" => rgb <= "000000";
					when "01100101001110111" => rgb <= "000000";
					when "01100101001111000" => rgb <= "000000";
					when "01100101001111001" => rgb <= "000000";
					when "01100101001111010" => rgb <= "000000";
					when "01100101001111011" => rgb <= "000000";
					when "01100101001111100" => rgb <= "000000";
					when "01100101001111101" => rgb <= "000000";
					when "01100101001111110" => rgb <= "000000";
					when "01100101001111111" => rgb <= "000000";
					when "01100101010000000" => rgb <= "000000";
					when "01100101010000001" => rgb <= "000000";
					when "01100101010000010" => rgb <= "000000";
					when "01100101010000011" => rgb <= "000000";
					when "01100101010000100" => rgb <= "000000";
					when "01100101010000101" => rgb <= "000000";
					when "01100101010000110" => rgb <= "000000";
					when "01100101010000111" => rgb <= "000000";
					when "01100101010001000" => rgb <= "000000";
					when "01100101010001001" => rgb <= "000000";
					when "01100101010001010" => rgb <= "000000";
					when "01100101010001011" => rgb <= "000000";
					when "01100101010001100" => rgb <= "000000";
					when "01100101010001101" => rgb <= "000000";
					when "01100101010001110" => rgb <= "000000";
					when "01100101010001111" => rgb <= "000000";
					when "01100101010010000" => rgb <= "000000";
					when "01100101010010001" => rgb <= "000000";
					when "01100101010010010" => rgb <= "000000";
					when "01100101010010011" => rgb <= "010000";
					when "01100101010010100" => rgb <= "101000";
					when "01100101010010101" => rgb <= "101000";
					when "01100101010010110" => rgb <= "101000";
					when "01100101010010111" => rgb <= "101000";
					when "01100101010011000" => rgb <= "101000";
					when "01100101010011001" => rgb <= "101000";
					when "01100101010011010" => rgb <= "101000";
					when "01100101010011011" => rgb <= "101000";
					when "01100101010011100" => rgb <= "101000";
					when "01100101010011101" => rgb <= "101000";
					when "01100101010011110" => rgb <= "101000";
					when "01100101010011111" => rgb <= "101000";
					when "01100101010100000" => rgb <= "101000";
					when "01100101010100001" => rgb <= "101000";
					when "01100101010100010" => rgb <= "101000";
					when "01100101010100011" => rgb <= "101000";
					when "01100101010100100" => rgb <= "101000";
					when "01100101010100101" => rgb <= "101000";
					when "01100101010100110" => rgb <= "101000";
					when "01100101010100111" => rgb <= "101000";
					when "01100101010101000" => rgb <= "101000";
					when "01100101010101001" => rgb <= "101000";
					when "01100101010101010" => rgb <= "010000";
					when "01100101010101011" => rgb <= "000000";
					when "01100101010101100" => rgb <= "000000";
					when "01100101010101101" => rgb <= "000000";
					when "01100101010101110" => rgb <= "000000";
					when "01100101010101111" => rgb <= "000000";
					when "01100101010110000" => rgb <= "000000";
					when "01100101010110001" => rgb <= "000000";
					when "01100101010110010" => rgb <= "000000";
					when "01100101010110011" => rgb <= "000000";
					when "01100101010110100" => rgb <= "000000";
					when "01100101010110101" => rgb <= "000000";
					when "01100101010110110" => rgb <= "000000";
					when "01100101010110111" => rgb <= "000000";
					when "01100101010111000" => rgb <= "000000";
					when "01100101010111001" => rgb <= "000000";
					when "01100101010111010" => rgb <= "000000";
					when "01100101010111011" => rgb <= "000000";
					when "01100101010111100" => rgb <= "000000";
					when "01100101010111101" => rgb <= "000000";
					when "01100101010111110" => rgb <= "000000";
					when "01100101010111111" => rgb <= "000000";
					when "01100101011000000" => rgb <= "000000";
					when "01100101011000001" => rgb <= "000000";
					when "01100101011000010" => rgb <= "000000";
					when "01100101011000011" => rgb <= "000000";
					when "01100101011000100" => rgb <= "000000";
					when "01100101011000101" => rgb <= "000000";
					when "01100101011000110" => rgb <= "000000";
					when "01100101011000111" => rgb <= "000000";
					when "01100101011001000" => rgb <= "000000";
					when "01100101011001001" => rgb <= "000000";
					when "01100101011001010" => rgb <= "000000";
					when "01100101011001011" => rgb <= "000000";
					when "01100101011001100" => rgb <= "000000";
					when "01100101011001101" => rgb <= "000000";
					when "01100101011001110" => rgb <= "000000";
					when "01100101011001111" => rgb <= "000000";
					when "01100101011010000" => rgb <= "000000";
					when "01100101011010001" => rgb <= "000000";
					when "01100101011010010" => rgb <= "000000";
					when "01100101011010011" => rgb <= "000000";
					when "01100101011010100" => rgb <= "000000";
					when "01100101011010101" => rgb <= "000000";
					when "01100101011010110" => rgb <= "000000";
					when "01100101011010111" => rgb <= "000000";
					when "01100101011011000" => rgb <= "000000";
					when "01100101011011001" => rgb <= "000000";
					when "01100101011011010" => rgb <= "000000";
					when "01100101011011011" => rgb <= "000000";
					when "01100101011011100" => rgb <= "000000";
					when "01100101011011101" => rgb <= "000000";
					when "01100101011011110" => rgb <= "000000";
					when "01100101011011111" => rgb <= "000000";
					when "01100101011100000" => rgb <= "000000";
					when "01100101011100001" => rgb <= "000000";
					when "01100101011100010" => rgb <= "000000";
					when "01100101011100011" => rgb <= "000000";
					when "01100101011100100" => rgb <= "000000";
					when "01100101011100101" => rgb <= "000000";
					when "01100101011100110" => rgb <= "000000";
					when "01100101011100111" => rgb <= "000000";
					when "01100101011101000" => rgb <= "000000";
					when "01100101011101001" => rgb <= "000000";
					when "01100101011101010" => rgb <= "000000";
					when "01100101011101011" => rgb <= "000000";
					when "01100101011101100" => rgb <= "000000";
					when "01100101011101101" => rgb <= "000000";
					when "01100101011101110" => rgb <= "000000";
					when "01100101011101111" => rgb <= "000000";
					when "01100101011110000" => rgb <= "000000";
					when "01100101011110001" => rgb <= "000000";
					when "01100101011110010" => rgb <= "000000";
					when "01100101011110011" => rgb <= "000000";
					when "01100101011110100" => rgb <= "000000";
					when "01100101011110101" => rgb <= "000000";
					when "01100101011110110" => rgb <= "000000";
					when "01100101011110111" => rgb <= "000000";
					when "01100101011111000" => rgb <= "000000";
					when "01100101011111001" => rgb <= "000000";
					when "01100101011111010" => rgb <= "000000";
					when "01100101011111011" => rgb <= "000000";
					when "01100101011111100" => rgb <= "000000";
					when "01100101011111101" => rgb <= "000000";
					when "01100101011111110" => rgb <= "000000";
					when "01100101011111111" => rgb <= "000000";
					when "01100101100000000" => rgb <= "000000";
					when "01100101100000001" => rgb <= "000000";
					when "01100101100000010" => rgb <= "000000";
					when "01100101100000011" => rgb <= "000000";
					when "01100101100000100" => rgb <= "000000";
					when "01100101100000101" => rgb <= "000000";
					when "01100101100000110" => rgb <= "000000";
					when "01100101100000111" => rgb <= "000000";
					when "01100101100001000" => rgb <= "000000";
					when "01100101100001001" => rgb <= "000000";
					when "01100101100001010" => rgb <= "000000";
					when "01100101100001011" => rgb <= "000000";
					when "01100101100001100" => rgb <= "000000";
					when "01100101100001101" => rgb <= "000000";
					when "01100101100001110" => rgb <= "000000";
					when "01100101100001111" => rgb <= "000000";
					when "01100101100010000" => rgb <= "000000";
					when "01100101100010001" => rgb <= "000000";
					when "01100101100010010" => rgb <= "000000";
					when "01100101100010011" => rgb <= "000000";
					when "01100101100010100" => rgb <= "000000";
					when "01100101100010101" => rgb <= "000000";
					when "01100101100010110" => rgb <= "000000";
					when "01100101100010111" => rgb <= "000000";
					when "01100101100011000" => rgb <= "000000";
					when "01100101100011001" => rgb <= "000000";
					when "01100101100011010" => rgb <= "000000";
					when "01100101100011011" => rgb <= "000000";
					when "01100101100011100" => rgb <= "000000";
					when "01100101100011101" => rgb <= "000000";
					when "01100101100011110" => rgb <= "000000";
					when "01100101100011111" => rgb <= "000000";
					when "01100101100100000" => rgb <= "000000";
					when "01100101100100001" => rgb <= "000000";
					when "01100101100100010" => rgb <= "000000";
					when "01100101100100011" => rgb <= "000000";
					when "01100101100100100" => rgb <= "000000";
					when "01100101100100101" => rgb <= "000000";
					when "01100101100100110" => rgb <= "000000";
					when "01100101100100111" => rgb <= "000000";
					when "01100101100101000" => rgb <= "000000";
					when "01100101100101001" => rgb <= "000000";
					when "01100101100101010" => rgb <= "000000";
					when "01100101100101011" => rgb <= "000000";
					when "01100101100101100" => rgb <= "000000";
					when "01100101100101101" => rgb <= "000000";
					when "01100101100101110" => rgb <= "000000";
					when "01100101100101111" => rgb <= "000000";
					when "01100101100110000" => rgb <= "000000";
					when "01100101100110001" => rgb <= "000000";
					when "01100101100110010" => rgb <= "000000";
					when "01100101100110011" => rgb <= "000000";
					when "01100101100110100" => rgb <= "000000";
					when "01100101100110101" => rgb <= "000000";
					when "01100101100110110" => rgb <= "000000";
					when "01100101100110111" => rgb <= "000000";
					when "01100101100111000" => rgb <= "000000";
					when "01100101100111001" => rgb <= "000000";
					when "01100101100111010" => rgb <= "000000";
					when "01100101100111011" => rgb <= "000000";
					when "01100101100111100" => rgb <= "000000";
					when "01100101100111101" => rgb <= "000000";
					when "01100101100111110" => rgb <= "000000";
					when "01100101100111111" => rgb <= "000000";
					when "01100110000000000" => rgb <= "000000";
					when "01100110000000001" => rgb <= "000000";
					when "01100110000000010" => rgb <= "000000";
					when "01100110000000011" => rgb <= "000000";
					when "01100110000000100" => rgb <= "000000";
					when "01100110000000101" => rgb <= "000000";
					when "01100110000000110" => rgb <= "000000";
					when "01100110000000111" => rgb <= "000000";
					when "01100110000001000" => rgb <= "000000";
					when "01100110000001001" => rgb <= "000000";
					when "01100110000001010" => rgb <= "000000";
					when "01100110000001011" => rgb <= "000000";
					when "01100110000001100" => rgb <= "000000";
					when "01100110000001101" => rgb <= "000000";
					when "01100110000001110" => rgb <= "000000";
					when "01100110000001111" => rgb <= "000000";
					when "01100110000010000" => rgb <= "000000";
					when "01100110000010001" => rgb <= "000000";
					when "01100110000010010" => rgb <= "000000";
					when "01100110000010011" => rgb <= "000000";
					when "01100110000010100" => rgb <= "000000";
					when "01100110000010101" => rgb <= "000000";
					when "01100110000010110" => rgb <= "000000";
					when "01100110000010111" => rgb <= "000000";
					when "01100110000011000" => rgb <= "000000";
					when "01100110000011001" => rgb <= "000000";
					when "01100110000011010" => rgb <= "000000";
					when "01100110000011011" => rgb <= "000000";
					when "01100110000011100" => rgb <= "000000";
					when "01100110000011101" => rgb <= "000000";
					when "01100110000011110" => rgb <= "000000";
					when "01100110000011111" => rgb <= "000000";
					when "01100110000100000" => rgb <= "000000";
					when "01100110000100001" => rgb <= "000000";
					when "01100110000100010" => rgb <= "000000";
					when "01100110000100011" => rgb <= "000000";
					when "01100110000100100" => rgb <= "000000";
					when "01100110000100101" => rgb <= "000000";
					when "01100110000100110" => rgb <= "000000";
					when "01100110000100111" => rgb <= "000000";
					when "01100110000101000" => rgb <= "000000";
					when "01100110000101001" => rgb <= "000000";
					when "01100110000101010" => rgb <= "000000";
					when "01100110000101011" => rgb <= "000000";
					when "01100110000101100" => rgb <= "000000";
					when "01100110000101101" => rgb <= "000000";
					when "01100110000101110" => rgb <= "000000";
					when "01100110000101111" => rgb <= "000000";
					when "01100110000110000" => rgb <= "000000";
					when "01100110000110001" => rgb <= "000000";
					when "01100110000110010" => rgb <= "000000";
					when "01100110000110011" => rgb <= "000000";
					when "01100110000110100" => rgb <= "000000";
					when "01100110000110101" => rgb <= "000000";
					when "01100110000110110" => rgb <= "000000";
					when "01100110000110111" => rgb <= "000000";
					when "01100110000111000" => rgb <= "000000";
					when "01100110000111001" => rgb <= "000000";
					when "01100110000111010" => rgb <= "000000";
					when "01100110000111011" => rgb <= "000000";
					when "01100110000111100" => rgb <= "000000";
					when "01100110000111101" => rgb <= "000000";
					when "01100110000111110" => rgb <= "000000";
					when "01100110000111111" => rgb <= "000000";
					when "01100110001000000" => rgb <= "000000";
					when "01100110001000001" => rgb <= "000000";
					when "01100110001000010" => rgb <= "000000";
					when "01100110001000011" => rgb <= "000000";
					when "01100110001000100" => rgb <= "000000";
					when "01100110001000101" => rgb <= "000000";
					when "01100110001000110" => rgb <= "000000";
					when "01100110001000111" => rgb <= "000000";
					when "01100110001001000" => rgb <= "000000";
					when "01100110001001001" => rgb <= "000000";
					when "01100110001001010" => rgb <= "000000";
					when "01100110001001011" => rgb <= "000000";
					when "01100110001001100" => rgb <= "000000";
					when "01100110001001101" => rgb <= "000000";
					when "01100110001001110" => rgb <= "000000";
					when "01100110001001111" => rgb <= "000000";
					when "01100110001010000" => rgb <= "000000";
					when "01100110001010001" => rgb <= "000000";
					when "01100110001010010" => rgb <= "000000";
					when "01100110001010011" => rgb <= "000000";
					when "01100110001010100" => rgb <= "000000";
					when "01100110001010101" => rgb <= "000000";
					when "01100110001010110" => rgb <= "000000";
					when "01100110001010111" => rgb <= "000000";
					when "01100110001011000" => rgb <= "000000";
					when "01100110001011001" => rgb <= "000000";
					when "01100110001011010" => rgb <= "000000";
					when "01100110001011011" => rgb <= "000000";
					when "01100110001011100" => rgb <= "000000";
					when "01100110001011101" => rgb <= "000000";
					when "01100110001011110" => rgb <= "000000";
					when "01100110001011111" => rgb <= "000000";
					when "01100110001100000" => rgb <= "000000";
					when "01100110001100001" => rgb <= "000000";
					when "01100110001100010" => rgb <= "000000";
					when "01100110001100011" => rgb <= "000000";
					when "01100110001100100" => rgb <= "000000";
					when "01100110001100101" => rgb <= "000000";
					when "01100110001100110" => rgb <= "000000";
					when "01100110001100111" => rgb <= "000000";
					when "01100110001101000" => rgb <= "000000";
					when "01100110001101001" => rgb <= "000000";
					when "01100110001101010" => rgb <= "000000";
					when "01100110001101011" => rgb <= "000000";
					when "01100110001101100" => rgb <= "000000";
					when "01100110001101101" => rgb <= "000000";
					when "01100110001101110" => rgb <= "000000";
					when "01100110001101111" => rgb <= "000000";
					when "01100110001110000" => rgb <= "000000";
					when "01100110001110001" => rgb <= "000000";
					when "01100110001110010" => rgb <= "000000";
					when "01100110001110011" => rgb <= "000000";
					when "01100110001110100" => rgb <= "000000";
					when "01100110001110101" => rgb <= "000000";
					when "01100110001110110" => rgb <= "000000";
					when "01100110001110111" => rgb <= "000000";
					when "01100110001111000" => rgb <= "000000";
					when "01100110001111001" => rgb <= "000000";
					when "01100110001111010" => rgb <= "000000";
					when "01100110001111011" => rgb <= "000000";
					when "01100110001111100" => rgb <= "000000";
					when "01100110001111101" => rgb <= "000000";
					when "01100110001111110" => rgb <= "000000";
					when "01100110001111111" => rgb <= "000000";
					when "01100110010000000" => rgb <= "000000";
					when "01100110010000001" => rgb <= "000000";
					when "01100110010000010" => rgb <= "000000";
					when "01100110010000011" => rgb <= "000000";
					when "01100110010000100" => rgb <= "000000";
					when "01100110010000101" => rgb <= "000000";
					when "01100110010000110" => rgb <= "000000";
					when "01100110010000111" => rgb <= "000000";
					when "01100110010001000" => rgb <= "000000";
					when "01100110010001001" => rgb <= "000000";
					when "01100110010001010" => rgb <= "000000";
					when "01100110010001011" => rgb <= "000000";
					when "01100110010001100" => rgb <= "000000";
					when "01100110010001101" => rgb <= "000000";
					when "01100110010001110" => rgb <= "000000";
					when "01100110010001111" => rgb <= "000000";
					when "01100110010010000" => rgb <= "000000";
					when "01100110010010001" => rgb <= "000000";
					when "01100110010010010" => rgb <= "000000";
					when "01100110010010011" => rgb <= "010000";
					when "01100110010010100" => rgb <= "101000";
					when "01100110010010101" => rgb <= "101000";
					when "01100110010010110" => rgb <= "101000";
					when "01100110010010111" => rgb <= "101000";
					when "01100110010011000" => rgb <= "101000";
					when "01100110010011001" => rgb <= "101000";
					when "01100110010011010" => rgb <= "101000";
					when "01100110010011011" => rgb <= "101000";
					when "01100110010011100" => rgb <= "101000";
					when "01100110010011101" => rgb <= "101000";
					when "01100110010011110" => rgb <= "101000";
					when "01100110010011111" => rgb <= "101000";
					when "01100110010100000" => rgb <= "101000";
					when "01100110010100001" => rgb <= "101000";
					when "01100110010100010" => rgb <= "101000";
					when "01100110010100011" => rgb <= "101000";
					when "01100110010100100" => rgb <= "101000";
					when "01100110010100101" => rgb <= "101000";
					when "01100110010100110" => rgb <= "101000";
					when "01100110010100111" => rgb <= "101000";
					when "01100110010101000" => rgb <= "101000";
					when "01100110010101001" => rgb <= "101000";
					when "01100110010101010" => rgb <= "010000";
					when "01100110010101011" => rgb <= "000000";
					when "01100110010101100" => rgb <= "000000";
					when "01100110010101101" => rgb <= "000000";
					when "01100110010101110" => rgb <= "000000";
					when "01100110010101111" => rgb <= "000000";
					when "01100110010110000" => rgb <= "000000";
					when "01100110010110001" => rgb <= "000000";
					when "01100110010110010" => rgb <= "000000";
					when "01100110010110011" => rgb <= "000000";
					when "01100110010110100" => rgb <= "000000";
					when "01100110010110101" => rgb <= "000000";
					when "01100110010110110" => rgb <= "000000";
					when "01100110010110111" => rgb <= "000000";
					when "01100110010111000" => rgb <= "000000";
					when "01100110010111001" => rgb <= "000000";
					when "01100110010111010" => rgb <= "000000";
					when "01100110010111011" => rgb <= "000000";
					when "01100110010111100" => rgb <= "000000";
					when "01100110010111101" => rgb <= "000000";
					when "01100110010111110" => rgb <= "000000";
					when "01100110010111111" => rgb <= "000000";
					when "01100110011000000" => rgb <= "000000";
					when "01100110011000001" => rgb <= "000000";
					when "01100110011000010" => rgb <= "000000";
					when "01100110011000011" => rgb <= "000000";
					when "01100110011000100" => rgb <= "000000";
					when "01100110011000101" => rgb <= "000000";
					when "01100110011000110" => rgb <= "000000";
					when "01100110011000111" => rgb <= "000000";
					when "01100110011001000" => rgb <= "000000";
					when "01100110011001001" => rgb <= "000000";
					when "01100110011001010" => rgb <= "000000";
					when "01100110011001011" => rgb <= "000000";
					when "01100110011001100" => rgb <= "000000";
					when "01100110011001101" => rgb <= "000000";
					when "01100110011001110" => rgb <= "000000";
					when "01100110011001111" => rgb <= "000000";
					when "01100110011010000" => rgb <= "000000";
					when "01100110011010001" => rgb <= "000000";
					when "01100110011010010" => rgb <= "000000";
					when "01100110011010011" => rgb <= "000000";
					when "01100110011010100" => rgb <= "000000";
					when "01100110011010101" => rgb <= "000000";
					when "01100110011010110" => rgb <= "000000";
					when "01100110011010111" => rgb <= "000000";
					when "01100110011011000" => rgb <= "000000";
					when "01100110011011001" => rgb <= "000000";
					when "01100110011011010" => rgb <= "000000";
					when "01100110011011011" => rgb <= "000000";
					when "01100110011011100" => rgb <= "000000";
					when "01100110011011101" => rgb <= "000000";
					when "01100110011011110" => rgb <= "000000";
					when "01100110011011111" => rgb <= "000000";
					when "01100110011100000" => rgb <= "000000";
					when "01100110011100001" => rgb <= "000000";
					when "01100110011100010" => rgb <= "000000";
					when "01100110011100011" => rgb <= "000000";
					when "01100110011100100" => rgb <= "000000";
					when "01100110011100101" => rgb <= "000000";
					when "01100110011100110" => rgb <= "000000";
					when "01100110011100111" => rgb <= "000000";
					when "01100110011101000" => rgb <= "000000";
					when "01100110011101001" => rgb <= "000000";
					when "01100110011101010" => rgb <= "000000";
					when "01100110011101011" => rgb <= "000000";
					when "01100110011101100" => rgb <= "000000";
					when "01100110011101101" => rgb <= "000000";
					when "01100110011101110" => rgb <= "000000";
					when "01100110011101111" => rgb <= "000000";
					when "01100110011110000" => rgb <= "000000";
					when "01100110011110001" => rgb <= "000000";
					when "01100110011110010" => rgb <= "000000";
					when "01100110011110011" => rgb <= "000000";
					when "01100110011110100" => rgb <= "000000";
					when "01100110011110101" => rgb <= "000000";
					when "01100110011110110" => rgb <= "000000";
					when "01100110011110111" => rgb <= "000000";
					when "01100110011111000" => rgb <= "000000";
					when "01100110011111001" => rgb <= "000000";
					when "01100110011111010" => rgb <= "000000";
					when "01100110011111011" => rgb <= "000000";
					when "01100110011111100" => rgb <= "000000";
					when "01100110011111101" => rgb <= "000000";
					when "01100110011111110" => rgb <= "000000";
					when "01100110011111111" => rgb <= "000000";
					when "01100110100000000" => rgb <= "000000";
					when "01100110100000001" => rgb <= "000000";
					when "01100110100000010" => rgb <= "000000";
					when "01100110100000011" => rgb <= "000000";
					when "01100110100000100" => rgb <= "000000";
					when "01100110100000101" => rgb <= "000000";
					when "01100110100000110" => rgb <= "000000";
					when "01100110100000111" => rgb <= "000000";
					when "01100110100001000" => rgb <= "000000";
					when "01100110100001001" => rgb <= "000000";
					when "01100110100001010" => rgb <= "000000";
					when "01100110100001011" => rgb <= "000000";
					when "01100110100001100" => rgb <= "000000";
					when "01100110100001101" => rgb <= "000000";
					when "01100110100001110" => rgb <= "000000";
					when "01100110100001111" => rgb <= "000000";
					when "01100110100010000" => rgb <= "000000";
					when "01100110100010001" => rgb <= "000000";
					when "01100110100010010" => rgb <= "000000";
					when "01100110100010011" => rgb <= "000000";
					when "01100110100010100" => rgb <= "000000";
					when "01100110100010101" => rgb <= "000000";
					when "01100110100010110" => rgb <= "000000";
					when "01100110100010111" => rgb <= "000000";
					when "01100110100011000" => rgb <= "000000";
					when "01100110100011001" => rgb <= "000000";
					when "01100110100011010" => rgb <= "000000";
					when "01100110100011011" => rgb <= "000000";
					when "01100110100011100" => rgb <= "000000";
					when "01100110100011101" => rgb <= "000000";
					when "01100110100011110" => rgb <= "000000";
					when "01100110100011111" => rgb <= "000000";
					when "01100110100100000" => rgb <= "000000";
					when "01100110100100001" => rgb <= "000000";
					when "01100110100100010" => rgb <= "000000";
					when "01100110100100011" => rgb <= "000000";
					when "01100110100100100" => rgb <= "000000";
					when "01100110100100101" => rgb <= "000000";
					when "01100110100100110" => rgb <= "000000";
					when "01100110100100111" => rgb <= "000000";
					when "01100110100101000" => rgb <= "000000";
					when "01100110100101001" => rgb <= "000000";
					when "01100110100101010" => rgb <= "000000";
					when "01100110100101011" => rgb <= "000000";
					when "01100110100101100" => rgb <= "000000";
					when "01100110100101101" => rgb <= "000000";
					when "01100110100101110" => rgb <= "000000";
					when "01100110100101111" => rgb <= "000000";
					when "01100110100110000" => rgb <= "000000";
					when "01100110100110001" => rgb <= "000000";
					when "01100110100110010" => rgb <= "000000";
					when "01100110100110011" => rgb <= "000000";
					when "01100110100110100" => rgb <= "000000";
					when "01100110100110101" => rgb <= "000000";
					when "01100110100110110" => rgb <= "000000";
					when "01100110100110111" => rgb <= "000000";
					when "01100110100111000" => rgb <= "000000";
					when "01100110100111001" => rgb <= "000000";
					when "01100110100111010" => rgb <= "000000";
					when "01100110100111011" => rgb <= "000000";
					when "01100110100111100" => rgb <= "000000";
					when "01100110100111101" => rgb <= "000000";
					when "01100110100111110" => rgb <= "000000";
					when "01100110100111111" => rgb <= "000000";
					when "01100111000000000" => rgb <= "000000";
					when "01100111000000001" => rgb <= "000000";
					when "01100111000000010" => rgb <= "000000";
					when "01100111000000011" => rgb <= "000000";
					when "01100111000000100" => rgb <= "000000";
					when "01100111000000101" => rgb <= "000000";
					when "01100111000000110" => rgb <= "000000";
					when "01100111000000111" => rgb <= "000000";
					when "01100111000001000" => rgb <= "000000";
					when "01100111000001001" => rgb <= "000000";
					when "01100111000001010" => rgb <= "000000";
					when "01100111000001011" => rgb <= "000000";
					when "01100111000001100" => rgb <= "000000";
					when "01100111000001101" => rgb <= "000000";
					when "01100111000001110" => rgb <= "000000";
					when "01100111000001111" => rgb <= "000000";
					when "01100111000010000" => rgb <= "000000";
					when "01100111000010001" => rgb <= "000000";
					when "01100111000010010" => rgb <= "000000";
					when "01100111000010011" => rgb <= "000000";
					when "01100111000010100" => rgb <= "000000";
					when "01100111000010101" => rgb <= "000000";
					when "01100111000010110" => rgb <= "000000";
					when "01100111000010111" => rgb <= "000000";
					when "01100111000011000" => rgb <= "000000";
					when "01100111000011001" => rgb <= "000000";
					when "01100111000011010" => rgb <= "000000";
					when "01100111000011011" => rgb <= "000000";
					when "01100111000011100" => rgb <= "000000";
					when "01100111000011101" => rgb <= "000000";
					when "01100111000011110" => rgb <= "000000";
					when "01100111000011111" => rgb <= "000000";
					when "01100111000100000" => rgb <= "000000";
					when "01100111000100001" => rgb <= "000000";
					when "01100111000100010" => rgb <= "000000";
					when "01100111000100011" => rgb <= "000000";
					when "01100111000100100" => rgb <= "000000";
					when "01100111000100101" => rgb <= "000000";
					when "01100111000100110" => rgb <= "000000";
					when "01100111000100111" => rgb <= "000000";
					when "01100111000101000" => rgb <= "000000";
					when "01100111000101001" => rgb <= "000000";
					when "01100111000101010" => rgb <= "000000";
					when "01100111000101011" => rgb <= "000000";
					when "01100111000101100" => rgb <= "000000";
					when "01100111000101101" => rgb <= "000000";
					when "01100111000101110" => rgb <= "000000";
					when "01100111000101111" => rgb <= "000000";
					when "01100111000110000" => rgb <= "000000";
					when "01100111000110001" => rgb <= "000000";
					when "01100111000110010" => rgb <= "000000";
					when "01100111000110011" => rgb <= "000000";
					when "01100111000110100" => rgb <= "000000";
					when "01100111000110101" => rgb <= "000000";
					when "01100111000110110" => rgb <= "000000";
					when "01100111000110111" => rgb <= "000000";
					when "01100111000111000" => rgb <= "000000";
					when "01100111000111001" => rgb <= "000000";
					when "01100111000111010" => rgb <= "000000";
					when "01100111000111011" => rgb <= "000000";
					when "01100111000111100" => rgb <= "000000";
					when "01100111000111101" => rgb <= "000000";
					when "01100111000111110" => rgb <= "000000";
					when "01100111000111111" => rgb <= "000000";
					when "01100111001000000" => rgb <= "000000";
					when "01100111001000001" => rgb <= "000000";
					when "01100111001000010" => rgb <= "000000";
					when "01100111001000011" => rgb <= "000000";
					when "01100111001000100" => rgb <= "000000";
					when "01100111001000101" => rgb <= "000000";
					when "01100111001000110" => rgb <= "000000";
					when "01100111001000111" => rgb <= "000000";
					when "01100111001001000" => rgb <= "000000";
					when "01100111001001001" => rgb <= "000000";
					when "01100111001001010" => rgb <= "000000";
					when "01100111001001011" => rgb <= "000000";
					when "01100111001001100" => rgb <= "000000";
					when "01100111001001101" => rgb <= "000000";
					when "01100111001001110" => rgb <= "000000";
					when "01100111001001111" => rgb <= "000000";
					when "01100111001010000" => rgb <= "000000";
					when "01100111001010001" => rgb <= "000000";
					when "01100111001010010" => rgb <= "000000";
					when "01100111001010011" => rgb <= "000000";
					when "01100111001010100" => rgb <= "000000";
					when "01100111001010101" => rgb <= "000000";
					when "01100111001010110" => rgb <= "000000";
					when "01100111001010111" => rgb <= "000000";
					when "01100111001011000" => rgb <= "000000";
					when "01100111001011001" => rgb <= "000000";
					when "01100111001011010" => rgb <= "000000";
					when "01100111001011011" => rgb <= "000000";
					when "01100111001011100" => rgb <= "000000";
					when "01100111001011101" => rgb <= "000000";
					when "01100111001011110" => rgb <= "000000";
					when "01100111001011111" => rgb <= "000000";
					when "01100111001100000" => rgb <= "000000";
					when "01100111001100001" => rgb <= "000000";
					when "01100111001100010" => rgb <= "000000";
					when "01100111001100011" => rgb <= "000000";
					when "01100111001100100" => rgb <= "000000";
					when "01100111001100101" => rgb <= "000000";
					when "01100111001100110" => rgb <= "000000";
					when "01100111001100111" => rgb <= "000000";
					when "01100111001101000" => rgb <= "000000";
					when "01100111001101001" => rgb <= "000000";
					when "01100111001101010" => rgb <= "000000";
					when "01100111001101011" => rgb <= "000000";
					when "01100111001101100" => rgb <= "000000";
					when "01100111001101101" => rgb <= "000000";
					when "01100111001101110" => rgb <= "000000";
					when "01100111001101111" => rgb <= "000000";
					when "01100111001110000" => rgb <= "000000";
					when "01100111001110001" => rgb <= "000000";
					when "01100111001110010" => rgb <= "000000";
					when "01100111001110011" => rgb <= "000000";
					when "01100111001110100" => rgb <= "000000";
					when "01100111001110101" => rgb <= "000000";
					when "01100111001110110" => rgb <= "000000";
					when "01100111001110111" => rgb <= "000000";
					when "01100111001111000" => rgb <= "000000";
					when "01100111001111001" => rgb <= "000000";
					when "01100111001111010" => rgb <= "000000";
					when "01100111001111011" => rgb <= "000000";
					when "01100111001111100" => rgb <= "000000";
					when "01100111001111101" => rgb <= "000000";
					when "01100111001111110" => rgb <= "000000";
					when "01100111001111111" => rgb <= "000000";
					when "01100111010000000" => rgb <= "000000";
					when "01100111010000001" => rgb <= "000000";
					when "01100111010000010" => rgb <= "000000";
					when "01100111010000011" => rgb <= "000000";
					when "01100111010000100" => rgb <= "000000";
					when "01100111010000101" => rgb <= "000000";
					when "01100111010000110" => rgb <= "000000";
					when "01100111010000111" => rgb <= "000000";
					when "01100111010001000" => rgb <= "000000";
					when "01100111010001001" => rgb <= "000000";
					when "01100111010001010" => rgb <= "000000";
					when "01100111010001011" => rgb <= "000000";
					when "01100111010001100" => rgb <= "000000";
					when "01100111010001101" => rgb <= "000000";
					when "01100111010001110" => rgb <= "000000";
					when "01100111010001111" => rgb <= "000000";
					when "01100111010010000" => rgb <= "000000";
					when "01100111010010001" => rgb <= "000000";
					when "01100111010010010" => rgb <= "000000";
					when "01100111010010011" => rgb <= "010000";
					when "01100111010010100" => rgb <= "101000";
					when "01100111010010101" => rgb <= "101000";
					when "01100111010010110" => rgb <= "101000";
					when "01100111010010111" => rgb <= "101000";
					when "01100111010011000" => rgb <= "101000";
					when "01100111010011001" => rgb <= "101000";
					when "01100111010011010" => rgb <= "101000";
					when "01100111010011011" => rgb <= "101000";
					when "01100111010011100" => rgb <= "101000";
					when "01100111010011101" => rgb <= "101000";
					when "01100111010011110" => rgb <= "101000";
					when "01100111010011111" => rgb <= "101000";
					when "01100111010100000" => rgb <= "101000";
					when "01100111010100001" => rgb <= "101000";
					when "01100111010100010" => rgb <= "101000";
					when "01100111010100011" => rgb <= "101000";
					when "01100111010100100" => rgb <= "101000";
					when "01100111010100101" => rgb <= "101000";
					when "01100111010100110" => rgb <= "101000";
					when "01100111010100111" => rgb <= "101000";
					when "01100111010101000" => rgb <= "101000";
					when "01100111010101001" => rgb <= "101000";
					when "01100111010101010" => rgb <= "010000";
					when "01100111010101011" => rgb <= "000000";
					when "01100111010101100" => rgb <= "000000";
					when "01100111010101101" => rgb <= "000000";
					when "01100111010101110" => rgb <= "000000";
					when "01100111010101111" => rgb <= "000000";
					when "01100111010110000" => rgb <= "000000";
					when "01100111010110001" => rgb <= "000000";
					when "01100111010110010" => rgb <= "000000";
					when "01100111010110011" => rgb <= "000000";
					when "01100111010110100" => rgb <= "000000";
					when "01100111010110101" => rgb <= "000000";
					when "01100111010110110" => rgb <= "000000";
					when "01100111010110111" => rgb <= "000000";
					when "01100111010111000" => rgb <= "000000";
					when "01100111010111001" => rgb <= "000000";
					when "01100111010111010" => rgb <= "000000";
					when "01100111010111011" => rgb <= "000000";
					when "01100111010111100" => rgb <= "000000";
					when "01100111010111101" => rgb <= "000000";
					when "01100111010111110" => rgb <= "000000";
					when "01100111010111111" => rgb <= "000000";
					when "01100111011000000" => rgb <= "000000";
					when "01100111011000001" => rgb <= "000000";
					when "01100111011000010" => rgb <= "000000";
					when "01100111011000011" => rgb <= "000000";
					when "01100111011000100" => rgb <= "000000";
					when "01100111011000101" => rgb <= "000000";
					when "01100111011000110" => rgb <= "000000";
					when "01100111011000111" => rgb <= "000000";
					when "01100111011001000" => rgb <= "000000";
					when "01100111011001001" => rgb <= "000000";
					when "01100111011001010" => rgb <= "000000";
					when "01100111011001011" => rgb <= "000000";
					when "01100111011001100" => rgb <= "000000";
					when "01100111011001101" => rgb <= "000000";
					when "01100111011001110" => rgb <= "000000";
					when "01100111011001111" => rgb <= "000000";
					when "01100111011010000" => rgb <= "000000";
					when "01100111011010001" => rgb <= "000000";
					when "01100111011010010" => rgb <= "000000";
					when "01100111011010011" => rgb <= "000000";
					when "01100111011010100" => rgb <= "000000";
					when "01100111011010101" => rgb <= "000000";
					when "01100111011010110" => rgb <= "000000";
					when "01100111011010111" => rgb <= "000000";
					when "01100111011011000" => rgb <= "000000";
					when "01100111011011001" => rgb <= "000000";
					when "01100111011011010" => rgb <= "000000";
					when "01100111011011011" => rgb <= "000000";
					when "01100111011011100" => rgb <= "000000";
					when "01100111011011101" => rgb <= "000000";
					when "01100111011011110" => rgb <= "000000";
					when "01100111011011111" => rgb <= "000000";
					when "01100111011100000" => rgb <= "000000";
					when "01100111011100001" => rgb <= "000000";
					when "01100111011100010" => rgb <= "000000";
					when "01100111011100011" => rgb <= "000000";
					when "01100111011100100" => rgb <= "000000";
					when "01100111011100101" => rgb <= "000000";
					when "01100111011100110" => rgb <= "000000";
					when "01100111011100111" => rgb <= "000000";
					when "01100111011101000" => rgb <= "000000";
					when "01100111011101001" => rgb <= "000000";
					when "01100111011101010" => rgb <= "000000";
					when "01100111011101011" => rgb <= "000000";
					when "01100111011101100" => rgb <= "000000";
					when "01100111011101101" => rgb <= "000000";
					when "01100111011101110" => rgb <= "000000";
					when "01100111011101111" => rgb <= "000000";
					when "01100111011110000" => rgb <= "000000";
					when "01100111011110001" => rgb <= "000000";
					when "01100111011110010" => rgb <= "000000";
					when "01100111011110011" => rgb <= "000000";
					when "01100111011110100" => rgb <= "000000";
					when "01100111011110101" => rgb <= "000000";
					when "01100111011110110" => rgb <= "000000";
					when "01100111011110111" => rgb <= "000000";
					when "01100111011111000" => rgb <= "000000";
					when "01100111011111001" => rgb <= "000000";
					when "01100111011111010" => rgb <= "000000";
					when "01100111011111011" => rgb <= "000000";
					when "01100111011111100" => rgb <= "000000";
					when "01100111011111101" => rgb <= "000000";
					when "01100111011111110" => rgb <= "000000";
					when "01100111011111111" => rgb <= "000000";
					when "01100111100000000" => rgb <= "000000";
					when "01100111100000001" => rgb <= "000000";
					when "01100111100000010" => rgb <= "000000";
					when "01100111100000011" => rgb <= "000000";
					when "01100111100000100" => rgb <= "000000";
					when "01100111100000101" => rgb <= "000000";
					when "01100111100000110" => rgb <= "000000";
					when "01100111100000111" => rgb <= "000000";
					when "01100111100001000" => rgb <= "000000";
					when "01100111100001001" => rgb <= "000000";
					when "01100111100001010" => rgb <= "000000";
					when "01100111100001011" => rgb <= "000000";
					when "01100111100001100" => rgb <= "000000";
					when "01100111100001101" => rgb <= "000000";
					when "01100111100001110" => rgb <= "000000";
					when "01100111100001111" => rgb <= "000000";
					when "01100111100010000" => rgb <= "000000";
					when "01100111100010001" => rgb <= "000000";
					when "01100111100010010" => rgb <= "000000";
					when "01100111100010011" => rgb <= "000000";
					when "01100111100010100" => rgb <= "000000";
					when "01100111100010101" => rgb <= "000000";
					when "01100111100010110" => rgb <= "000000";
					when "01100111100010111" => rgb <= "000000";
					when "01100111100011000" => rgb <= "000000";
					when "01100111100011001" => rgb <= "000000";
					when "01100111100011010" => rgb <= "000000";
					when "01100111100011011" => rgb <= "000000";
					when "01100111100011100" => rgb <= "000000";
					when "01100111100011101" => rgb <= "000000";
					when "01100111100011110" => rgb <= "000000";
					when "01100111100011111" => rgb <= "000000";
					when "01100111100100000" => rgb <= "000000";
					when "01100111100100001" => rgb <= "000000";
					when "01100111100100010" => rgb <= "000000";
					when "01100111100100011" => rgb <= "000000";
					when "01100111100100100" => rgb <= "000000";
					when "01100111100100101" => rgb <= "000000";
					when "01100111100100110" => rgb <= "000000";
					when "01100111100100111" => rgb <= "000000";
					when "01100111100101000" => rgb <= "000000";
					when "01100111100101001" => rgb <= "000000";
					when "01100111100101010" => rgb <= "000000";
					when "01100111100101011" => rgb <= "000000";
					when "01100111100101100" => rgb <= "000000";
					when "01100111100101101" => rgb <= "000000";
					when "01100111100101110" => rgb <= "000000";
					when "01100111100101111" => rgb <= "000000";
					when "01100111100110000" => rgb <= "000000";
					when "01100111100110001" => rgb <= "000000";
					when "01100111100110010" => rgb <= "000000";
					when "01100111100110011" => rgb <= "000000";
					when "01100111100110100" => rgb <= "000000";
					when "01100111100110101" => rgb <= "000000";
					when "01100111100110110" => rgb <= "000000";
					when "01100111100110111" => rgb <= "000000";
					when "01100111100111000" => rgb <= "000000";
					when "01100111100111001" => rgb <= "000000";
					when "01100111100111010" => rgb <= "000000";
					when "01100111100111011" => rgb <= "000000";
					when "01100111100111100" => rgb <= "000000";
					when "01100111100111101" => rgb <= "000000";
					when "01100111100111110" => rgb <= "000000";
					when "01100111100111111" => rgb <= "000000";
					when "01101000000000000" => rgb <= "000000";
					when "01101000000000001" => rgb <= "000000";
					when "01101000000000010" => rgb <= "000000";
					when "01101000000000011" => rgb <= "000000";
					when "01101000000000100" => rgb <= "000000";
					when "01101000000000101" => rgb <= "000000";
					when "01101000000000110" => rgb <= "000000";
					when "01101000000000111" => rgb <= "000000";
					when "01101000000001000" => rgb <= "000000";
					when "01101000000001001" => rgb <= "000000";
					when "01101000000001010" => rgb <= "000000";
					when "01101000000001011" => rgb <= "000000";
					when "01101000000001100" => rgb <= "000000";
					when "01101000000001101" => rgb <= "000000";
					when "01101000000001110" => rgb <= "000000";
					when "01101000000001111" => rgb <= "000000";
					when "01101000000010000" => rgb <= "000000";
					when "01101000000010001" => rgb <= "000000";
					when "01101000000010010" => rgb <= "000000";
					when "01101000000010011" => rgb <= "000000";
					when "01101000000010100" => rgb <= "000000";
					when "01101000000010101" => rgb <= "000000";
					when "01101000000010110" => rgb <= "000000";
					when "01101000000010111" => rgb <= "000000";
					when "01101000000011000" => rgb <= "000000";
					when "01101000000011001" => rgb <= "000000";
					when "01101000000011010" => rgb <= "000000";
					when "01101000000011011" => rgb <= "000000";
					when "01101000000011100" => rgb <= "000000";
					when "01101000000011101" => rgb <= "000000";
					when "01101000000011110" => rgb <= "000000";
					when "01101000000011111" => rgb <= "000000";
					when "01101000000100000" => rgb <= "000000";
					when "01101000000100001" => rgb <= "000000";
					when "01101000000100010" => rgb <= "000000";
					when "01101000000100011" => rgb <= "000000";
					when "01101000000100100" => rgb <= "000000";
					when "01101000000100101" => rgb <= "000000";
					when "01101000000100110" => rgb <= "000000";
					when "01101000000100111" => rgb <= "000000";
					when "01101000000101000" => rgb <= "000000";
					when "01101000000101001" => rgb <= "000000";
					when "01101000000101010" => rgb <= "000000";
					when "01101000000101011" => rgb <= "000000";
					when "01101000000101100" => rgb <= "000000";
					when "01101000000101101" => rgb <= "000000";
					when "01101000000101110" => rgb <= "000000";
					when "01101000000101111" => rgb <= "000000";
					when "01101000000110000" => rgb <= "000000";
					when "01101000000110001" => rgb <= "000000";
					when "01101000000110010" => rgb <= "000000";
					when "01101000000110011" => rgb <= "000000";
					when "01101000000110100" => rgb <= "000000";
					when "01101000000110101" => rgb <= "000000";
					when "01101000000110110" => rgb <= "000000";
					when "01101000000110111" => rgb <= "000000";
					when "01101000000111000" => rgb <= "000000";
					when "01101000000111001" => rgb <= "000000";
					when "01101000000111010" => rgb <= "000000";
					when "01101000000111011" => rgb <= "000000";
					when "01101000000111100" => rgb <= "000000";
					when "01101000000111101" => rgb <= "000000";
					when "01101000000111110" => rgb <= "000000";
					when "01101000000111111" => rgb <= "000000";
					when "01101000001000000" => rgb <= "000000";
					when "01101000001000001" => rgb <= "000000";
					when "01101000001000010" => rgb <= "000000";
					when "01101000001000011" => rgb <= "000000";
					when "01101000001000100" => rgb <= "000000";
					when "01101000001000101" => rgb <= "000000";
					when "01101000001000110" => rgb <= "000000";
					when "01101000001000111" => rgb <= "000000";
					when "01101000001001000" => rgb <= "000000";
					when "01101000001001001" => rgb <= "000000";
					when "01101000001001010" => rgb <= "000000";
					when "01101000001001011" => rgb <= "000000";
					when "01101000001001100" => rgb <= "000000";
					when "01101000001001101" => rgb <= "000000";
					when "01101000001001110" => rgb <= "000000";
					when "01101000001001111" => rgb <= "000000";
					when "01101000001010000" => rgb <= "000000";
					when "01101000001010001" => rgb <= "000000";
					when "01101000001010010" => rgb <= "000000";
					when "01101000001010011" => rgb <= "000000";
					when "01101000001010100" => rgb <= "000000";
					when "01101000001010101" => rgb <= "000000";
					when "01101000001010110" => rgb <= "000000";
					when "01101000001010111" => rgb <= "000000";
					when "01101000001011000" => rgb <= "000000";
					when "01101000001011001" => rgb <= "000000";
					when "01101000001011010" => rgb <= "000000";
					when "01101000001011011" => rgb <= "000000";
					when "01101000001011100" => rgb <= "000000";
					when "01101000001011101" => rgb <= "000000";
					when "01101000001011110" => rgb <= "000000";
					when "01101000001011111" => rgb <= "000000";
					when "01101000001100000" => rgb <= "000000";
					when "01101000001100001" => rgb <= "000000";
					when "01101000001100010" => rgb <= "000000";
					when "01101000001100011" => rgb <= "000000";
					when "01101000001100100" => rgb <= "000000";
					when "01101000001100101" => rgb <= "000000";
					when "01101000001100110" => rgb <= "000000";
					when "01101000001100111" => rgb <= "000000";
					when "01101000001101000" => rgb <= "000000";
					when "01101000001101001" => rgb <= "000000";
					when "01101000001101010" => rgb <= "000000";
					when "01101000001101011" => rgb <= "000000";
					when "01101000001101100" => rgb <= "000000";
					when "01101000001101101" => rgb <= "000000";
					when "01101000001101110" => rgb <= "000000";
					when "01101000001101111" => rgb <= "000000";
					when "01101000001110000" => rgb <= "000000";
					when "01101000001110001" => rgb <= "000000";
					when "01101000001110010" => rgb <= "000000";
					when "01101000001110011" => rgb <= "000000";
					when "01101000001110100" => rgb <= "000000";
					when "01101000001110101" => rgb <= "000000";
					when "01101000001110110" => rgb <= "000000";
					when "01101000001110111" => rgb <= "000000";
					when "01101000001111000" => rgb <= "000000";
					when "01101000001111001" => rgb <= "000000";
					when "01101000001111010" => rgb <= "000000";
					when "01101000001111011" => rgb <= "000000";
					when "01101000001111100" => rgb <= "000000";
					when "01101000001111101" => rgb <= "000000";
					when "01101000001111110" => rgb <= "000000";
					when "01101000001111111" => rgb <= "000000";
					when "01101000010000000" => rgb <= "000000";
					when "01101000010000001" => rgb <= "000000";
					when "01101000010000010" => rgb <= "000000";
					when "01101000010000011" => rgb <= "000000";
					when "01101000010000100" => rgb <= "000000";
					when "01101000010000101" => rgb <= "000000";
					when "01101000010000110" => rgb <= "000000";
					when "01101000010000111" => rgb <= "000000";
					when "01101000010001000" => rgb <= "000000";
					when "01101000010001001" => rgb <= "000000";
					when "01101000010001010" => rgb <= "000000";
					when "01101000010001011" => rgb <= "000000";
					when "01101000010001100" => rgb <= "000000";
					when "01101000010001101" => rgb <= "000000";
					when "01101000010001110" => rgb <= "000000";
					when "01101000010001111" => rgb <= "000000";
					when "01101000010010000" => rgb <= "000000";
					when "01101000010010001" => rgb <= "000000";
					when "01101000010010010" => rgb <= "000000";
					when "01101000010010011" => rgb <= "010000";
					when "01101000010010100" => rgb <= "101000";
					when "01101000010010101" => rgb <= "101000";
					when "01101000010010110" => rgb <= "101000";
					when "01101000010010111" => rgb <= "101000";
					when "01101000010011000" => rgb <= "101000";
					when "01101000010011001" => rgb <= "101000";
					when "01101000010011010" => rgb <= "101000";
					when "01101000010011011" => rgb <= "101000";
					when "01101000010011100" => rgb <= "101000";
					when "01101000010011101" => rgb <= "101000";
					when "01101000010011110" => rgb <= "101000";
					when "01101000010011111" => rgb <= "101000";
					when "01101000010100000" => rgb <= "101000";
					when "01101000010100001" => rgb <= "101000";
					when "01101000010100010" => rgb <= "101000";
					when "01101000010100011" => rgb <= "101000";
					when "01101000010100100" => rgb <= "101000";
					when "01101000010100101" => rgb <= "101000";
					when "01101000010100110" => rgb <= "101000";
					when "01101000010100111" => rgb <= "101000";
					when "01101000010101000" => rgb <= "101000";
					when "01101000010101001" => rgb <= "101000";
					when "01101000010101010" => rgb <= "010000";
					when "01101000010101011" => rgb <= "000000";
					when "01101000010101100" => rgb <= "000000";
					when "01101000010101101" => rgb <= "000000";
					when "01101000010101110" => rgb <= "000000";
					when "01101000010101111" => rgb <= "000000";
					when "01101000010110000" => rgb <= "000000";
					when "01101000010110001" => rgb <= "000000";
					when "01101000010110010" => rgb <= "000000";
					when "01101000010110011" => rgb <= "000000";
					when "01101000010110100" => rgb <= "000000";
					when "01101000010110101" => rgb <= "000000";
					when "01101000010110110" => rgb <= "000000";
					when "01101000010110111" => rgb <= "000000";
					when "01101000010111000" => rgb <= "000000";
					when "01101000010111001" => rgb <= "000000";
					when "01101000010111010" => rgb <= "000000";
					when "01101000010111011" => rgb <= "000000";
					when "01101000010111100" => rgb <= "000000";
					when "01101000010111101" => rgb <= "000000";
					when "01101000010111110" => rgb <= "000000";
					when "01101000010111111" => rgb <= "000000";
					when "01101000011000000" => rgb <= "000000";
					when "01101000011000001" => rgb <= "000000";
					when "01101000011000010" => rgb <= "000000";
					when "01101000011000011" => rgb <= "000000";
					when "01101000011000100" => rgb <= "000000";
					when "01101000011000101" => rgb <= "000000";
					when "01101000011000110" => rgb <= "000000";
					when "01101000011000111" => rgb <= "000000";
					when "01101000011001000" => rgb <= "000000";
					when "01101000011001001" => rgb <= "000000";
					when "01101000011001010" => rgb <= "000000";
					when "01101000011001011" => rgb <= "000000";
					when "01101000011001100" => rgb <= "000000";
					when "01101000011001101" => rgb <= "000000";
					when "01101000011001110" => rgb <= "000000";
					when "01101000011001111" => rgb <= "000000";
					when "01101000011010000" => rgb <= "000000";
					when "01101000011010001" => rgb <= "000000";
					when "01101000011010010" => rgb <= "000000";
					when "01101000011010011" => rgb <= "000000";
					when "01101000011010100" => rgb <= "000000";
					when "01101000011010101" => rgb <= "000000";
					when "01101000011010110" => rgb <= "000000";
					when "01101000011010111" => rgb <= "000000";
					when "01101000011011000" => rgb <= "000000";
					when "01101000011011001" => rgb <= "000000";
					when "01101000011011010" => rgb <= "000000";
					when "01101000011011011" => rgb <= "000000";
					when "01101000011011100" => rgb <= "000000";
					when "01101000011011101" => rgb <= "000000";
					when "01101000011011110" => rgb <= "000000";
					when "01101000011011111" => rgb <= "000000";
					when "01101000011100000" => rgb <= "000000";
					when "01101000011100001" => rgb <= "000000";
					when "01101000011100010" => rgb <= "000000";
					when "01101000011100011" => rgb <= "000000";
					when "01101000011100100" => rgb <= "000000";
					when "01101000011100101" => rgb <= "000000";
					when "01101000011100110" => rgb <= "000000";
					when "01101000011100111" => rgb <= "000000";
					when "01101000011101000" => rgb <= "000000";
					when "01101000011101001" => rgb <= "000000";
					when "01101000011101010" => rgb <= "000000";
					when "01101000011101011" => rgb <= "000000";
					when "01101000011101100" => rgb <= "000000";
					when "01101000011101101" => rgb <= "000000";
					when "01101000011101110" => rgb <= "000000";
					when "01101000011101111" => rgb <= "000000";
					when "01101000011110000" => rgb <= "000000";
					when "01101000011110001" => rgb <= "000000";
					when "01101000011110010" => rgb <= "000000";
					when "01101000011110011" => rgb <= "000000";
					when "01101000011110100" => rgb <= "000000";
					when "01101000011110101" => rgb <= "000000";
					when "01101000011110110" => rgb <= "000000";
					when "01101000011110111" => rgb <= "000000";
					when "01101000011111000" => rgb <= "000000";
					when "01101000011111001" => rgb <= "000000";
					when "01101000011111010" => rgb <= "000000";
					when "01101000011111011" => rgb <= "000000";
					when "01101000011111100" => rgb <= "000000";
					when "01101000011111101" => rgb <= "000000";
					when "01101000011111110" => rgb <= "000000";
					when "01101000011111111" => rgb <= "000000";
					when "01101000100000000" => rgb <= "000000";
					when "01101000100000001" => rgb <= "000000";
					when "01101000100000010" => rgb <= "000000";
					when "01101000100000011" => rgb <= "000000";
					when "01101000100000100" => rgb <= "000000";
					when "01101000100000101" => rgb <= "000000";
					when "01101000100000110" => rgb <= "000000";
					when "01101000100000111" => rgb <= "000000";
					when "01101000100001000" => rgb <= "000000";
					when "01101000100001001" => rgb <= "000000";
					when "01101000100001010" => rgb <= "000000";
					when "01101000100001011" => rgb <= "000000";
					when "01101000100001100" => rgb <= "000000";
					when "01101000100001101" => rgb <= "000000";
					when "01101000100001110" => rgb <= "000000";
					when "01101000100001111" => rgb <= "000000";
					when "01101000100010000" => rgb <= "000000";
					when "01101000100010001" => rgb <= "000000";
					when "01101000100010010" => rgb <= "000000";
					when "01101000100010011" => rgb <= "000000";
					when "01101000100010100" => rgb <= "000000";
					when "01101000100010101" => rgb <= "000000";
					when "01101000100010110" => rgb <= "000000";
					when "01101000100010111" => rgb <= "000000";
					when "01101000100011000" => rgb <= "000000";
					when "01101000100011001" => rgb <= "000000";
					when "01101000100011010" => rgb <= "000000";
					when "01101000100011011" => rgb <= "000000";
					when "01101000100011100" => rgb <= "000000";
					when "01101000100011101" => rgb <= "000000";
					when "01101000100011110" => rgb <= "000000";
					when "01101000100011111" => rgb <= "000000";
					when "01101000100100000" => rgb <= "000000";
					when "01101000100100001" => rgb <= "000000";
					when "01101000100100010" => rgb <= "000000";
					when "01101000100100011" => rgb <= "000000";
					when "01101000100100100" => rgb <= "000000";
					when "01101000100100101" => rgb <= "000000";
					when "01101000100100110" => rgb <= "000000";
					when "01101000100100111" => rgb <= "000000";
					when "01101000100101000" => rgb <= "000000";
					when "01101000100101001" => rgb <= "000000";
					when "01101000100101010" => rgb <= "000000";
					when "01101000100101011" => rgb <= "000000";
					when "01101000100101100" => rgb <= "000000";
					when "01101000100101101" => rgb <= "000000";
					when "01101000100101110" => rgb <= "000000";
					when "01101000100101111" => rgb <= "000000";
					when "01101000100110000" => rgb <= "000000";
					when "01101000100110001" => rgb <= "000000";
					when "01101000100110010" => rgb <= "000000";
					when "01101000100110011" => rgb <= "000000";
					when "01101000100110100" => rgb <= "000000";
					when "01101000100110101" => rgb <= "000000";
					when "01101000100110110" => rgb <= "000000";
					when "01101000100110111" => rgb <= "000000";
					when "01101000100111000" => rgb <= "000000";
					when "01101000100111001" => rgb <= "000000";
					when "01101000100111010" => rgb <= "000000";
					when "01101000100111011" => rgb <= "000000";
					when "01101000100111100" => rgb <= "000000";
					when "01101000100111101" => rgb <= "000000";
					when "01101000100111110" => rgb <= "000000";
					when "01101000100111111" => rgb <= "000000";
					when "01101001000000000" => rgb <= "000000";
					when "01101001000000001" => rgb <= "000000";
					when "01101001000000010" => rgb <= "000000";
					when "01101001000000011" => rgb <= "000000";
					when "01101001000000100" => rgb <= "000000";
					when "01101001000000101" => rgb <= "000000";
					when "01101001000000110" => rgb <= "000000";
					when "01101001000000111" => rgb <= "000000";
					when "01101001000001000" => rgb <= "000000";
					when "01101001000001001" => rgb <= "000000";
					when "01101001000001010" => rgb <= "000000";
					when "01101001000001011" => rgb <= "000000";
					when "01101001000001100" => rgb <= "000000";
					when "01101001000001101" => rgb <= "000000";
					when "01101001000001110" => rgb <= "000000";
					when "01101001000001111" => rgb <= "000000";
					when "01101001000010000" => rgb <= "000000";
					when "01101001000010001" => rgb <= "000000";
					when "01101001000010010" => rgb <= "000000";
					when "01101001000010011" => rgb <= "000000";
					when "01101001000010100" => rgb <= "000000";
					when "01101001000010101" => rgb <= "000000";
					when "01101001000010110" => rgb <= "000000";
					when "01101001000010111" => rgb <= "000000";
					when "01101001000011000" => rgb <= "000000";
					when "01101001000011001" => rgb <= "000000";
					when "01101001000011010" => rgb <= "000000";
					when "01101001000011011" => rgb <= "000000";
					when "01101001000011100" => rgb <= "000000";
					when "01101001000011101" => rgb <= "000000";
					when "01101001000011110" => rgb <= "000000";
					when "01101001000011111" => rgb <= "000000";
					when "01101001000100000" => rgb <= "000000";
					when "01101001000100001" => rgb <= "000000";
					when "01101001000100010" => rgb <= "000000";
					when "01101001000100011" => rgb <= "000000";
					when "01101001000100100" => rgb <= "000000";
					when "01101001000100101" => rgb <= "000000";
					when "01101001000100110" => rgb <= "000000";
					when "01101001000100111" => rgb <= "000000";
					when "01101001000101000" => rgb <= "000000";
					when "01101001000101001" => rgb <= "000000";
					when "01101001000101010" => rgb <= "000000";
					when "01101001000101011" => rgb <= "000000";
					when "01101001000101100" => rgb <= "000000";
					when "01101001000101101" => rgb <= "000000";
					when "01101001000101110" => rgb <= "000000";
					when "01101001000101111" => rgb <= "000000";
					when "01101001000110000" => rgb <= "000000";
					when "01101001000110001" => rgb <= "000000";
					when "01101001000110010" => rgb <= "000000";
					when "01101001000110011" => rgb <= "000000";
					when "01101001000110100" => rgb <= "000000";
					when "01101001000110101" => rgb <= "000000";
					when "01101001000110110" => rgb <= "000000";
					when "01101001000110111" => rgb <= "000000";
					when "01101001000111000" => rgb <= "000000";
					when "01101001000111001" => rgb <= "000000";
					when "01101001000111010" => rgb <= "000000";
					when "01101001000111011" => rgb <= "000000";
					when "01101001000111100" => rgb <= "000000";
					when "01101001000111101" => rgb <= "000000";
					when "01101001000111110" => rgb <= "000000";
					when "01101001000111111" => rgb <= "000000";
					when "01101001001000000" => rgb <= "000000";
					when "01101001001000001" => rgb <= "000000";
					when "01101001001000010" => rgb <= "000000";
					when "01101001001000011" => rgb <= "000000";
					when "01101001001000100" => rgb <= "000000";
					when "01101001001000101" => rgb <= "000000";
					when "01101001001000110" => rgb <= "000000";
					when "01101001001000111" => rgb <= "000000";
					when "01101001001001000" => rgb <= "000000";
					when "01101001001001001" => rgb <= "000000";
					when "01101001001001010" => rgb <= "000000";
					when "01101001001001011" => rgb <= "000000";
					when "01101001001001100" => rgb <= "000000";
					when "01101001001001101" => rgb <= "000000";
					when "01101001001001110" => rgb <= "000000";
					when "01101001001001111" => rgb <= "000000";
					when "01101001001010000" => rgb <= "000000";
					when "01101001001010001" => rgb <= "000000";
					when "01101001001010010" => rgb <= "000000";
					when "01101001001010011" => rgb <= "000000";
					when "01101001001010100" => rgb <= "000000";
					when "01101001001010101" => rgb <= "000000";
					when "01101001001010110" => rgb <= "000000";
					when "01101001001010111" => rgb <= "000000";
					when "01101001001011000" => rgb <= "000000";
					when "01101001001011001" => rgb <= "000000";
					when "01101001001011010" => rgb <= "000000";
					when "01101001001011011" => rgb <= "000000";
					when "01101001001011100" => rgb <= "000000";
					when "01101001001011101" => rgb <= "000000";
					when "01101001001011110" => rgb <= "000000";
					when "01101001001011111" => rgb <= "000000";
					when "01101001001100000" => rgb <= "000000";
					when "01101001001100001" => rgb <= "000000";
					when "01101001001100010" => rgb <= "000000";
					when "01101001001100011" => rgb <= "000000";
					when "01101001001100100" => rgb <= "000000";
					when "01101001001100101" => rgb <= "000000";
					when "01101001001100110" => rgb <= "000000";
					when "01101001001100111" => rgb <= "000000";
					when "01101001001101000" => rgb <= "000000";
					when "01101001001101001" => rgb <= "000000";
					when "01101001001101010" => rgb <= "000000";
					when "01101001001101011" => rgb <= "000000";
					when "01101001001101100" => rgb <= "000000";
					when "01101001001101101" => rgb <= "000000";
					when "01101001001101110" => rgb <= "000000";
					when "01101001001101111" => rgb <= "000000";
					when "01101001001110000" => rgb <= "000000";
					when "01101001001110001" => rgb <= "000000";
					when "01101001001110010" => rgb <= "000000";
					when "01101001001110011" => rgb <= "000000";
					when "01101001001110100" => rgb <= "000000";
					when "01101001001110101" => rgb <= "000000";
					when "01101001001110110" => rgb <= "000000";
					when "01101001001110111" => rgb <= "000000";
					when "01101001001111000" => rgb <= "000000";
					when "01101001001111001" => rgb <= "000000";
					when "01101001001111010" => rgb <= "000000";
					when "01101001001111011" => rgb <= "000000";
					when "01101001001111100" => rgb <= "000000";
					when "01101001001111101" => rgb <= "000000";
					when "01101001001111110" => rgb <= "000000";
					when "01101001001111111" => rgb <= "000000";
					when "01101001010000000" => rgb <= "000000";
					when "01101001010000001" => rgb <= "000000";
					when "01101001010000010" => rgb <= "000000";
					when "01101001010000011" => rgb <= "000000";
					when "01101001010000100" => rgb <= "000000";
					when "01101001010000101" => rgb <= "000000";
					when "01101001010000110" => rgb <= "000000";
					when "01101001010000111" => rgb <= "000000";
					when "01101001010001000" => rgb <= "000000";
					when "01101001010001001" => rgb <= "000000";
					when "01101001010001010" => rgb <= "000000";
					when "01101001010001011" => rgb <= "000000";
					when "01101001010001100" => rgb <= "000000";
					when "01101001010001101" => rgb <= "000000";
					when "01101001010001110" => rgb <= "000000";
					when "01101001010001111" => rgb <= "000000";
					when "01101001010010000" => rgb <= "000000";
					when "01101001010010001" => rgb <= "000000";
					when "01101001010010010" => rgb <= "000000";
					when "01101001010010011" => rgb <= "010000";
					when "01101001010010100" => rgb <= "101000";
					when "01101001010010101" => rgb <= "101000";
					when "01101001010010110" => rgb <= "101000";
					when "01101001010010111" => rgb <= "101000";
					when "01101001010011000" => rgb <= "101000";
					when "01101001010011001" => rgb <= "101000";
					when "01101001010011010" => rgb <= "101000";
					when "01101001010011011" => rgb <= "101000";
					when "01101001010011100" => rgb <= "101000";
					when "01101001010011101" => rgb <= "101000";
					when "01101001010011110" => rgb <= "101000";
					when "01101001010011111" => rgb <= "101000";
					when "01101001010100000" => rgb <= "101000";
					when "01101001010100001" => rgb <= "101000";
					when "01101001010100010" => rgb <= "101000";
					when "01101001010100011" => rgb <= "101000";
					when "01101001010100100" => rgb <= "101000";
					when "01101001010100101" => rgb <= "101000";
					when "01101001010100110" => rgb <= "101000";
					when "01101001010100111" => rgb <= "101000";
					when "01101001010101000" => rgb <= "101000";
					when "01101001010101001" => rgb <= "101000";
					when "01101001010101010" => rgb <= "010000";
					when "01101001010101011" => rgb <= "000000";
					when "01101001010101100" => rgb <= "000000";
					when "01101001010101101" => rgb <= "000000";
					when "01101001010101110" => rgb <= "000000";
					when "01101001010101111" => rgb <= "000000";
					when "01101001010110000" => rgb <= "000000";
					when "01101001010110001" => rgb <= "000000";
					when "01101001010110010" => rgb <= "000000";
					when "01101001010110011" => rgb <= "000000";
					when "01101001010110100" => rgb <= "000000";
					when "01101001010110101" => rgb <= "000000";
					when "01101001010110110" => rgb <= "000000";
					when "01101001010110111" => rgb <= "000000";
					when "01101001010111000" => rgb <= "000000";
					when "01101001010111001" => rgb <= "000000";
					when "01101001010111010" => rgb <= "000000";
					when "01101001010111011" => rgb <= "000000";
					when "01101001010111100" => rgb <= "000000";
					when "01101001010111101" => rgb <= "000000";
					when "01101001010111110" => rgb <= "000000";
					when "01101001010111111" => rgb <= "000000";
					when "01101001011000000" => rgb <= "000000";
					when "01101001011000001" => rgb <= "000000";
					when "01101001011000010" => rgb <= "000000";
					when "01101001011000011" => rgb <= "000000";
					when "01101001011000100" => rgb <= "000000";
					when "01101001011000101" => rgb <= "000000";
					when "01101001011000110" => rgb <= "000000";
					when "01101001011000111" => rgb <= "000000";
					when "01101001011001000" => rgb <= "000000";
					when "01101001011001001" => rgb <= "000000";
					when "01101001011001010" => rgb <= "000000";
					when "01101001011001011" => rgb <= "000000";
					when "01101001011001100" => rgb <= "000000";
					when "01101001011001101" => rgb <= "000000";
					when "01101001011001110" => rgb <= "000000";
					when "01101001011001111" => rgb <= "000000";
					when "01101001011010000" => rgb <= "000000";
					when "01101001011010001" => rgb <= "000000";
					when "01101001011010010" => rgb <= "000000";
					when "01101001011010011" => rgb <= "000000";
					when "01101001011010100" => rgb <= "000000";
					when "01101001011010101" => rgb <= "000000";
					when "01101001011010110" => rgb <= "000000";
					when "01101001011010111" => rgb <= "000000";
					when "01101001011011000" => rgb <= "000000";
					when "01101001011011001" => rgb <= "000000";
					when "01101001011011010" => rgb <= "000000";
					when "01101001011011011" => rgb <= "000000";
					when "01101001011011100" => rgb <= "000000";
					when "01101001011011101" => rgb <= "000000";
					when "01101001011011110" => rgb <= "000000";
					when "01101001011011111" => rgb <= "000000";
					when "01101001011100000" => rgb <= "000000";
					when "01101001011100001" => rgb <= "000000";
					when "01101001011100010" => rgb <= "000000";
					when "01101001011100011" => rgb <= "000000";
					when "01101001011100100" => rgb <= "000000";
					when "01101001011100101" => rgb <= "000000";
					when "01101001011100110" => rgb <= "000000";
					when "01101001011100111" => rgb <= "000000";
					when "01101001011101000" => rgb <= "000000";
					when "01101001011101001" => rgb <= "000000";
					when "01101001011101010" => rgb <= "000000";
					when "01101001011101011" => rgb <= "000000";
					when "01101001011101100" => rgb <= "000000";
					when "01101001011101101" => rgb <= "000000";
					when "01101001011101110" => rgb <= "000000";
					when "01101001011101111" => rgb <= "000000";
					when "01101001011110000" => rgb <= "000000";
					when "01101001011110001" => rgb <= "000000";
					when "01101001011110010" => rgb <= "000000";
					when "01101001011110011" => rgb <= "000000";
					when "01101001011110100" => rgb <= "000000";
					when "01101001011110101" => rgb <= "000000";
					when "01101001011110110" => rgb <= "000000";
					when "01101001011110111" => rgb <= "000000";
					when "01101001011111000" => rgb <= "000000";
					when "01101001011111001" => rgb <= "000000";
					when "01101001011111010" => rgb <= "000000";
					when "01101001011111011" => rgb <= "000000";
					when "01101001011111100" => rgb <= "000000";
					when "01101001011111101" => rgb <= "000000";
					when "01101001011111110" => rgb <= "000000";
					when "01101001011111111" => rgb <= "000000";
					when "01101001100000000" => rgb <= "000000";
					when "01101001100000001" => rgb <= "000000";
					when "01101001100000010" => rgb <= "000000";
					when "01101001100000011" => rgb <= "000000";
					when "01101001100000100" => rgb <= "000000";
					when "01101001100000101" => rgb <= "000000";
					when "01101001100000110" => rgb <= "000000";
					when "01101001100000111" => rgb <= "000000";
					when "01101001100001000" => rgb <= "000000";
					when "01101001100001001" => rgb <= "000000";
					when "01101001100001010" => rgb <= "000000";
					when "01101001100001011" => rgb <= "000000";
					when "01101001100001100" => rgb <= "000000";
					when "01101001100001101" => rgb <= "000000";
					when "01101001100001110" => rgb <= "000000";
					when "01101001100001111" => rgb <= "000000";
					when "01101001100010000" => rgb <= "000000";
					when "01101001100010001" => rgb <= "000000";
					when "01101001100010010" => rgb <= "000000";
					when "01101001100010011" => rgb <= "000000";
					when "01101001100010100" => rgb <= "000000";
					when "01101001100010101" => rgb <= "000000";
					when "01101001100010110" => rgb <= "000000";
					when "01101001100010111" => rgb <= "000000";
					when "01101001100011000" => rgb <= "000000";
					when "01101001100011001" => rgb <= "000000";
					when "01101001100011010" => rgb <= "000000";
					when "01101001100011011" => rgb <= "000000";
					when "01101001100011100" => rgb <= "000000";
					when "01101001100011101" => rgb <= "000000";
					when "01101001100011110" => rgb <= "000000";
					when "01101001100011111" => rgb <= "000000";
					when "01101001100100000" => rgb <= "000000";
					when "01101001100100001" => rgb <= "000000";
					when "01101001100100010" => rgb <= "000000";
					when "01101001100100011" => rgb <= "000000";
					when "01101001100100100" => rgb <= "000000";
					when "01101001100100101" => rgb <= "000000";
					when "01101001100100110" => rgb <= "000000";
					when "01101001100100111" => rgb <= "000000";
					when "01101001100101000" => rgb <= "000000";
					when "01101001100101001" => rgb <= "000000";
					when "01101001100101010" => rgb <= "000000";
					when "01101001100101011" => rgb <= "000000";
					when "01101001100101100" => rgb <= "000000";
					when "01101001100101101" => rgb <= "000000";
					when "01101001100101110" => rgb <= "000000";
					when "01101001100101111" => rgb <= "000000";
					when "01101001100110000" => rgb <= "000000";
					when "01101001100110001" => rgb <= "000000";
					when "01101001100110010" => rgb <= "000000";
					when "01101001100110011" => rgb <= "000000";
					when "01101001100110100" => rgb <= "000000";
					when "01101001100110101" => rgb <= "000000";
					when "01101001100110110" => rgb <= "000000";
					when "01101001100110111" => rgb <= "000000";
					when "01101001100111000" => rgb <= "000000";
					when "01101001100111001" => rgb <= "000000";
					when "01101001100111010" => rgb <= "000000";
					when "01101001100111011" => rgb <= "000000";
					when "01101001100111100" => rgb <= "000000";
					when "01101001100111101" => rgb <= "000000";
					when "01101001100111110" => rgb <= "000000";
					when "01101001100111111" => rgb <= "000000";
					when "01101010000000000" => rgb <= "000000";
					when "01101010000000001" => rgb <= "000000";
					when "01101010000000010" => rgb <= "000000";
					when "01101010000000011" => rgb <= "000000";
					when "01101010000000100" => rgb <= "000000";
					when "01101010000000101" => rgb <= "000000";
					when "01101010000000110" => rgb <= "000000";
					when "01101010000000111" => rgb <= "000000";
					when "01101010000001000" => rgb <= "000000";
					when "01101010000001001" => rgb <= "000000";
					when "01101010000001010" => rgb <= "000000";
					when "01101010000001011" => rgb <= "000000";
					when "01101010000001100" => rgb <= "000000";
					when "01101010000001101" => rgb <= "000000";
					when "01101010000001110" => rgb <= "000000";
					when "01101010000001111" => rgb <= "000000";
					when "01101010000010000" => rgb <= "000000";
					when "01101010000010001" => rgb <= "000000";
					when "01101010000010010" => rgb <= "000000";
					when "01101010000010011" => rgb <= "000000";
					when "01101010000010100" => rgb <= "000000";
					when "01101010000010101" => rgb <= "000000";
					when "01101010000010110" => rgb <= "000000";
					when "01101010000010111" => rgb <= "000000";
					when "01101010000011000" => rgb <= "000000";
					when "01101010000011001" => rgb <= "000000";
					when "01101010000011010" => rgb <= "000000";
					when "01101010000011011" => rgb <= "000000";
					when "01101010000011100" => rgb <= "000000";
					when "01101010000011101" => rgb <= "000000";
					when "01101010000011110" => rgb <= "000000";
					when "01101010000011111" => rgb <= "000000";
					when "01101010000100000" => rgb <= "000000";
					when "01101010000100001" => rgb <= "000000";
					when "01101010000100010" => rgb <= "000000";
					when "01101010000100011" => rgb <= "000000";
					when "01101010000100100" => rgb <= "000000";
					when "01101010000100101" => rgb <= "000000";
					when "01101010000100110" => rgb <= "000000";
					when "01101010000100111" => rgb <= "000000";
					when "01101010000101000" => rgb <= "000000";
					when "01101010000101001" => rgb <= "000000";
					when "01101010000101010" => rgb <= "000000";
					when "01101010000101011" => rgb <= "000000";
					when "01101010000101100" => rgb <= "000000";
					when "01101010000101101" => rgb <= "000000";
					when "01101010000101110" => rgb <= "000000";
					when "01101010000101111" => rgb <= "000000";
					when "01101010000110000" => rgb <= "000000";
					when "01101010000110001" => rgb <= "000000";
					when "01101010000110010" => rgb <= "000000";
					when "01101010000110011" => rgb <= "000000";
					when "01101010000110100" => rgb <= "000000";
					when "01101010000110101" => rgb <= "000000";
					when "01101010000110110" => rgb <= "000000";
					when "01101010000110111" => rgb <= "000000";
					when "01101010000111000" => rgb <= "000000";
					when "01101010000111001" => rgb <= "000000";
					when "01101010000111010" => rgb <= "000000";
					when "01101010000111011" => rgb <= "000000";
					when "01101010000111100" => rgb <= "000000";
					when "01101010000111101" => rgb <= "000000";
					when "01101010000111110" => rgb <= "000000";
					when "01101010000111111" => rgb <= "000000";
					when "01101010001000000" => rgb <= "000000";
					when "01101010001000001" => rgb <= "000000";
					when "01101010001000010" => rgb <= "000000";
					when "01101010001000011" => rgb <= "000000";
					when "01101010001000100" => rgb <= "000000";
					when "01101010001000101" => rgb <= "000000";
					when "01101010001000110" => rgb <= "000000";
					when "01101010001000111" => rgb <= "000000";
					when "01101010001001000" => rgb <= "000000";
					when "01101010001001001" => rgb <= "000000";
					when "01101010001001010" => rgb <= "000000";
					when "01101010001001011" => rgb <= "000000";
					when "01101010001001100" => rgb <= "000000";
					when "01101010001001101" => rgb <= "000000";
					when "01101010001001110" => rgb <= "000000";
					when "01101010001001111" => rgb <= "000000";
					when "01101010001010000" => rgb <= "000000";
					when "01101010001010001" => rgb <= "000000";
					when "01101010001010010" => rgb <= "000000";
					when "01101010001010011" => rgb <= "000000";
					when "01101010001010100" => rgb <= "000000";
					when "01101010001010101" => rgb <= "000000";
					when "01101010001010110" => rgb <= "000000";
					when "01101010001010111" => rgb <= "000000";
					when "01101010001011000" => rgb <= "000000";
					when "01101010001011001" => rgb <= "000000";
					when "01101010001011010" => rgb <= "000000";
					when "01101010001011011" => rgb <= "000000";
					when "01101010001011100" => rgb <= "000000";
					when "01101010001011101" => rgb <= "000000";
					when "01101010001011110" => rgb <= "000000";
					when "01101010001011111" => rgb <= "000000";
					when "01101010001100000" => rgb <= "000000";
					when "01101010001100001" => rgb <= "000000";
					when "01101010001100010" => rgb <= "000000";
					when "01101010001100011" => rgb <= "000000";
					when "01101010001100100" => rgb <= "000000";
					when "01101010001100101" => rgb <= "000000";
					when "01101010001100110" => rgb <= "000000";
					when "01101010001100111" => rgb <= "000000";
					when "01101010001101000" => rgb <= "000000";
					when "01101010001101001" => rgb <= "000000";
					when "01101010001101010" => rgb <= "000000";
					when "01101010001101011" => rgb <= "000000";
					when "01101010001101100" => rgb <= "000000";
					when "01101010001101101" => rgb <= "000000";
					when "01101010001101110" => rgb <= "000000";
					when "01101010001101111" => rgb <= "000000";
					when "01101010001110000" => rgb <= "000000";
					when "01101010001110001" => rgb <= "000000";
					when "01101010001110010" => rgb <= "000000";
					when "01101010001110011" => rgb <= "000000";
					when "01101010001110100" => rgb <= "000000";
					when "01101010001110101" => rgb <= "000000";
					when "01101010001110110" => rgb <= "000000";
					when "01101010001110111" => rgb <= "000000";
					when "01101010001111000" => rgb <= "000000";
					when "01101010001111001" => rgb <= "000000";
					when "01101010001111010" => rgb <= "000000";
					when "01101010001111011" => rgb <= "000000";
					when "01101010001111100" => rgb <= "000000";
					when "01101010001111101" => rgb <= "000000";
					when "01101010001111110" => rgb <= "000000";
					when "01101010001111111" => rgb <= "000000";
					when "01101010010000000" => rgb <= "000000";
					when "01101010010000001" => rgb <= "000000";
					when "01101010010000010" => rgb <= "000000";
					when "01101010010000011" => rgb <= "000000";
					when "01101010010000100" => rgb <= "000000";
					when "01101010010000101" => rgb <= "000000";
					when "01101010010000110" => rgb <= "000000";
					when "01101010010000111" => rgb <= "000000";
					when "01101010010001000" => rgb <= "000000";
					when "01101010010001001" => rgb <= "000000";
					when "01101010010001010" => rgb <= "000000";
					when "01101010010001011" => rgb <= "000000";
					when "01101010010001100" => rgb <= "000000";
					when "01101010010001101" => rgb <= "000000";
					when "01101010010001110" => rgb <= "000000";
					when "01101010010001111" => rgb <= "000000";
					when "01101010010010000" => rgb <= "000000";
					when "01101010010010001" => rgb <= "000000";
					when "01101010010010010" => rgb <= "000000";
					when "01101010010010011" => rgb <= "010000";
					when "01101010010010100" => rgb <= "101000";
					when "01101010010010101" => rgb <= "101000";
					when "01101010010010110" => rgb <= "101000";
					when "01101010010010111" => rgb <= "101000";
					when "01101010010011000" => rgb <= "101000";
					when "01101010010011001" => rgb <= "101000";
					when "01101010010011010" => rgb <= "101000";
					when "01101010010011011" => rgb <= "101000";
					when "01101010010011100" => rgb <= "101000";
					when "01101010010011101" => rgb <= "101000";
					when "01101010010011110" => rgb <= "101000";
					when "01101010010011111" => rgb <= "101000";
					when "01101010010100000" => rgb <= "101000";
					when "01101010010100001" => rgb <= "101000";
					when "01101010010100010" => rgb <= "101000";
					when "01101010010100011" => rgb <= "101000";
					when "01101010010100100" => rgb <= "101000";
					when "01101010010100101" => rgb <= "101000";
					when "01101010010100110" => rgb <= "101000";
					when "01101010010100111" => rgb <= "101000";
					when "01101010010101000" => rgb <= "101000";
					when "01101010010101001" => rgb <= "101000";
					when "01101010010101010" => rgb <= "010000";
					when "01101010010101011" => rgb <= "000000";
					when "01101010010101100" => rgb <= "000000";
					when "01101010010101101" => rgb <= "000000";
					when "01101010010101110" => rgb <= "000000";
					when "01101010010101111" => rgb <= "000000";
					when "01101010010110000" => rgb <= "000000";
					when "01101010010110001" => rgb <= "000000";
					when "01101010010110010" => rgb <= "000000";
					when "01101010010110011" => rgb <= "000000";
					when "01101010010110100" => rgb <= "000000";
					when "01101010010110101" => rgb <= "000000";
					when "01101010010110110" => rgb <= "000000";
					when "01101010010110111" => rgb <= "000000";
					when "01101010010111000" => rgb <= "000000";
					when "01101010010111001" => rgb <= "000000";
					when "01101010010111010" => rgb <= "000000";
					when "01101010010111011" => rgb <= "000000";
					when "01101010010111100" => rgb <= "000000";
					when "01101010010111101" => rgb <= "000000";
					when "01101010010111110" => rgb <= "000000";
					when "01101010010111111" => rgb <= "000000";
					when "01101010011000000" => rgb <= "000000";
					when "01101010011000001" => rgb <= "000000";
					when "01101010011000010" => rgb <= "000000";
					when "01101010011000011" => rgb <= "000000";
					when "01101010011000100" => rgb <= "000000";
					when "01101010011000101" => rgb <= "000000";
					when "01101010011000110" => rgb <= "000000";
					when "01101010011000111" => rgb <= "000000";
					when "01101010011001000" => rgb <= "000000";
					when "01101010011001001" => rgb <= "000000";
					when "01101010011001010" => rgb <= "000000";
					when "01101010011001011" => rgb <= "000000";
					when "01101010011001100" => rgb <= "000000";
					when "01101010011001101" => rgb <= "000000";
					when "01101010011001110" => rgb <= "000000";
					when "01101010011001111" => rgb <= "000000";
					when "01101010011010000" => rgb <= "000000";
					when "01101010011010001" => rgb <= "000000";
					when "01101010011010010" => rgb <= "000000";
					when "01101010011010011" => rgb <= "000000";
					when "01101010011010100" => rgb <= "000000";
					when "01101010011010101" => rgb <= "000000";
					when "01101010011010110" => rgb <= "000000";
					when "01101010011010111" => rgb <= "000000";
					when "01101010011011000" => rgb <= "000000";
					when "01101010011011001" => rgb <= "000000";
					when "01101010011011010" => rgb <= "000000";
					when "01101010011011011" => rgb <= "000000";
					when "01101010011011100" => rgb <= "000000";
					when "01101010011011101" => rgb <= "000000";
					when "01101010011011110" => rgb <= "000000";
					when "01101010011011111" => rgb <= "000000";
					when "01101010011100000" => rgb <= "000000";
					when "01101010011100001" => rgb <= "000000";
					when "01101010011100010" => rgb <= "000000";
					when "01101010011100011" => rgb <= "000000";
					when "01101010011100100" => rgb <= "000000";
					when "01101010011100101" => rgb <= "000000";
					when "01101010011100110" => rgb <= "000000";
					when "01101010011100111" => rgb <= "000000";
					when "01101010011101000" => rgb <= "000000";
					when "01101010011101001" => rgb <= "000000";
					when "01101010011101010" => rgb <= "000000";
					when "01101010011101011" => rgb <= "000000";
					when "01101010011101100" => rgb <= "000000";
					when "01101010011101101" => rgb <= "000000";
					when "01101010011101110" => rgb <= "000000";
					when "01101010011101111" => rgb <= "000000";
					when "01101010011110000" => rgb <= "000000";
					when "01101010011110001" => rgb <= "000000";
					when "01101010011110010" => rgb <= "000000";
					when "01101010011110011" => rgb <= "000000";
					when "01101010011110100" => rgb <= "000000";
					when "01101010011110101" => rgb <= "000000";
					when "01101010011110110" => rgb <= "000000";
					when "01101010011110111" => rgb <= "000000";
					when "01101010011111000" => rgb <= "000000";
					when "01101010011111001" => rgb <= "000000";
					when "01101010011111010" => rgb <= "000000";
					when "01101010011111011" => rgb <= "000000";
					when "01101010011111100" => rgb <= "000000";
					when "01101010011111101" => rgb <= "000000";
					when "01101010011111110" => rgb <= "000000";
					when "01101010011111111" => rgb <= "000000";
					when "01101010100000000" => rgb <= "000000";
					when "01101010100000001" => rgb <= "000000";
					when "01101010100000010" => rgb <= "000000";
					when "01101010100000011" => rgb <= "000000";
					when "01101010100000100" => rgb <= "000000";
					when "01101010100000101" => rgb <= "000000";
					when "01101010100000110" => rgb <= "000000";
					when "01101010100000111" => rgb <= "000000";
					when "01101010100001000" => rgb <= "000000";
					when "01101010100001001" => rgb <= "000000";
					when "01101010100001010" => rgb <= "000000";
					when "01101010100001011" => rgb <= "000000";
					when "01101010100001100" => rgb <= "000000";
					when "01101010100001101" => rgb <= "000000";
					when "01101010100001110" => rgb <= "000000";
					when "01101010100001111" => rgb <= "000000";
					when "01101010100010000" => rgb <= "000000";
					when "01101010100010001" => rgb <= "000000";
					when "01101010100010010" => rgb <= "000000";
					when "01101010100010011" => rgb <= "000000";
					when "01101010100010100" => rgb <= "000000";
					when "01101010100010101" => rgb <= "000000";
					when "01101010100010110" => rgb <= "000000";
					when "01101010100010111" => rgb <= "000000";
					when "01101010100011000" => rgb <= "000000";
					when "01101010100011001" => rgb <= "000000";
					when "01101010100011010" => rgb <= "000000";
					when "01101010100011011" => rgb <= "000000";
					when "01101010100011100" => rgb <= "000000";
					when "01101010100011101" => rgb <= "000000";
					when "01101010100011110" => rgb <= "000000";
					when "01101010100011111" => rgb <= "000000";
					when "01101010100100000" => rgb <= "000000";
					when "01101010100100001" => rgb <= "000000";
					when "01101010100100010" => rgb <= "000000";
					when "01101010100100011" => rgb <= "000000";
					when "01101010100100100" => rgb <= "000000";
					when "01101010100100101" => rgb <= "000000";
					when "01101010100100110" => rgb <= "000000";
					when "01101010100100111" => rgb <= "000000";
					when "01101010100101000" => rgb <= "000000";
					when "01101010100101001" => rgb <= "000000";
					when "01101010100101010" => rgb <= "000000";
					when "01101010100101011" => rgb <= "000000";
					when "01101010100101100" => rgb <= "000000";
					when "01101010100101101" => rgb <= "000000";
					when "01101010100101110" => rgb <= "000000";
					when "01101010100101111" => rgb <= "000000";
					when "01101010100110000" => rgb <= "000000";
					when "01101010100110001" => rgb <= "000000";
					when "01101010100110010" => rgb <= "000000";
					when "01101010100110011" => rgb <= "000000";
					when "01101010100110100" => rgb <= "000000";
					when "01101010100110101" => rgb <= "000000";
					when "01101010100110110" => rgb <= "000000";
					when "01101010100110111" => rgb <= "000000";
					when "01101010100111000" => rgb <= "000000";
					when "01101010100111001" => rgb <= "000000";
					when "01101010100111010" => rgb <= "000000";
					when "01101010100111011" => rgb <= "000000";
					when "01101010100111100" => rgb <= "000000";
					when "01101010100111101" => rgb <= "000000";
					when "01101010100111110" => rgb <= "000000";
					when "01101010100111111" => rgb <= "000000";
					when "01101011000000000" => rgb <= "000000";
					when "01101011000000001" => rgb <= "000000";
					when "01101011000000010" => rgb <= "000000";
					when "01101011000000011" => rgb <= "000000";
					when "01101011000000100" => rgb <= "000000";
					when "01101011000000101" => rgb <= "000000";
					when "01101011000000110" => rgb <= "000000";
					when "01101011000000111" => rgb <= "000000";
					when "01101011000001000" => rgb <= "000000";
					when "01101011000001001" => rgb <= "000000";
					when "01101011000001010" => rgb <= "000000";
					when "01101011000001011" => rgb <= "000000";
					when "01101011000001100" => rgb <= "000000";
					when "01101011000001101" => rgb <= "000000";
					when "01101011000001110" => rgb <= "000000";
					when "01101011000001111" => rgb <= "000000";
					when "01101011000010000" => rgb <= "000000";
					when "01101011000010001" => rgb <= "000000";
					when "01101011000010010" => rgb <= "000000";
					when "01101011000010011" => rgb <= "000000";
					when "01101011000010100" => rgb <= "000000";
					when "01101011000010101" => rgb <= "000000";
					when "01101011000010110" => rgb <= "000000";
					when "01101011000010111" => rgb <= "000000";
					when "01101011000011000" => rgb <= "000000";
					when "01101011000011001" => rgb <= "000000";
					when "01101011000011010" => rgb <= "000000";
					when "01101011000011011" => rgb <= "000000";
					when "01101011000011100" => rgb <= "000000";
					when "01101011000011101" => rgb <= "000000";
					when "01101011000011110" => rgb <= "000000";
					when "01101011000011111" => rgb <= "000000";
					when "01101011000100000" => rgb <= "000000";
					when "01101011000100001" => rgb <= "000000";
					when "01101011000100010" => rgb <= "000000";
					when "01101011000100011" => rgb <= "000000";
					when "01101011000100100" => rgb <= "000000";
					when "01101011000100101" => rgb <= "000000";
					when "01101011000100110" => rgb <= "000000";
					when "01101011000100111" => rgb <= "000000";
					when "01101011000101000" => rgb <= "000000";
					when "01101011000101001" => rgb <= "000000";
					when "01101011000101010" => rgb <= "000000";
					when "01101011000101011" => rgb <= "000000";
					when "01101011000101100" => rgb <= "000000";
					when "01101011000101101" => rgb <= "000000";
					when "01101011000101110" => rgb <= "000000";
					when "01101011000101111" => rgb <= "000000";
					when "01101011000110000" => rgb <= "000000";
					when "01101011000110001" => rgb <= "000000";
					when "01101011000110010" => rgb <= "000000";
					when "01101011000110011" => rgb <= "000000";
					when "01101011000110100" => rgb <= "000000";
					when "01101011000110101" => rgb <= "000000";
					when "01101011000110110" => rgb <= "000000";
					when "01101011000110111" => rgb <= "000000";
					when "01101011000111000" => rgb <= "000000";
					when "01101011000111001" => rgb <= "000000";
					when "01101011000111010" => rgb <= "000000";
					when "01101011000111011" => rgb <= "000000";
					when "01101011000111100" => rgb <= "000000";
					when "01101011000111101" => rgb <= "000000";
					when "01101011000111110" => rgb <= "000000";
					when "01101011000111111" => rgb <= "000000";
					when "01101011001000000" => rgb <= "000000";
					when "01101011001000001" => rgb <= "000000";
					when "01101011001000010" => rgb <= "000000";
					when "01101011001000011" => rgb <= "000000";
					when "01101011001000100" => rgb <= "000000";
					when "01101011001000101" => rgb <= "000000";
					when "01101011001000110" => rgb <= "000000";
					when "01101011001000111" => rgb <= "000000";
					when "01101011001001000" => rgb <= "000000";
					when "01101011001001001" => rgb <= "000000";
					when "01101011001001010" => rgb <= "000000";
					when "01101011001001011" => rgb <= "000000";
					when "01101011001001100" => rgb <= "000000";
					when "01101011001001101" => rgb <= "000000";
					when "01101011001001110" => rgb <= "000000";
					when "01101011001001111" => rgb <= "000000";
					when "01101011001010000" => rgb <= "000000";
					when "01101011001010001" => rgb <= "000000";
					when "01101011001010010" => rgb <= "000000";
					when "01101011001010011" => rgb <= "000000";
					when "01101011001010100" => rgb <= "000000";
					when "01101011001010101" => rgb <= "000000";
					when "01101011001010110" => rgb <= "000000";
					when "01101011001010111" => rgb <= "000000";
					when "01101011001011000" => rgb <= "000000";
					when "01101011001011001" => rgb <= "000000";
					when "01101011001011010" => rgb <= "000000";
					when "01101011001011011" => rgb <= "000000";
					when "01101011001011100" => rgb <= "000000";
					when "01101011001011101" => rgb <= "000000";
					when "01101011001011110" => rgb <= "000000";
					when "01101011001011111" => rgb <= "000000";
					when "01101011001100000" => rgb <= "000000";
					when "01101011001100001" => rgb <= "000000";
					when "01101011001100010" => rgb <= "000000";
					when "01101011001100011" => rgb <= "000000";
					when "01101011001100100" => rgb <= "000000";
					when "01101011001100101" => rgb <= "000000";
					when "01101011001100110" => rgb <= "000000";
					when "01101011001100111" => rgb <= "000000";
					when "01101011001101000" => rgb <= "000000";
					when "01101011001101001" => rgb <= "000000";
					when "01101011001101010" => rgb <= "000000";
					when "01101011001101011" => rgb <= "000000";
					when "01101011001101100" => rgb <= "000000";
					when "01101011001101101" => rgb <= "000000";
					when "01101011001101110" => rgb <= "000000";
					when "01101011001101111" => rgb <= "000000";
					when "01101011001110000" => rgb <= "000000";
					when "01101011001110001" => rgb <= "000000";
					when "01101011001110010" => rgb <= "000000";
					when "01101011001110011" => rgb <= "000000";
					when "01101011001110100" => rgb <= "000000";
					when "01101011001110101" => rgb <= "000000";
					when "01101011001110110" => rgb <= "000000";
					when "01101011001110111" => rgb <= "000000";
					when "01101011001111000" => rgb <= "000000";
					when "01101011001111001" => rgb <= "000000";
					when "01101011001111010" => rgb <= "000000";
					when "01101011001111011" => rgb <= "000000";
					when "01101011001111100" => rgb <= "000000";
					when "01101011001111101" => rgb <= "000000";
					when "01101011001111110" => rgb <= "000000";
					when "01101011001111111" => rgb <= "000000";
					when "01101011010000000" => rgb <= "000000";
					when "01101011010000001" => rgb <= "000000";
					when "01101011010000010" => rgb <= "000000";
					when "01101011010000011" => rgb <= "000000";
					when "01101011010000100" => rgb <= "000000";
					when "01101011010000101" => rgb <= "000000";
					when "01101011010000110" => rgb <= "000000";
					when "01101011010000111" => rgb <= "000000";
					when "01101011010001000" => rgb <= "000000";
					when "01101011010001001" => rgb <= "000000";
					when "01101011010001010" => rgb <= "000000";
					when "01101011010001011" => rgb <= "000000";
					when "01101011010001100" => rgb <= "000000";
					when "01101011010001101" => rgb <= "000000";
					when "01101011010001110" => rgb <= "000000";
					when "01101011010001111" => rgb <= "000000";
					when "01101011010010000" => rgb <= "000000";
					when "01101011010010001" => rgb <= "000000";
					when "01101011010010010" => rgb <= "000000";
					when "01101011010010011" => rgb <= "010100";
					when "01101011010010100" => rgb <= "101000";
					when "01101011010010101" => rgb <= "101000";
					when "01101011010010110" => rgb <= "101000";
					when "01101011010010111" => rgb <= "101000";
					when "01101011010011000" => rgb <= "101000";
					when "01101011010011001" => rgb <= "101000";
					when "01101011010011010" => rgb <= "101000";
					when "01101011010011011" => rgb <= "101000";
					when "01101011010011100" => rgb <= "101000";
					when "01101011010011101" => rgb <= "101000";
					when "01101011010011110" => rgb <= "101000";
					when "01101011010011111" => rgb <= "101000";
					when "01101011010100000" => rgb <= "101000";
					when "01101011010100001" => rgb <= "101000";
					when "01101011010100010" => rgb <= "101000";
					when "01101011010100011" => rgb <= "101000";
					when "01101011010100100" => rgb <= "101000";
					when "01101011010100101" => rgb <= "101000";
					when "01101011010100110" => rgb <= "101000";
					when "01101011010100111" => rgb <= "101000";
					when "01101011010101000" => rgb <= "101000";
					when "01101011010101001" => rgb <= "101000";
					when "01101011010101010" => rgb <= "010100";
					when "01101011010101011" => rgb <= "000000";
					when "01101011010101100" => rgb <= "000000";
					when "01101011010101101" => rgb <= "000000";
					when "01101011010101110" => rgb <= "010000";
					when "01101011010101111" => rgb <= "000000";
					when "01101011010110000" => rgb <= "000000";
					when "01101011010110001" => rgb <= "000000";
					when "01101011010110010" => rgb <= "000000";
					when "01101011010110011" => rgb <= "000000";
					when "01101011010110100" => rgb <= "010000";
					when "01101011010110101" => rgb <= "000000";
					when "01101011010110110" => rgb <= "000000";
					when "01101011010110111" => rgb <= "000000";
					when "01101011010111000" => rgb <= "000000";
					when "01101011010111001" => rgb <= "000000";
					when "01101011010111010" => rgb <= "000000";
					when "01101011010111011" => rgb <= "000000";
					when "01101011010111100" => rgb <= "000000";
					when "01101011010111101" => rgb <= "000000";
					when "01101011010111110" => rgb <= "000000";
					when "01101011010111111" => rgb <= "000000";
					when "01101011011000000" => rgb <= "000000";
					when "01101011011000001" => rgb <= "000000";
					when "01101011011000010" => rgb <= "000000";
					when "01101011011000011" => rgb <= "000000";
					when "01101011011000100" => rgb <= "000000";
					when "01101011011000101" => rgb <= "000000";
					when "01101011011000110" => rgb <= "000000";
					when "01101011011000111" => rgb <= "000000";
					when "01101011011001000" => rgb <= "000000";
					when "01101011011001001" => rgb <= "000000";
					when "01101011011001010" => rgb <= "000000";
					when "01101011011001011" => rgb <= "000000";
					when "01101011011001100" => rgb <= "000000";
					when "01101011011001101" => rgb <= "000000";
					when "01101011011001110" => rgb <= "000000";
					when "01101011011001111" => rgb <= "000000";
					when "01101011011010000" => rgb <= "000000";
					when "01101011011010001" => rgb <= "000000";
					when "01101011011010010" => rgb <= "000000";
					when "01101011011010011" => rgb <= "000000";
					when "01101011011010100" => rgb <= "000000";
					when "01101011011010101" => rgb <= "000000";
					when "01101011011010110" => rgb <= "000000";
					when "01101011011010111" => rgb <= "000000";
					when "01101011011011000" => rgb <= "000000";
					when "01101011011011001" => rgb <= "000000";
					when "01101011011011010" => rgb <= "000000";
					when "01101011011011011" => rgb <= "000000";
					when "01101011011011100" => rgb <= "000000";
					when "01101011011011101" => rgb <= "000000";
					when "01101011011011110" => rgb <= "000000";
					when "01101011011011111" => rgb <= "000000";
					when "01101011011100000" => rgb <= "000000";
					when "01101011011100001" => rgb <= "000000";
					when "01101011011100010" => rgb <= "000000";
					when "01101011011100011" => rgb <= "000000";
					when "01101011011100100" => rgb <= "000000";
					when "01101011011100101" => rgb <= "000000";
					when "01101011011100110" => rgb <= "000000";
					when "01101011011100111" => rgb <= "000000";
					when "01101011011101000" => rgb <= "000000";
					when "01101011011101001" => rgb <= "000000";
					when "01101011011101010" => rgb <= "000000";
					when "01101011011101011" => rgb <= "000000";
					when "01101011011101100" => rgb <= "000000";
					when "01101011011101101" => rgb <= "000000";
					when "01101011011101110" => rgb <= "000000";
					when "01101011011101111" => rgb <= "000000";
					when "01101011011110000" => rgb <= "000000";
					when "01101011011110001" => rgb <= "000000";
					when "01101011011110010" => rgb <= "000000";
					when "01101011011110011" => rgb <= "000000";
					when "01101011011110100" => rgb <= "000000";
					when "01101011011110101" => rgb <= "000000";
					when "01101011011110110" => rgb <= "000000";
					when "01101011011110111" => rgb <= "000000";
					when "01101011011111000" => rgb <= "000000";
					when "01101011011111001" => rgb <= "000000";
					when "01101011011111010" => rgb <= "000000";
					when "01101011011111011" => rgb <= "000000";
					when "01101011011111100" => rgb <= "000000";
					when "01101011011111101" => rgb <= "000000";
					when "01101011011111110" => rgb <= "000000";
					when "01101011011111111" => rgb <= "000000";
					when "01101011100000000" => rgb <= "000000";
					when "01101011100000001" => rgb <= "000000";
					when "01101011100000010" => rgb <= "000000";
					when "01101011100000011" => rgb <= "000000";
					when "01101011100000100" => rgb <= "000000";
					when "01101011100000101" => rgb <= "000000";
					when "01101011100000110" => rgb <= "000000";
					when "01101011100000111" => rgb <= "000000";
					when "01101011100001000" => rgb <= "000000";
					when "01101011100001001" => rgb <= "000000";
					when "01101011100001010" => rgb <= "000000";
					when "01101011100001011" => rgb <= "000000";
					when "01101011100001100" => rgb <= "000000";
					when "01101011100001101" => rgb <= "000000";
					when "01101011100001110" => rgb <= "000000";
					when "01101011100001111" => rgb <= "000000";
					when "01101011100010000" => rgb <= "000000";
					when "01101011100010001" => rgb <= "000000";
					when "01101011100010010" => rgb <= "000000";
					when "01101011100010011" => rgb <= "000000";
					when "01101011100010100" => rgb <= "000000";
					when "01101011100010101" => rgb <= "000000";
					when "01101011100010110" => rgb <= "000000";
					when "01101011100010111" => rgb <= "000000";
					when "01101011100011000" => rgb <= "000000";
					when "01101011100011001" => rgb <= "000000";
					when "01101011100011010" => rgb <= "000000";
					when "01101011100011011" => rgb <= "000000";
					when "01101011100011100" => rgb <= "000000";
					when "01101011100011101" => rgb <= "000000";
					when "01101011100011110" => rgb <= "000000";
					when "01101011100011111" => rgb <= "000000";
					when "01101011100100000" => rgb <= "000000";
					when "01101011100100001" => rgb <= "000000";
					when "01101011100100010" => rgb <= "000000";
					when "01101011100100011" => rgb <= "000000";
					when "01101011100100100" => rgb <= "000000";
					when "01101011100100101" => rgb <= "000000";
					when "01101011100100110" => rgb <= "000000";
					when "01101011100100111" => rgb <= "000000";
					when "01101011100101000" => rgb <= "000000";
					when "01101011100101001" => rgb <= "000000";
					when "01101011100101010" => rgb <= "000000";
					when "01101011100101011" => rgb <= "000000";
					when "01101011100101100" => rgb <= "000000";
					when "01101011100101101" => rgb <= "000000";
					when "01101011100101110" => rgb <= "000000";
					when "01101011100101111" => rgb <= "000000";
					when "01101011100110000" => rgb <= "000000";
					when "01101011100110001" => rgb <= "000000";
					when "01101011100110010" => rgb <= "000000";
					when "01101011100110011" => rgb <= "000000";
					when "01101011100110100" => rgb <= "000000";
					when "01101011100110101" => rgb <= "000000";
					when "01101011100110110" => rgb <= "000000";
					when "01101011100110111" => rgb <= "000000";
					when "01101011100111000" => rgb <= "000000";
					when "01101011100111001" => rgb <= "000000";
					when "01101011100111010" => rgb <= "000000";
					when "01101011100111011" => rgb <= "000000";
					when "01101011100111100" => rgb <= "000000";
					when "01101011100111101" => rgb <= "000000";
					when "01101011100111110" => rgb <= "000000";
					when "01101011100111111" => rgb <= "000000";
					when "01101100000000000" => rgb <= "000000";
					when "01101100000000001" => rgb <= "000000";
					when "01101100000000010" => rgb <= "000000";
					when "01101100000000011" => rgb <= "000000";
					when "01101100000000100" => rgb <= "000000";
					when "01101100000000101" => rgb <= "000000";
					when "01101100000000110" => rgb <= "000000";
					when "01101100000000111" => rgb <= "000000";
					when "01101100000001000" => rgb <= "000000";
					when "01101100000001001" => rgb <= "000000";
					when "01101100000001010" => rgb <= "000000";
					when "01101100000001011" => rgb <= "000000";
					when "01101100000001100" => rgb <= "000000";
					when "01101100000001101" => rgb <= "000000";
					when "01101100000001110" => rgb <= "000000";
					when "01101100000001111" => rgb <= "000000";
					when "01101100000010000" => rgb <= "000000";
					when "01101100000010001" => rgb <= "000000";
					when "01101100000010010" => rgb <= "000000";
					when "01101100000010011" => rgb <= "000000";
					when "01101100000010100" => rgb <= "000000";
					when "01101100000010101" => rgb <= "000000";
					when "01101100000010110" => rgb <= "000000";
					when "01101100000010111" => rgb <= "000000";
					when "01101100000011000" => rgb <= "000000";
					when "01101100000011001" => rgb <= "000000";
					when "01101100000011010" => rgb <= "000000";
					when "01101100000011011" => rgb <= "000000";
					when "01101100000011100" => rgb <= "000000";
					when "01101100000011101" => rgb <= "000000";
					when "01101100000011110" => rgb <= "000000";
					when "01101100000011111" => rgb <= "000000";
					when "01101100000100000" => rgb <= "000000";
					when "01101100000100001" => rgb <= "000000";
					when "01101100000100010" => rgb <= "000000";
					when "01101100000100011" => rgb <= "000000";
					when "01101100000100100" => rgb <= "000000";
					when "01101100000100101" => rgb <= "000000";
					when "01101100000100110" => rgb <= "000000";
					when "01101100000100111" => rgb <= "000000";
					when "01101100000101000" => rgb <= "000000";
					when "01101100000101001" => rgb <= "000000";
					when "01101100000101010" => rgb <= "000000";
					when "01101100000101011" => rgb <= "000000";
					when "01101100000101100" => rgb <= "000000";
					when "01101100000101101" => rgb <= "000000";
					when "01101100000101110" => rgb <= "000000";
					when "01101100000101111" => rgb <= "000000";
					when "01101100000110000" => rgb <= "000000";
					when "01101100000110001" => rgb <= "000000";
					when "01101100000110010" => rgb <= "000000";
					when "01101100000110011" => rgb <= "000000";
					when "01101100000110100" => rgb <= "000000";
					when "01101100000110101" => rgb <= "000000";
					when "01101100000110110" => rgb <= "000000";
					when "01101100000110111" => rgb <= "000000";
					when "01101100000111000" => rgb <= "000000";
					when "01101100000111001" => rgb <= "000000";
					when "01101100000111010" => rgb <= "000000";
					when "01101100000111011" => rgb <= "000000";
					when "01101100000111100" => rgb <= "000000";
					when "01101100000111101" => rgb <= "000000";
					when "01101100000111110" => rgb <= "000000";
					when "01101100000111111" => rgb <= "000000";
					when "01101100001000000" => rgb <= "000000";
					when "01101100001000001" => rgb <= "000000";
					when "01101100001000010" => rgb <= "000000";
					when "01101100001000011" => rgb <= "000000";
					when "01101100001000100" => rgb <= "000000";
					when "01101100001000101" => rgb <= "000000";
					when "01101100001000110" => rgb <= "000000";
					when "01101100001000111" => rgb <= "000000";
					when "01101100001001000" => rgb <= "000000";
					when "01101100001001001" => rgb <= "000000";
					when "01101100001001010" => rgb <= "000000";
					when "01101100001001011" => rgb <= "000000";
					when "01101100001001100" => rgb <= "000000";
					when "01101100001001101" => rgb <= "000000";
					when "01101100001001110" => rgb <= "000000";
					when "01101100001001111" => rgb <= "000000";
					when "01101100001010000" => rgb <= "000000";
					when "01101100001010001" => rgb <= "000000";
					when "01101100001010010" => rgb <= "000000";
					when "01101100001010011" => rgb <= "000000";
					when "01101100001010100" => rgb <= "000000";
					when "01101100001010101" => rgb <= "000000";
					when "01101100001010110" => rgb <= "000000";
					when "01101100001010111" => rgb <= "000000";
					when "01101100001011000" => rgb <= "000000";
					when "01101100001011001" => rgb <= "000000";
					when "01101100001011010" => rgb <= "000000";
					when "01101100001011011" => rgb <= "000000";
					when "01101100001011100" => rgb <= "000000";
					when "01101100001011101" => rgb <= "000000";
					when "01101100001011110" => rgb <= "000000";
					when "01101100001011111" => rgb <= "000000";
					when "01101100001100000" => rgb <= "000000";
					when "01101100001100001" => rgb <= "000000";
					when "01101100001100010" => rgb <= "000000";
					when "01101100001100011" => rgb <= "000000";
					when "01101100001100100" => rgb <= "000000";
					when "01101100001100101" => rgb <= "000000";
					when "01101100001100110" => rgb <= "000000";
					when "01101100001100111" => rgb <= "000000";
					when "01101100001101000" => rgb <= "000000";
					when "01101100001101001" => rgb <= "000000";
					when "01101100001101010" => rgb <= "000000";
					when "01101100001101011" => rgb <= "000000";
					when "01101100001101100" => rgb <= "000000";
					when "01101100001101101" => rgb <= "000000";
					when "01101100001101110" => rgb <= "000000";
					when "01101100001101111" => rgb <= "000000";
					when "01101100001110000" => rgb <= "000000";
					when "01101100001110001" => rgb <= "000000";
					when "01101100001110010" => rgb <= "000000";
					when "01101100001110011" => rgb <= "000000";
					when "01101100001110100" => rgb <= "000000";
					when "01101100001110101" => rgb <= "000000";
					when "01101100001110110" => rgb <= "000000";
					when "01101100001110111" => rgb <= "000000";
					when "01101100001111000" => rgb <= "000000";
					when "01101100001111001" => rgb <= "000000";
					when "01101100001111010" => rgb <= "000000";
					when "01101100001111011" => rgb <= "000000";
					when "01101100001111100" => rgb <= "000000";
					when "01101100001111101" => rgb <= "000000";
					when "01101100001111110" => rgb <= "000000";
					when "01101100001111111" => rgb <= "000000";
					when "01101100010000000" => rgb <= "000000";
					when "01101100010000001" => rgb <= "000000";
					when "01101100010000010" => rgb <= "000000";
					when "01101100010000011" => rgb <= "000000";
					when "01101100010000100" => rgb <= "000000";
					when "01101100010000101" => rgb <= "000000";
					when "01101100010000110" => rgb <= "000000";
					when "01101100010000111" => rgb <= "000000";
					when "01101100010001000" => rgb <= "100100";
					when "01101100010001001" => rgb <= "101000";
					when "01101100010001010" => rgb <= "101000";
					when "01101100010001011" => rgb <= "101000";
					when "01101100010001100" => rgb <= "101000";
					when "01101100010001101" => rgb <= "101000";
					when "01101100010001110" => rgb <= "101000";
					when "01101100010001111" => rgb <= "101000";
					when "01101100010010000" => rgb <= "101000";
					when "01101100010010001" => rgb <= "101000";
					when "01101100010010010" => rgb <= "101000";
					when "01101100010010011" => rgb <= "101000";
					when "01101100010010100" => rgb <= "101000";
					when "01101100010010101" => rgb <= "101000";
					when "01101100010010110" => rgb <= "101000";
					when "01101100010010111" => rgb <= "101000";
					when "01101100010011000" => rgb <= "101000";
					when "01101100010011001" => rgb <= "101000";
					when "01101100010011010" => rgb <= "101000";
					when "01101100010011011" => rgb <= "101000";
					when "01101100010011100" => rgb <= "101000";
					when "01101100010011101" => rgb <= "101000";
					when "01101100010011110" => rgb <= "101000";
					when "01101100010011111" => rgb <= "101000";
					when "01101100010100000" => rgb <= "101000";
					when "01101100010100001" => rgb <= "101000";
					when "01101100010100010" => rgb <= "101000";
					when "01101100010100011" => rgb <= "101000";
					when "01101100010100100" => rgb <= "101000";
					when "01101100010100101" => rgb <= "101000";
					when "01101100010100110" => rgb <= "101000";
					when "01101100010100111" => rgb <= "101000";
					when "01101100010101000" => rgb <= "101000";
					when "01101100010101001" => rgb <= "101000";
					when "01101100010101010" => rgb <= "101000";
					when "01101100010101011" => rgb <= "101000";
					when "01101100010101100" => rgb <= "101000";
					when "01101100010101101" => rgb <= "101000";
					when "01101100010101110" => rgb <= "101000";
					when "01101100010101111" => rgb <= "101000";
					when "01101100010110000" => rgb <= "101000";
					when "01101100010110001" => rgb <= "101000";
					when "01101100010110010" => rgb <= "101000";
					when "01101100010110011" => rgb <= "101000";
					when "01101100010110100" => rgb <= "101000";
					when "01101100010110101" => rgb <= "010100";
					when "01101100010110110" => rgb <= "000000";
					when "01101100010110111" => rgb <= "000000";
					when "01101100010111000" => rgb <= "000000";
					when "01101100010111001" => rgb <= "000000";
					when "01101100010111010" => rgb <= "000000";
					when "01101100010111011" => rgb <= "000000";
					when "01101100010111100" => rgb <= "000000";
					when "01101100010111101" => rgb <= "000000";
					when "01101100010111110" => rgb <= "000000";
					when "01101100010111111" => rgb <= "000000";
					when "01101100011000000" => rgb <= "000000";
					when "01101100011000001" => rgb <= "000000";
					when "01101100011000010" => rgb <= "000000";
					when "01101100011000011" => rgb <= "000000";
					when "01101100011000100" => rgb <= "000000";
					when "01101100011000101" => rgb <= "000000";
					when "01101100011000110" => rgb <= "000000";
					when "01101100011000111" => rgb <= "000000";
					when "01101100011001000" => rgb <= "000000";
					when "01101100011001001" => rgb <= "000000";
					when "01101100011001010" => rgb <= "000000";
					when "01101100011001011" => rgb <= "000000";
					when "01101100011001100" => rgb <= "000000";
					when "01101100011001101" => rgb <= "000000";
					when "01101100011001110" => rgb <= "000000";
					when "01101100011001111" => rgb <= "000000";
					when "01101100011010000" => rgb <= "000000";
					when "01101100011010001" => rgb <= "000000";
					when "01101100011010010" => rgb <= "000000";
					when "01101100011010011" => rgb <= "000000";
					when "01101100011010100" => rgb <= "000000";
					when "01101100011010101" => rgb <= "000000";
					when "01101100011010110" => rgb <= "000000";
					when "01101100011010111" => rgb <= "000000";
					when "01101100011011000" => rgb <= "000000";
					when "01101100011011001" => rgb <= "000000";
					when "01101100011011010" => rgb <= "000000";
					when "01101100011011011" => rgb <= "000000";
					when "01101100011011100" => rgb <= "000000";
					when "01101100011011101" => rgb <= "000000";
					when "01101100011011110" => rgb <= "000000";
					when "01101100011011111" => rgb <= "000000";
					when "01101100011100000" => rgb <= "000000";
					when "01101100011100001" => rgb <= "000000";
					when "01101100011100010" => rgb <= "000000";
					when "01101100011100011" => rgb <= "000000";
					when "01101100011100100" => rgb <= "000000";
					when "01101100011100101" => rgb <= "000000";
					when "01101100011100110" => rgb <= "000000";
					when "01101100011100111" => rgb <= "000000";
					when "01101100011101000" => rgb <= "000000";
					when "01101100011101001" => rgb <= "000000";
					when "01101100011101010" => rgb <= "000000";
					when "01101100011101011" => rgb <= "000000";
					when "01101100011101100" => rgb <= "000000";
					when "01101100011101101" => rgb <= "000000";
					when "01101100011101110" => rgb <= "000000";
					when "01101100011101111" => rgb <= "000000";
					when "01101100011110000" => rgb <= "000000";
					when "01101100011110001" => rgb <= "000000";
					when "01101100011110010" => rgb <= "000000";
					when "01101100011110011" => rgb <= "000000";
					when "01101100011110100" => rgb <= "000000";
					when "01101100011110101" => rgb <= "000000";
					when "01101100011110110" => rgb <= "000000";
					when "01101100011110111" => rgb <= "000000";
					when "01101100011111000" => rgb <= "000000";
					when "01101100011111001" => rgb <= "000000";
					when "01101100011111010" => rgb <= "000000";
					when "01101100011111011" => rgb <= "000000";
					when "01101100011111100" => rgb <= "000000";
					when "01101100011111101" => rgb <= "000000";
					when "01101100011111110" => rgb <= "000000";
					when "01101100011111111" => rgb <= "000000";
					when "01101100100000000" => rgb <= "000000";
					when "01101100100000001" => rgb <= "000000";
					when "01101100100000010" => rgb <= "000000";
					when "01101100100000011" => rgb <= "000000";
					when "01101100100000100" => rgb <= "000000";
					when "01101100100000101" => rgb <= "000000";
					when "01101100100000110" => rgb <= "000000";
					when "01101100100000111" => rgb <= "000000";
					when "01101100100001000" => rgb <= "000000";
					when "01101100100001001" => rgb <= "000000";
					when "01101100100001010" => rgb <= "000000";
					when "01101100100001011" => rgb <= "000000";
					when "01101100100001100" => rgb <= "000000";
					when "01101100100001101" => rgb <= "000000";
					when "01101100100001110" => rgb <= "000000";
					when "01101100100001111" => rgb <= "000000";
					when "01101100100010000" => rgb <= "000000";
					when "01101100100010001" => rgb <= "000000";
					when "01101100100010010" => rgb <= "000000";
					when "01101100100010011" => rgb <= "000000";
					when "01101100100010100" => rgb <= "000000";
					when "01101100100010101" => rgb <= "000000";
					when "01101100100010110" => rgb <= "000000";
					when "01101100100010111" => rgb <= "000000";
					when "01101100100011000" => rgb <= "000000";
					when "01101100100011001" => rgb <= "000000";
					when "01101100100011010" => rgb <= "000000";
					when "01101100100011011" => rgb <= "000000";
					when "01101100100011100" => rgb <= "000000";
					when "01101100100011101" => rgb <= "000000";
					when "01101100100011110" => rgb <= "000000";
					when "01101100100011111" => rgb <= "000000";
					when "01101100100100000" => rgb <= "000000";
					when "01101100100100001" => rgb <= "000000";
					when "01101100100100010" => rgb <= "000000";
					when "01101100100100011" => rgb <= "000000";
					when "01101100100100100" => rgb <= "000000";
					when "01101100100100101" => rgb <= "000000";
					when "01101100100100110" => rgb <= "000000";
					when "01101100100100111" => rgb <= "000000";
					when "01101100100101000" => rgb <= "000000";
					when "01101100100101001" => rgb <= "000000";
					when "01101100100101010" => rgb <= "000000";
					when "01101100100101011" => rgb <= "000000";
					when "01101100100101100" => rgb <= "000000";
					when "01101100100101101" => rgb <= "000000";
					when "01101100100101110" => rgb <= "000000";
					when "01101100100101111" => rgb <= "000000";
					when "01101100100110000" => rgb <= "000000";
					when "01101100100110001" => rgb <= "000000";
					when "01101100100110010" => rgb <= "000000";
					when "01101100100110011" => rgb <= "000000";
					when "01101100100110100" => rgb <= "000000";
					when "01101100100110101" => rgb <= "000000";
					when "01101100100110110" => rgb <= "000000";
					when "01101100100110111" => rgb <= "000000";
					when "01101100100111000" => rgb <= "000000";
					when "01101100100111001" => rgb <= "000000";
					when "01101100100111010" => rgb <= "000000";
					when "01101100100111011" => rgb <= "000000";
					when "01101100100111100" => rgb <= "000000";
					when "01101100100111101" => rgb <= "000000";
					when "01101100100111110" => rgb <= "000000";
					when "01101100100111111" => rgb <= "000000";
					when "01101101000000000" => rgb <= "000000";
					when "01101101000000001" => rgb <= "000000";
					when "01101101000000010" => rgb <= "000000";
					when "01101101000000011" => rgb <= "000000";
					when "01101101000000100" => rgb <= "000000";
					when "01101101000000101" => rgb <= "000000";
					when "01101101000000110" => rgb <= "000000";
					when "01101101000000111" => rgb <= "000000";
					when "01101101000001000" => rgb <= "000000";
					when "01101101000001001" => rgb <= "000000";
					when "01101101000001010" => rgb <= "000000";
					when "01101101000001011" => rgb <= "000000";
					when "01101101000001100" => rgb <= "000000";
					when "01101101000001101" => rgb <= "000000";
					when "01101101000001110" => rgb <= "000000";
					when "01101101000001111" => rgb <= "000000";
					when "01101101000010000" => rgb <= "000000";
					when "01101101000010001" => rgb <= "000000";
					when "01101101000010010" => rgb <= "000000";
					when "01101101000010011" => rgb <= "000000";
					when "01101101000010100" => rgb <= "000000";
					when "01101101000010101" => rgb <= "000000";
					when "01101101000010110" => rgb <= "000000";
					when "01101101000010111" => rgb <= "000000";
					when "01101101000011000" => rgb <= "000000";
					when "01101101000011001" => rgb <= "000000";
					when "01101101000011010" => rgb <= "000000";
					when "01101101000011011" => rgb <= "000000";
					when "01101101000011100" => rgb <= "000000";
					when "01101101000011101" => rgb <= "000000";
					when "01101101000011110" => rgb <= "000000";
					when "01101101000011111" => rgb <= "000000";
					when "01101101000100000" => rgb <= "000000";
					when "01101101000100001" => rgb <= "000000";
					when "01101101000100010" => rgb <= "000000";
					when "01101101000100011" => rgb <= "000000";
					when "01101101000100100" => rgb <= "000000";
					when "01101101000100101" => rgb <= "000000";
					when "01101101000100110" => rgb <= "000000";
					when "01101101000100111" => rgb <= "000000";
					when "01101101000101000" => rgb <= "000000";
					when "01101101000101001" => rgb <= "000000";
					when "01101101000101010" => rgb <= "000000";
					when "01101101000101011" => rgb <= "000000";
					when "01101101000101100" => rgb <= "000000";
					when "01101101000101101" => rgb <= "000000";
					when "01101101000101110" => rgb <= "000000";
					when "01101101000101111" => rgb <= "000000";
					when "01101101000110000" => rgb <= "000000";
					when "01101101000110001" => rgb <= "000000";
					when "01101101000110010" => rgb <= "000000";
					when "01101101000110011" => rgb <= "000000";
					when "01101101000110100" => rgb <= "000000";
					when "01101101000110101" => rgb <= "000000";
					when "01101101000110110" => rgb <= "000000";
					when "01101101000110111" => rgb <= "000000";
					when "01101101000111000" => rgb <= "000000";
					when "01101101000111001" => rgb <= "000000";
					when "01101101000111010" => rgb <= "000000";
					when "01101101000111011" => rgb <= "000000";
					when "01101101000111100" => rgb <= "000000";
					when "01101101000111101" => rgb <= "000000";
					when "01101101000111110" => rgb <= "000000";
					when "01101101000111111" => rgb <= "000000";
					when "01101101001000000" => rgb <= "000000";
					when "01101101001000001" => rgb <= "000000";
					when "01101101001000010" => rgb <= "000000";
					when "01101101001000011" => rgb <= "000000";
					when "01101101001000100" => rgb <= "000000";
					when "01101101001000101" => rgb <= "000000";
					when "01101101001000110" => rgb <= "000000";
					when "01101101001000111" => rgb <= "000000";
					when "01101101001001000" => rgb <= "000000";
					when "01101101001001001" => rgb <= "000000";
					when "01101101001001010" => rgb <= "000000";
					when "01101101001001011" => rgb <= "000000";
					when "01101101001001100" => rgb <= "000000";
					when "01101101001001101" => rgb <= "000000";
					when "01101101001001110" => rgb <= "000000";
					when "01101101001001111" => rgb <= "000000";
					when "01101101001010000" => rgb <= "000000";
					when "01101101001010001" => rgb <= "000000";
					when "01101101001010010" => rgb <= "000000";
					when "01101101001010011" => rgb <= "000000";
					when "01101101001010100" => rgb <= "000000";
					when "01101101001010101" => rgb <= "000000";
					when "01101101001010110" => rgb <= "000000";
					when "01101101001010111" => rgb <= "000000";
					when "01101101001011000" => rgb <= "000000";
					when "01101101001011001" => rgb <= "000000";
					when "01101101001011010" => rgb <= "000000";
					when "01101101001011011" => rgb <= "000000";
					when "01101101001011100" => rgb <= "000000";
					when "01101101001011101" => rgb <= "000000";
					when "01101101001011110" => rgb <= "000000";
					when "01101101001011111" => rgb <= "000000";
					when "01101101001100000" => rgb <= "000000";
					when "01101101001100001" => rgb <= "000000";
					when "01101101001100010" => rgb <= "000000";
					when "01101101001100011" => rgb <= "000000";
					when "01101101001100100" => rgb <= "000000";
					when "01101101001100101" => rgb <= "000000";
					when "01101101001100110" => rgb <= "000000";
					when "01101101001100111" => rgb <= "000000";
					when "01101101001101000" => rgb <= "000000";
					when "01101101001101001" => rgb <= "000000";
					when "01101101001101010" => rgb <= "000000";
					when "01101101001101011" => rgb <= "000000";
					when "01101101001101100" => rgb <= "000000";
					when "01101101001101101" => rgb <= "000000";
					when "01101101001101110" => rgb <= "000000";
					when "01101101001101111" => rgb <= "000000";
					when "01101101001110000" => rgb <= "000000";
					when "01101101001110001" => rgb <= "000000";
					when "01101101001110010" => rgb <= "000000";
					when "01101101001110011" => rgb <= "000000";
					when "01101101001110100" => rgb <= "000000";
					when "01101101001110101" => rgb <= "000000";
					when "01101101001110110" => rgb <= "000000";
					when "01101101001110111" => rgb <= "000000";
					when "01101101001111000" => rgb <= "000000";
					when "01101101001111001" => rgb <= "000000";
					when "01101101001111010" => rgb <= "000000";
					when "01101101001111011" => rgb <= "000000";
					when "01101101001111100" => rgb <= "000000";
					when "01101101001111101" => rgb <= "000000";
					when "01101101001111110" => rgb <= "000000";
					when "01101101001111111" => rgb <= "000000";
					when "01101101010000000" => rgb <= "000000";
					when "01101101010000001" => rgb <= "000000";
					when "01101101010000010" => rgb <= "000000";
					when "01101101010000011" => rgb <= "000000";
					when "01101101010000100" => rgb <= "000000";
					when "01101101010000101" => rgb <= "000000";
					when "01101101010000110" => rgb <= "000000";
					when "01101101010000111" => rgb <= "000000";
					when "01101101010001000" => rgb <= "010100";
					when "01101101010001001" => rgb <= "101000";
					when "01101101010001010" => rgb <= "101000";
					when "01101101010001011" => rgb <= "101000";
					when "01101101010001100" => rgb <= "101000";
					when "01101101010001101" => rgb <= "101000";
					when "01101101010001110" => rgb <= "101000";
					when "01101101010001111" => rgb <= "101000";
					when "01101101010010000" => rgb <= "101000";
					when "01101101010010001" => rgb <= "101000";
					when "01101101010010010" => rgb <= "101000";
					when "01101101010010011" => rgb <= "101000";
					when "01101101010010100" => rgb <= "101000";
					when "01101101010010101" => rgb <= "101000";
					when "01101101010010110" => rgb <= "101000";
					when "01101101010010111" => rgb <= "101000";
					when "01101101010011000" => rgb <= "101000";
					when "01101101010011001" => rgb <= "101000";
					when "01101101010011010" => rgb <= "101000";
					when "01101101010011011" => rgb <= "101000";
					when "01101101010011100" => rgb <= "101000";
					when "01101101010011101" => rgb <= "101000";
					when "01101101010011110" => rgb <= "101000";
					when "01101101010011111" => rgb <= "101000";
					when "01101101010100000" => rgb <= "101000";
					when "01101101010100001" => rgb <= "101000";
					when "01101101010100010" => rgb <= "101000";
					when "01101101010100011" => rgb <= "101000";
					when "01101101010100100" => rgb <= "101000";
					when "01101101010100101" => rgb <= "101000";
					when "01101101010100110" => rgb <= "101000";
					when "01101101010100111" => rgb <= "101000";
					when "01101101010101000" => rgb <= "101000";
					when "01101101010101001" => rgb <= "101000";
					when "01101101010101010" => rgb <= "101000";
					when "01101101010101011" => rgb <= "101000";
					when "01101101010101100" => rgb <= "101000";
					when "01101101010101101" => rgb <= "101000";
					when "01101101010101110" => rgb <= "101000";
					when "01101101010101111" => rgb <= "101000";
					when "01101101010110000" => rgb <= "101000";
					when "01101101010110001" => rgb <= "101000";
					when "01101101010110010" => rgb <= "101000";
					when "01101101010110011" => rgb <= "101000";
					when "01101101010110100" => rgb <= "101000";
					when "01101101010110101" => rgb <= "010100";
					when "01101101010110110" => rgb <= "000000";
					when "01101101010110111" => rgb <= "000000";
					when "01101101010111000" => rgb <= "000000";
					when "01101101010111001" => rgb <= "000000";
					when "01101101010111010" => rgb <= "000000";
					when "01101101010111011" => rgb <= "000000";
					when "01101101010111100" => rgb <= "000000";
					when "01101101010111101" => rgb <= "000000";
					when "01101101010111110" => rgb <= "000000";
					when "01101101010111111" => rgb <= "000000";
					when "01101101011000000" => rgb <= "000000";
					when "01101101011000001" => rgb <= "000000";
					when "01101101011000010" => rgb <= "000000";
					when "01101101011000011" => rgb <= "000000";
					when "01101101011000100" => rgb <= "000000";
					when "01101101011000101" => rgb <= "000000";
					when "01101101011000110" => rgb <= "000000";
					when "01101101011000111" => rgb <= "000000";
					when "01101101011001000" => rgb <= "000000";
					when "01101101011001001" => rgb <= "000000";
					when "01101101011001010" => rgb <= "000000";
					when "01101101011001011" => rgb <= "000000";
					when "01101101011001100" => rgb <= "000000";
					when "01101101011001101" => rgb <= "000000";
					when "01101101011001110" => rgb <= "000000";
					when "01101101011001111" => rgb <= "000000";
					when "01101101011010000" => rgb <= "000000";
					when "01101101011010001" => rgb <= "000000";
					when "01101101011010010" => rgb <= "000000";
					when "01101101011010011" => rgb <= "000000";
					when "01101101011010100" => rgb <= "000000";
					when "01101101011010101" => rgb <= "000000";
					when "01101101011010110" => rgb <= "000000";
					when "01101101011010111" => rgb <= "000000";
					when "01101101011011000" => rgb <= "000000";
					when "01101101011011001" => rgb <= "000000";
					when "01101101011011010" => rgb <= "000000";
					when "01101101011011011" => rgb <= "000000";
					when "01101101011011100" => rgb <= "000000";
					when "01101101011011101" => rgb <= "000000";
					when "01101101011011110" => rgb <= "000000";
					when "01101101011011111" => rgb <= "000000";
					when "01101101011100000" => rgb <= "000000";
					when "01101101011100001" => rgb <= "000000";
					when "01101101011100010" => rgb <= "000000";
					when "01101101011100011" => rgb <= "000000";
					when "01101101011100100" => rgb <= "000000";
					when "01101101011100101" => rgb <= "000000";
					when "01101101011100110" => rgb <= "000000";
					when "01101101011100111" => rgb <= "000000";
					when "01101101011101000" => rgb <= "000000";
					when "01101101011101001" => rgb <= "000000";
					when "01101101011101010" => rgb <= "000000";
					when "01101101011101011" => rgb <= "000000";
					when "01101101011101100" => rgb <= "000000";
					when "01101101011101101" => rgb <= "000000";
					when "01101101011101110" => rgb <= "000000";
					when "01101101011101111" => rgb <= "000000";
					when "01101101011110000" => rgb <= "000000";
					when "01101101011110001" => rgb <= "000000";
					when "01101101011110010" => rgb <= "000000";
					when "01101101011110011" => rgb <= "000000";
					when "01101101011110100" => rgb <= "000000";
					when "01101101011110101" => rgb <= "000000";
					when "01101101011110110" => rgb <= "000000";
					when "01101101011110111" => rgb <= "000000";
					when "01101101011111000" => rgb <= "000000";
					when "01101101011111001" => rgb <= "000000";
					when "01101101011111010" => rgb <= "000000";
					when "01101101011111011" => rgb <= "000000";
					when "01101101011111100" => rgb <= "000000";
					when "01101101011111101" => rgb <= "000000";
					when "01101101011111110" => rgb <= "000000";
					when "01101101011111111" => rgb <= "000000";
					when "01101101100000000" => rgb <= "000000";
					when "01101101100000001" => rgb <= "000000";
					when "01101101100000010" => rgb <= "000000";
					when "01101101100000011" => rgb <= "000000";
					when "01101101100000100" => rgb <= "000000";
					when "01101101100000101" => rgb <= "000000";
					when "01101101100000110" => rgb <= "000000";
					when "01101101100000111" => rgb <= "000000";
					when "01101101100001000" => rgb <= "000000";
					when "01101101100001001" => rgb <= "000000";
					when "01101101100001010" => rgb <= "000000";
					when "01101101100001011" => rgb <= "000000";
					when "01101101100001100" => rgb <= "000000";
					when "01101101100001101" => rgb <= "000000";
					when "01101101100001110" => rgb <= "000000";
					when "01101101100001111" => rgb <= "000000";
					when "01101101100010000" => rgb <= "000000";
					when "01101101100010001" => rgb <= "000000";
					when "01101101100010010" => rgb <= "000000";
					when "01101101100010011" => rgb <= "000000";
					when "01101101100010100" => rgb <= "000000";
					when "01101101100010101" => rgb <= "000000";
					when "01101101100010110" => rgb <= "000000";
					when "01101101100010111" => rgb <= "000000";
					when "01101101100011000" => rgb <= "000000";
					when "01101101100011001" => rgb <= "000000";
					when "01101101100011010" => rgb <= "000000";
					when "01101101100011011" => rgb <= "000000";
					when "01101101100011100" => rgb <= "000000";
					when "01101101100011101" => rgb <= "000000";
					when "01101101100011110" => rgb <= "000000";
					when "01101101100011111" => rgb <= "000000";
					when "01101101100100000" => rgb <= "000000";
					when "01101101100100001" => rgb <= "000000";
					when "01101101100100010" => rgb <= "000000";
					when "01101101100100011" => rgb <= "000000";
					when "01101101100100100" => rgb <= "000000";
					when "01101101100100101" => rgb <= "000000";
					when "01101101100100110" => rgb <= "000000";
					when "01101101100100111" => rgb <= "000000";
					when "01101101100101000" => rgb <= "000000";
					when "01101101100101001" => rgb <= "000000";
					when "01101101100101010" => rgb <= "000000";
					when "01101101100101011" => rgb <= "000000";
					when "01101101100101100" => rgb <= "000000";
					when "01101101100101101" => rgb <= "000000";
					when "01101101100101110" => rgb <= "000000";
					when "01101101100101111" => rgb <= "000000";
					when "01101101100110000" => rgb <= "000000";
					when "01101101100110001" => rgb <= "000000";
					when "01101101100110010" => rgb <= "000000";
					when "01101101100110011" => rgb <= "000000";
					when "01101101100110100" => rgb <= "000000";
					when "01101101100110101" => rgb <= "000000";
					when "01101101100110110" => rgb <= "000000";
					when "01101101100110111" => rgb <= "000000";
					when "01101101100111000" => rgb <= "000000";
					when "01101101100111001" => rgb <= "000000";
					when "01101101100111010" => rgb <= "000000";
					when "01101101100111011" => rgb <= "000000";
					when "01101101100111100" => rgb <= "000000";
					when "01101101100111101" => rgb <= "000000";
					when "01101101100111110" => rgb <= "000000";
					when "01101101100111111" => rgb <= "000000";
					when "01101110000000000" => rgb <= "000000";
					when "01101110000000001" => rgb <= "000000";
					when "01101110000000010" => rgb <= "000000";
					when "01101110000000011" => rgb <= "000000";
					when "01101110000000100" => rgb <= "000000";
					when "01101110000000101" => rgb <= "000000";
					when "01101110000000110" => rgb <= "000000";
					when "01101110000000111" => rgb <= "000000";
					when "01101110000001000" => rgb <= "000000";
					when "01101110000001001" => rgb <= "000000";
					when "01101110000001010" => rgb <= "000000";
					when "01101110000001011" => rgb <= "000000";
					when "01101110000001100" => rgb <= "000000";
					when "01101110000001101" => rgb <= "000000";
					when "01101110000001110" => rgb <= "000000";
					when "01101110000001111" => rgb <= "000000";
					when "01101110000010000" => rgb <= "000000";
					when "01101110000010001" => rgb <= "000000";
					when "01101110000010010" => rgb <= "000000";
					when "01101110000010011" => rgb <= "000000";
					when "01101110000010100" => rgb <= "000000";
					when "01101110000010101" => rgb <= "000000";
					when "01101110000010110" => rgb <= "000000";
					when "01101110000010111" => rgb <= "000000";
					when "01101110000011000" => rgb <= "000000";
					when "01101110000011001" => rgb <= "000000";
					when "01101110000011010" => rgb <= "000000";
					when "01101110000011011" => rgb <= "000000";
					when "01101110000011100" => rgb <= "000000";
					when "01101110000011101" => rgb <= "000000";
					when "01101110000011110" => rgb <= "000000";
					when "01101110000011111" => rgb <= "000000";
					when "01101110000100000" => rgb <= "000000";
					when "01101110000100001" => rgb <= "000000";
					when "01101110000100010" => rgb <= "000000";
					when "01101110000100011" => rgb <= "000000";
					when "01101110000100100" => rgb <= "000000";
					when "01101110000100101" => rgb <= "000000";
					when "01101110000100110" => rgb <= "000000";
					when "01101110000100111" => rgb <= "000000";
					when "01101110000101000" => rgb <= "000000";
					when "01101110000101001" => rgb <= "000000";
					when "01101110000101010" => rgb <= "000000";
					when "01101110000101011" => rgb <= "000000";
					when "01101110000101100" => rgb <= "000000";
					when "01101110000101101" => rgb <= "000000";
					when "01101110000101110" => rgb <= "000000";
					when "01101110000101111" => rgb <= "000000";
					when "01101110000110000" => rgb <= "000000";
					when "01101110000110001" => rgb <= "000000";
					when "01101110000110010" => rgb <= "000000";
					when "01101110000110011" => rgb <= "000000";
					when "01101110000110100" => rgb <= "000000";
					when "01101110000110101" => rgb <= "000000";
					when "01101110000110110" => rgb <= "000000";
					when "01101110000110111" => rgb <= "000000";
					when "01101110000111000" => rgb <= "000000";
					when "01101110000111001" => rgb <= "000000";
					when "01101110000111010" => rgb <= "000000";
					when "01101110000111011" => rgb <= "000000";
					when "01101110000111100" => rgb <= "000000";
					when "01101110000111101" => rgb <= "000000";
					when "01101110000111110" => rgb <= "000000";
					when "01101110000111111" => rgb <= "000000";
					when "01101110001000000" => rgb <= "000000";
					when "01101110001000001" => rgb <= "000000";
					when "01101110001000010" => rgb <= "000000";
					when "01101110001000011" => rgb <= "000000";
					when "01101110001000100" => rgb <= "000000";
					when "01101110001000101" => rgb <= "000000";
					when "01101110001000110" => rgb <= "000000";
					when "01101110001000111" => rgb <= "000000";
					when "01101110001001000" => rgb <= "000000";
					when "01101110001001001" => rgb <= "000000";
					when "01101110001001010" => rgb <= "000000";
					when "01101110001001011" => rgb <= "000000";
					when "01101110001001100" => rgb <= "000000";
					when "01101110001001101" => rgb <= "000000";
					when "01101110001001110" => rgb <= "000000";
					when "01101110001001111" => rgb <= "000000";
					when "01101110001010000" => rgb <= "000000";
					when "01101110001010001" => rgb <= "000000";
					when "01101110001010010" => rgb <= "000000";
					when "01101110001010011" => rgb <= "000000";
					when "01101110001010100" => rgb <= "000000";
					when "01101110001010101" => rgb <= "000000";
					when "01101110001010110" => rgb <= "000000";
					when "01101110001010111" => rgb <= "000000";
					when "01101110001011000" => rgb <= "000000";
					when "01101110001011001" => rgb <= "000000";
					when "01101110001011010" => rgb <= "000000";
					when "01101110001011011" => rgb <= "000000";
					when "01101110001011100" => rgb <= "000000";
					when "01101110001011101" => rgb <= "000000";
					when "01101110001011110" => rgb <= "000000";
					when "01101110001011111" => rgb <= "000000";
					when "01101110001100000" => rgb <= "000000";
					when "01101110001100001" => rgb <= "000000";
					when "01101110001100010" => rgb <= "000000";
					when "01101110001100011" => rgb <= "000000";
					when "01101110001100100" => rgb <= "000000";
					when "01101110001100101" => rgb <= "000000";
					when "01101110001100110" => rgb <= "000000";
					when "01101110001100111" => rgb <= "000000";
					when "01101110001101000" => rgb <= "000000";
					when "01101110001101001" => rgb <= "000000";
					when "01101110001101010" => rgb <= "000000";
					when "01101110001101011" => rgb <= "000000";
					when "01101110001101100" => rgb <= "000000";
					when "01101110001101101" => rgb <= "000000";
					when "01101110001101110" => rgb <= "000000";
					when "01101110001101111" => rgb <= "000000";
					when "01101110001110000" => rgb <= "000000";
					when "01101110001110001" => rgb <= "000000";
					when "01101110001110010" => rgb <= "000000";
					when "01101110001110011" => rgb <= "000000";
					when "01101110001110100" => rgb <= "000000";
					when "01101110001110101" => rgb <= "000000";
					when "01101110001110110" => rgb <= "000000";
					when "01101110001110111" => rgb <= "000000";
					when "01101110001111000" => rgb <= "000000";
					when "01101110001111001" => rgb <= "000000";
					when "01101110001111010" => rgb <= "000000";
					when "01101110001111011" => rgb <= "000000";
					when "01101110001111100" => rgb <= "000000";
					when "01101110001111101" => rgb <= "000000";
					when "01101110001111110" => rgb <= "000000";
					when "01101110001111111" => rgb <= "000000";
					when "01101110010000000" => rgb <= "000000";
					when "01101110010000001" => rgb <= "000000";
					when "01101110010000010" => rgb <= "000000";
					when "01101110010000011" => rgb <= "000000";
					when "01101110010000100" => rgb <= "000000";
					when "01101110010000101" => rgb <= "000000";
					when "01101110010000110" => rgb <= "000000";
					when "01101110010000111" => rgb <= "000000";
					when "01101110010001000" => rgb <= "010100";
					when "01101110010001001" => rgb <= "101000";
					when "01101110010001010" => rgb <= "101000";
					when "01101110010001011" => rgb <= "101000";
					when "01101110010001100" => rgb <= "101000";
					when "01101110010001101" => rgb <= "101000";
					when "01101110010001110" => rgb <= "101000";
					when "01101110010001111" => rgb <= "101000";
					when "01101110010010000" => rgb <= "101000";
					when "01101110010010001" => rgb <= "101000";
					when "01101110010010010" => rgb <= "101000";
					when "01101110010010011" => rgb <= "101000";
					when "01101110010010100" => rgb <= "101000";
					when "01101110010010101" => rgb <= "101000";
					when "01101110010010110" => rgb <= "101000";
					when "01101110010010111" => rgb <= "101000";
					when "01101110010011000" => rgb <= "101000";
					when "01101110010011001" => rgb <= "101000";
					when "01101110010011010" => rgb <= "101000";
					when "01101110010011011" => rgb <= "101000";
					when "01101110010011100" => rgb <= "101000";
					when "01101110010011101" => rgb <= "101000";
					when "01101110010011110" => rgb <= "101000";
					when "01101110010011111" => rgb <= "101000";
					when "01101110010100000" => rgb <= "101000";
					when "01101110010100001" => rgb <= "101000";
					when "01101110010100010" => rgb <= "101000";
					when "01101110010100011" => rgb <= "101000";
					when "01101110010100100" => rgb <= "101000";
					when "01101110010100101" => rgb <= "101000";
					when "01101110010100110" => rgb <= "101000";
					when "01101110010100111" => rgb <= "101000";
					when "01101110010101000" => rgb <= "101000";
					when "01101110010101001" => rgb <= "101000";
					when "01101110010101010" => rgb <= "101000";
					when "01101110010101011" => rgb <= "101000";
					when "01101110010101100" => rgb <= "101000";
					when "01101110010101101" => rgb <= "101000";
					when "01101110010101110" => rgb <= "101000";
					when "01101110010101111" => rgb <= "101000";
					when "01101110010110000" => rgb <= "101000";
					when "01101110010110001" => rgb <= "101000";
					when "01101110010110010" => rgb <= "101000";
					when "01101110010110011" => rgb <= "101000";
					when "01101110010110100" => rgb <= "101000";
					when "01101110010110101" => rgb <= "010100";
					when "01101110010110110" => rgb <= "000000";
					when "01101110010110111" => rgb <= "000000";
					when "01101110010111000" => rgb <= "000000";
					when "01101110010111001" => rgb <= "000000";
					when "01101110010111010" => rgb <= "000000";
					when "01101110010111011" => rgb <= "000000";
					when "01101110010111100" => rgb <= "000000";
					when "01101110010111101" => rgb <= "000000";
					when "01101110010111110" => rgb <= "000000";
					when "01101110010111111" => rgb <= "000000";
					when "01101110011000000" => rgb <= "000000";
					when "01101110011000001" => rgb <= "000000";
					when "01101110011000010" => rgb <= "000000";
					when "01101110011000011" => rgb <= "000000";
					when "01101110011000100" => rgb <= "000000";
					when "01101110011000101" => rgb <= "000000";
					when "01101110011000110" => rgb <= "000000";
					when "01101110011000111" => rgb <= "000000";
					when "01101110011001000" => rgb <= "000000";
					when "01101110011001001" => rgb <= "000000";
					when "01101110011001010" => rgb <= "000000";
					when "01101110011001011" => rgb <= "000000";
					when "01101110011001100" => rgb <= "000000";
					when "01101110011001101" => rgb <= "000000";
					when "01101110011001110" => rgb <= "000000";
					when "01101110011001111" => rgb <= "000000";
					when "01101110011010000" => rgb <= "000000";
					when "01101110011010001" => rgb <= "000000";
					when "01101110011010010" => rgb <= "000000";
					when "01101110011010011" => rgb <= "000000";
					when "01101110011010100" => rgb <= "000000";
					when "01101110011010101" => rgb <= "000000";
					when "01101110011010110" => rgb <= "000000";
					when "01101110011010111" => rgb <= "000000";
					when "01101110011011000" => rgb <= "000000";
					when "01101110011011001" => rgb <= "000000";
					when "01101110011011010" => rgb <= "000000";
					when "01101110011011011" => rgb <= "000000";
					when "01101110011011100" => rgb <= "000000";
					when "01101110011011101" => rgb <= "000000";
					when "01101110011011110" => rgb <= "000000";
					when "01101110011011111" => rgb <= "000000";
					when "01101110011100000" => rgb <= "000000";
					when "01101110011100001" => rgb <= "000000";
					when "01101110011100010" => rgb <= "000000";
					when "01101110011100011" => rgb <= "000000";
					when "01101110011100100" => rgb <= "000000";
					when "01101110011100101" => rgb <= "000000";
					when "01101110011100110" => rgb <= "000000";
					when "01101110011100111" => rgb <= "000000";
					when "01101110011101000" => rgb <= "000000";
					when "01101110011101001" => rgb <= "000000";
					when "01101110011101010" => rgb <= "000000";
					when "01101110011101011" => rgb <= "000000";
					when "01101110011101100" => rgb <= "000000";
					when "01101110011101101" => rgb <= "000000";
					when "01101110011101110" => rgb <= "000000";
					when "01101110011101111" => rgb <= "000000";
					when "01101110011110000" => rgb <= "000000";
					when "01101110011110001" => rgb <= "000000";
					when "01101110011110010" => rgb <= "000000";
					when "01101110011110011" => rgb <= "000000";
					when "01101110011110100" => rgb <= "000000";
					when "01101110011110101" => rgb <= "000000";
					when "01101110011110110" => rgb <= "000000";
					when "01101110011110111" => rgb <= "000000";
					when "01101110011111000" => rgb <= "000000";
					when "01101110011111001" => rgb <= "000000";
					when "01101110011111010" => rgb <= "000000";
					when "01101110011111011" => rgb <= "000000";
					when "01101110011111100" => rgb <= "000000";
					when "01101110011111101" => rgb <= "000000";
					when "01101110011111110" => rgb <= "000000";
					when "01101110011111111" => rgb <= "000000";
					when "01101110100000000" => rgb <= "000000";
					when "01101110100000001" => rgb <= "000000";
					when "01101110100000010" => rgb <= "000000";
					when "01101110100000011" => rgb <= "000000";
					when "01101110100000100" => rgb <= "000000";
					when "01101110100000101" => rgb <= "000000";
					when "01101110100000110" => rgb <= "000000";
					when "01101110100000111" => rgb <= "000000";
					when "01101110100001000" => rgb <= "000000";
					when "01101110100001001" => rgb <= "000000";
					when "01101110100001010" => rgb <= "000000";
					when "01101110100001011" => rgb <= "000000";
					when "01101110100001100" => rgb <= "000000";
					when "01101110100001101" => rgb <= "000000";
					when "01101110100001110" => rgb <= "000000";
					when "01101110100001111" => rgb <= "000000";
					when "01101110100010000" => rgb <= "000000";
					when "01101110100010001" => rgb <= "000000";
					when "01101110100010010" => rgb <= "000000";
					when "01101110100010011" => rgb <= "000000";
					when "01101110100010100" => rgb <= "000000";
					when "01101110100010101" => rgb <= "000000";
					when "01101110100010110" => rgb <= "000000";
					when "01101110100010111" => rgb <= "000000";
					when "01101110100011000" => rgb <= "000000";
					when "01101110100011001" => rgb <= "000000";
					when "01101110100011010" => rgb <= "000000";
					when "01101110100011011" => rgb <= "000000";
					when "01101110100011100" => rgb <= "000000";
					when "01101110100011101" => rgb <= "000000";
					when "01101110100011110" => rgb <= "000000";
					when "01101110100011111" => rgb <= "000000";
					when "01101110100100000" => rgb <= "000000";
					when "01101110100100001" => rgb <= "000000";
					when "01101110100100010" => rgb <= "000000";
					when "01101110100100011" => rgb <= "000000";
					when "01101110100100100" => rgb <= "000000";
					when "01101110100100101" => rgb <= "000000";
					when "01101110100100110" => rgb <= "000000";
					when "01101110100100111" => rgb <= "000000";
					when "01101110100101000" => rgb <= "000000";
					when "01101110100101001" => rgb <= "000000";
					when "01101110100101010" => rgb <= "000000";
					when "01101110100101011" => rgb <= "000000";
					when "01101110100101100" => rgb <= "000000";
					when "01101110100101101" => rgb <= "000000";
					when "01101110100101110" => rgb <= "000000";
					when "01101110100101111" => rgb <= "000000";
					when "01101110100110000" => rgb <= "000000";
					when "01101110100110001" => rgb <= "000000";
					when "01101110100110010" => rgb <= "000000";
					when "01101110100110011" => rgb <= "000000";
					when "01101110100110100" => rgb <= "000000";
					when "01101110100110101" => rgb <= "000000";
					when "01101110100110110" => rgb <= "000000";
					when "01101110100110111" => rgb <= "000000";
					when "01101110100111000" => rgb <= "000000";
					when "01101110100111001" => rgb <= "000000";
					when "01101110100111010" => rgb <= "000000";
					when "01101110100111011" => rgb <= "000000";
					when "01101110100111100" => rgb <= "000000";
					when "01101110100111101" => rgb <= "000000";
					when "01101110100111110" => rgb <= "000000";
					when "01101110100111111" => rgb <= "000000";
					when "01101111000000000" => rgb <= "000000";
					when "01101111000000001" => rgb <= "000000";
					when "01101111000000010" => rgb <= "000000";
					when "01101111000000011" => rgb <= "000000";
					when "01101111000000100" => rgb <= "000000";
					when "01101111000000101" => rgb <= "000000";
					when "01101111000000110" => rgb <= "000000";
					when "01101111000000111" => rgb <= "000000";
					when "01101111000001000" => rgb <= "000000";
					when "01101111000001001" => rgb <= "000000";
					when "01101111000001010" => rgb <= "000000";
					when "01101111000001011" => rgb <= "000000";
					when "01101111000001100" => rgb <= "000000";
					when "01101111000001101" => rgb <= "000000";
					when "01101111000001110" => rgb <= "000000";
					when "01101111000001111" => rgb <= "000000";
					when "01101111000010000" => rgb <= "000000";
					when "01101111000010001" => rgb <= "000000";
					when "01101111000010010" => rgb <= "000000";
					when "01101111000010011" => rgb <= "000000";
					when "01101111000010100" => rgb <= "000000";
					when "01101111000010101" => rgb <= "000000";
					when "01101111000010110" => rgb <= "000000";
					when "01101111000010111" => rgb <= "000000";
					when "01101111000011000" => rgb <= "000000";
					when "01101111000011001" => rgb <= "000000";
					when "01101111000011010" => rgb <= "000000";
					when "01101111000011011" => rgb <= "000000";
					when "01101111000011100" => rgb <= "000000";
					when "01101111000011101" => rgb <= "000000";
					when "01101111000011110" => rgb <= "000000";
					when "01101111000011111" => rgb <= "000000";
					when "01101111000100000" => rgb <= "000000";
					when "01101111000100001" => rgb <= "000000";
					when "01101111000100010" => rgb <= "000000";
					when "01101111000100011" => rgb <= "000000";
					when "01101111000100100" => rgb <= "000000";
					when "01101111000100101" => rgb <= "000000";
					when "01101111000100110" => rgb <= "000000";
					when "01101111000100111" => rgb <= "000000";
					when "01101111000101000" => rgb <= "000000";
					when "01101111000101001" => rgb <= "000000";
					when "01101111000101010" => rgb <= "000000";
					when "01101111000101011" => rgb <= "000000";
					when "01101111000101100" => rgb <= "000000";
					when "01101111000101101" => rgb <= "000000";
					when "01101111000101110" => rgb <= "000000";
					when "01101111000101111" => rgb <= "000000";
					when "01101111000110000" => rgb <= "000000";
					when "01101111000110001" => rgb <= "000000";
					when "01101111000110010" => rgb <= "000000";
					when "01101111000110011" => rgb <= "000000";
					when "01101111000110100" => rgb <= "000000";
					when "01101111000110101" => rgb <= "000000";
					when "01101111000110110" => rgb <= "000000";
					when "01101111000110111" => rgb <= "000000";
					when "01101111000111000" => rgb <= "000000";
					when "01101111000111001" => rgb <= "000000";
					when "01101111000111010" => rgb <= "000000";
					when "01101111000111011" => rgb <= "000000";
					when "01101111000111100" => rgb <= "000000";
					when "01101111000111101" => rgb <= "000000";
					when "01101111000111110" => rgb <= "000000";
					when "01101111000111111" => rgb <= "000000";
					when "01101111001000000" => rgb <= "000000";
					when "01101111001000001" => rgb <= "000000";
					when "01101111001000010" => rgb <= "000000";
					when "01101111001000011" => rgb <= "000000";
					when "01101111001000100" => rgb <= "000000";
					when "01101111001000101" => rgb <= "000000";
					when "01101111001000110" => rgb <= "000000";
					when "01101111001000111" => rgb <= "000000";
					when "01101111001001000" => rgb <= "000000";
					when "01101111001001001" => rgb <= "000000";
					when "01101111001001010" => rgb <= "000000";
					when "01101111001001011" => rgb <= "000000";
					when "01101111001001100" => rgb <= "000000";
					when "01101111001001101" => rgb <= "000000";
					when "01101111001001110" => rgb <= "000000";
					when "01101111001001111" => rgb <= "000000";
					when "01101111001010000" => rgb <= "000000";
					when "01101111001010001" => rgb <= "000000";
					when "01101111001010010" => rgb <= "000000";
					when "01101111001010011" => rgb <= "000000";
					when "01101111001010100" => rgb <= "000000";
					when "01101111001010101" => rgb <= "000000";
					when "01101111001010110" => rgb <= "000000";
					when "01101111001010111" => rgb <= "000000";
					when "01101111001011000" => rgb <= "000000";
					when "01101111001011001" => rgb <= "000000";
					when "01101111001011010" => rgb <= "000000";
					when "01101111001011011" => rgb <= "000000";
					when "01101111001011100" => rgb <= "000000";
					when "01101111001011101" => rgb <= "000000";
					when "01101111001011110" => rgb <= "000000";
					when "01101111001011111" => rgb <= "000000";
					when "01101111001100000" => rgb <= "000000";
					when "01101111001100001" => rgb <= "000000";
					when "01101111001100010" => rgb <= "000000";
					when "01101111001100011" => rgb <= "000000";
					when "01101111001100100" => rgb <= "000000";
					when "01101111001100101" => rgb <= "000000";
					when "01101111001100110" => rgb <= "000000";
					when "01101111001100111" => rgb <= "000000";
					when "01101111001101000" => rgb <= "000000";
					when "01101111001101001" => rgb <= "000000";
					when "01101111001101010" => rgb <= "000000";
					when "01101111001101011" => rgb <= "000000";
					when "01101111001101100" => rgb <= "000000";
					when "01101111001101101" => rgb <= "000000";
					when "01101111001101110" => rgb <= "000000";
					when "01101111001101111" => rgb <= "000000";
					when "01101111001110000" => rgb <= "000000";
					when "01101111001110001" => rgb <= "000000";
					when "01101111001110010" => rgb <= "000000";
					when "01101111001110011" => rgb <= "000000";
					when "01101111001110100" => rgb <= "000000";
					when "01101111001110101" => rgb <= "000000";
					when "01101111001110110" => rgb <= "000000";
					when "01101111001110111" => rgb <= "000000";
					when "01101111001111000" => rgb <= "000000";
					when "01101111001111001" => rgb <= "000000";
					when "01101111001111010" => rgb <= "000000";
					when "01101111001111011" => rgb <= "000000";
					when "01101111001111100" => rgb <= "000000";
					when "01101111001111101" => rgb <= "000000";
					when "01101111001111110" => rgb <= "000000";
					when "01101111001111111" => rgb <= "000000";
					when "01101111010000000" => rgb <= "000000";
					when "01101111010000001" => rgb <= "000000";
					when "01101111010000010" => rgb <= "000000";
					when "01101111010000011" => rgb <= "000000";
					when "01101111010000100" => rgb <= "000000";
					when "01101111010000101" => rgb <= "000000";
					when "01101111010000110" => rgb <= "000000";
					when "01101111010000111" => rgb <= "000000";
					when "01101111010001000" => rgb <= "010100";
					when "01101111010001001" => rgb <= "101000";
					when "01101111010001010" => rgb <= "101000";
					when "01101111010001011" => rgb <= "101000";
					when "01101111010001100" => rgb <= "101000";
					when "01101111010001101" => rgb <= "101000";
					when "01101111010001110" => rgb <= "101000";
					when "01101111010001111" => rgb <= "101000";
					when "01101111010010000" => rgb <= "101000";
					when "01101111010010001" => rgb <= "101000";
					when "01101111010010010" => rgb <= "101000";
					when "01101111010010011" => rgb <= "101000";
					when "01101111010010100" => rgb <= "101000";
					when "01101111010010101" => rgb <= "101000";
					when "01101111010010110" => rgb <= "101000";
					when "01101111010010111" => rgb <= "101000";
					when "01101111010011000" => rgb <= "101000";
					when "01101111010011001" => rgb <= "101000";
					when "01101111010011010" => rgb <= "101000";
					when "01101111010011011" => rgb <= "101000";
					when "01101111010011100" => rgb <= "101000";
					when "01101111010011101" => rgb <= "101000";
					when "01101111010011110" => rgb <= "101000";
					when "01101111010011111" => rgb <= "101000";
					when "01101111010100000" => rgb <= "101000";
					when "01101111010100001" => rgb <= "101000";
					when "01101111010100010" => rgb <= "101000";
					when "01101111010100011" => rgb <= "101000";
					when "01101111010100100" => rgb <= "101000";
					when "01101111010100101" => rgb <= "101000";
					when "01101111010100110" => rgb <= "101000";
					when "01101111010100111" => rgb <= "101000";
					when "01101111010101000" => rgb <= "101000";
					when "01101111010101001" => rgb <= "101000";
					when "01101111010101010" => rgb <= "101000";
					when "01101111010101011" => rgb <= "101000";
					when "01101111010101100" => rgb <= "101000";
					when "01101111010101101" => rgb <= "101000";
					when "01101111010101110" => rgb <= "101000";
					when "01101111010101111" => rgb <= "101000";
					when "01101111010110000" => rgb <= "101000";
					when "01101111010110001" => rgb <= "101000";
					when "01101111010110010" => rgb <= "101000";
					when "01101111010110011" => rgb <= "101000";
					when "01101111010110100" => rgb <= "101000";
					when "01101111010110101" => rgb <= "010100";
					when "01101111010110110" => rgb <= "000000";
					when "01101111010110111" => rgb <= "000000";
					when "01101111010111000" => rgb <= "000000";
					when "01101111010111001" => rgb <= "000000";
					when "01101111010111010" => rgb <= "000000";
					when "01101111010111011" => rgb <= "000000";
					when "01101111010111100" => rgb <= "000000";
					when "01101111010111101" => rgb <= "000000";
					when "01101111010111110" => rgb <= "000000";
					when "01101111010111111" => rgb <= "000000";
					when "01101111011000000" => rgb <= "000000";
					when "01101111011000001" => rgb <= "000000";
					when "01101111011000010" => rgb <= "000000";
					when "01101111011000011" => rgb <= "000000";
					when "01101111011000100" => rgb <= "000000";
					when "01101111011000101" => rgb <= "000000";
					when "01101111011000110" => rgb <= "000000";
					when "01101111011000111" => rgb <= "000000";
					when "01101111011001000" => rgb <= "000000";
					when "01101111011001001" => rgb <= "000000";
					when "01101111011001010" => rgb <= "000000";
					when "01101111011001011" => rgb <= "000000";
					when "01101111011001100" => rgb <= "000000";
					when "01101111011001101" => rgb <= "000000";
					when "01101111011001110" => rgb <= "000000";
					when "01101111011001111" => rgb <= "000000";
					when "01101111011010000" => rgb <= "000000";
					when "01101111011010001" => rgb <= "000000";
					when "01101111011010010" => rgb <= "000000";
					when "01101111011010011" => rgb <= "000000";
					when "01101111011010100" => rgb <= "000000";
					when "01101111011010101" => rgb <= "000000";
					when "01101111011010110" => rgb <= "000000";
					when "01101111011010111" => rgb <= "000000";
					when "01101111011011000" => rgb <= "000000";
					when "01101111011011001" => rgb <= "000000";
					when "01101111011011010" => rgb <= "000000";
					when "01101111011011011" => rgb <= "000000";
					when "01101111011011100" => rgb <= "000000";
					when "01101111011011101" => rgb <= "000000";
					when "01101111011011110" => rgb <= "000000";
					when "01101111011011111" => rgb <= "000000";
					when "01101111011100000" => rgb <= "000000";
					when "01101111011100001" => rgb <= "000000";
					when "01101111011100010" => rgb <= "000000";
					when "01101111011100011" => rgb <= "000000";
					when "01101111011100100" => rgb <= "000000";
					when "01101111011100101" => rgb <= "000000";
					when "01101111011100110" => rgb <= "000000";
					when "01101111011100111" => rgb <= "000000";
					when "01101111011101000" => rgb <= "000000";
					when "01101111011101001" => rgb <= "000000";
					when "01101111011101010" => rgb <= "000000";
					when "01101111011101011" => rgb <= "000000";
					when "01101111011101100" => rgb <= "000000";
					when "01101111011101101" => rgb <= "000000";
					when "01101111011101110" => rgb <= "000000";
					when "01101111011101111" => rgb <= "000000";
					when "01101111011110000" => rgb <= "000000";
					when "01101111011110001" => rgb <= "000000";
					when "01101111011110010" => rgb <= "000000";
					when "01101111011110011" => rgb <= "000000";
					when "01101111011110100" => rgb <= "000000";
					when "01101111011110101" => rgb <= "000000";
					when "01101111011110110" => rgb <= "000000";
					when "01101111011110111" => rgb <= "000000";
					when "01101111011111000" => rgb <= "000000";
					when "01101111011111001" => rgb <= "000000";
					when "01101111011111010" => rgb <= "000000";
					when "01101111011111011" => rgb <= "000000";
					when "01101111011111100" => rgb <= "000000";
					when "01101111011111101" => rgb <= "000000";
					when "01101111011111110" => rgb <= "000000";
					when "01101111011111111" => rgb <= "000000";
					when "01101111100000000" => rgb <= "000000";
					when "01101111100000001" => rgb <= "000000";
					when "01101111100000010" => rgb <= "000000";
					when "01101111100000011" => rgb <= "000000";
					when "01101111100000100" => rgb <= "000000";
					when "01101111100000101" => rgb <= "000000";
					when "01101111100000110" => rgb <= "000000";
					when "01101111100000111" => rgb <= "000000";
					when "01101111100001000" => rgb <= "000000";
					when "01101111100001001" => rgb <= "000000";
					when "01101111100001010" => rgb <= "000000";
					when "01101111100001011" => rgb <= "000000";
					when "01101111100001100" => rgb <= "000000";
					when "01101111100001101" => rgb <= "000000";
					when "01101111100001110" => rgb <= "000000";
					when "01101111100001111" => rgb <= "000000";
					when "01101111100010000" => rgb <= "000000";
					when "01101111100010001" => rgb <= "000000";
					when "01101111100010010" => rgb <= "000000";
					when "01101111100010011" => rgb <= "000000";
					when "01101111100010100" => rgb <= "000000";
					when "01101111100010101" => rgb <= "000000";
					when "01101111100010110" => rgb <= "000000";
					when "01101111100010111" => rgb <= "000000";
					when "01101111100011000" => rgb <= "000000";
					when "01101111100011001" => rgb <= "000000";
					when "01101111100011010" => rgb <= "000000";
					when "01101111100011011" => rgb <= "000000";
					when "01101111100011100" => rgb <= "000000";
					when "01101111100011101" => rgb <= "000000";
					when "01101111100011110" => rgb <= "000000";
					when "01101111100011111" => rgb <= "000000";
					when "01101111100100000" => rgb <= "000000";
					when "01101111100100001" => rgb <= "000000";
					when "01101111100100010" => rgb <= "000000";
					when "01101111100100011" => rgb <= "000000";
					when "01101111100100100" => rgb <= "000000";
					when "01101111100100101" => rgb <= "000000";
					when "01101111100100110" => rgb <= "000000";
					when "01101111100100111" => rgb <= "000000";
					when "01101111100101000" => rgb <= "000000";
					when "01101111100101001" => rgb <= "000000";
					when "01101111100101010" => rgb <= "000000";
					when "01101111100101011" => rgb <= "000000";
					when "01101111100101100" => rgb <= "000000";
					when "01101111100101101" => rgb <= "000000";
					when "01101111100101110" => rgb <= "000000";
					when "01101111100101111" => rgb <= "000000";
					when "01101111100110000" => rgb <= "000000";
					when "01101111100110001" => rgb <= "000000";
					when "01101111100110010" => rgb <= "000000";
					when "01101111100110011" => rgb <= "000000";
					when "01101111100110100" => rgb <= "000000";
					when "01101111100110101" => rgb <= "000000";
					when "01101111100110110" => rgb <= "000000";
					when "01101111100110111" => rgb <= "000000";
					when "01101111100111000" => rgb <= "000000";
					when "01101111100111001" => rgb <= "000000";
					when "01101111100111010" => rgb <= "000000";
					when "01101111100111011" => rgb <= "000000";
					when "01101111100111100" => rgb <= "000000";
					when "01101111100111101" => rgb <= "000000";
					when "01101111100111110" => rgb <= "000000";
					when "01101111100111111" => rgb <= "000000";
					when "01110000000000000" => rgb <= "000000";
					when "01110000000000001" => rgb <= "000000";
					when "01110000000000010" => rgb <= "000000";
					when "01110000000000011" => rgb <= "000000";
					when "01110000000000100" => rgb <= "000000";
					when "01110000000000101" => rgb <= "000000";
					when "01110000000000110" => rgb <= "000000";
					when "01110000000000111" => rgb <= "000000";
					when "01110000000001000" => rgb <= "000000";
					when "01110000000001001" => rgb <= "000000";
					when "01110000000001010" => rgb <= "000000";
					when "01110000000001011" => rgb <= "000000";
					when "01110000000001100" => rgb <= "000000";
					when "01110000000001101" => rgb <= "000000";
					when "01110000000001110" => rgb <= "000000";
					when "01110000000001111" => rgb <= "000000";
					when "01110000000010000" => rgb <= "000000";
					when "01110000000010001" => rgb <= "000000";
					when "01110000000010010" => rgb <= "000000";
					when "01110000000010011" => rgb <= "000000";
					when "01110000000010100" => rgb <= "000000";
					when "01110000000010101" => rgb <= "000000";
					when "01110000000010110" => rgb <= "000000";
					when "01110000000010111" => rgb <= "000000";
					when "01110000000011000" => rgb <= "000000";
					when "01110000000011001" => rgb <= "000000";
					when "01110000000011010" => rgb <= "000000";
					when "01110000000011011" => rgb <= "000000";
					when "01110000000011100" => rgb <= "000000";
					when "01110000000011101" => rgb <= "000000";
					when "01110000000011110" => rgb <= "000000";
					when "01110000000011111" => rgb <= "000000";
					when "01110000000100000" => rgb <= "000000";
					when "01110000000100001" => rgb <= "000000";
					when "01110000000100010" => rgb <= "000000";
					when "01110000000100011" => rgb <= "000000";
					when "01110000000100100" => rgb <= "000000";
					when "01110000000100101" => rgb <= "000000";
					when "01110000000100110" => rgb <= "000000";
					when "01110000000100111" => rgb <= "000000";
					when "01110000000101000" => rgb <= "000000";
					when "01110000000101001" => rgb <= "000000";
					when "01110000000101010" => rgb <= "000000";
					when "01110000000101011" => rgb <= "000000";
					when "01110000000101100" => rgb <= "000000";
					when "01110000000101101" => rgb <= "000000";
					when "01110000000101110" => rgb <= "000000";
					when "01110000000101111" => rgb <= "000000";
					when "01110000000110000" => rgb <= "000000";
					when "01110000000110001" => rgb <= "000000";
					when "01110000000110010" => rgb <= "000000";
					when "01110000000110011" => rgb <= "000000";
					when "01110000000110100" => rgb <= "000000";
					when "01110000000110101" => rgb <= "000000";
					when "01110000000110110" => rgb <= "000000";
					when "01110000000110111" => rgb <= "000000";
					when "01110000000111000" => rgb <= "000000";
					when "01110000000111001" => rgb <= "000000";
					when "01110000000111010" => rgb <= "000000";
					when "01110000000111011" => rgb <= "000000";
					when "01110000000111100" => rgb <= "000000";
					when "01110000000111101" => rgb <= "000000";
					when "01110000000111110" => rgb <= "000000";
					when "01110000000111111" => rgb <= "000000";
					when "01110000001000000" => rgb <= "000000";
					when "01110000001000001" => rgb <= "000000";
					when "01110000001000010" => rgb <= "000000";
					when "01110000001000011" => rgb <= "000000";
					when "01110000001000100" => rgb <= "000000";
					when "01110000001000101" => rgb <= "000000";
					when "01110000001000110" => rgb <= "000000";
					when "01110000001000111" => rgb <= "000000";
					when "01110000001001000" => rgb <= "000000";
					when "01110000001001001" => rgb <= "000000";
					when "01110000001001010" => rgb <= "000000";
					when "01110000001001011" => rgb <= "000000";
					when "01110000001001100" => rgb <= "000000";
					when "01110000001001101" => rgb <= "000000";
					when "01110000001001110" => rgb <= "000000";
					when "01110000001001111" => rgb <= "000000";
					when "01110000001010000" => rgb <= "000000";
					when "01110000001010001" => rgb <= "000000";
					when "01110000001010010" => rgb <= "000000";
					when "01110000001010011" => rgb <= "000000";
					when "01110000001010100" => rgb <= "000000";
					when "01110000001010101" => rgb <= "000000";
					when "01110000001010110" => rgb <= "000000";
					when "01110000001010111" => rgb <= "000000";
					when "01110000001011000" => rgb <= "000000";
					when "01110000001011001" => rgb <= "000000";
					when "01110000001011010" => rgb <= "000000";
					when "01110000001011011" => rgb <= "000000";
					when "01110000001011100" => rgb <= "000000";
					when "01110000001011101" => rgb <= "000000";
					when "01110000001011110" => rgb <= "000000";
					when "01110000001011111" => rgb <= "000000";
					when "01110000001100000" => rgb <= "000000";
					when "01110000001100001" => rgb <= "000000";
					when "01110000001100010" => rgb <= "000000";
					when "01110000001100011" => rgb <= "000000";
					when "01110000001100100" => rgb <= "000000";
					when "01110000001100101" => rgb <= "000000";
					when "01110000001100110" => rgb <= "000000";
					when "01110000001100111" => rgb <= "000000";
					when "01110000001101000" => rgb <= "000000";
					when "01110000001101001" => rgb <= "000000";
					when "01110000001101010" => rgb <= "000000";
					when "01110000001101011" => rgb <= "000000";
					when "01110000001101100" => rgb <= "000000";
					when "01110000001101101" => rgb <= "000000";
					when "01110000001101110" => rgb <= "000000";
					when "01110000001101111" => rgb <= "000000";
					when "01110000001110000" => rgb <= "000000";
					when "01110000001110001" => rgb <= "000000";
					when "01110000001110010" => rgb <= "000000";
					when "01110000001110011" => rgb <= "000000";
					when "01110000001110100" => rgb <= "000000";
					when "01110000001110101" => rgb <= "000000";
					when "01110000001110110" => rgb <= "000000";
					when "01110000001110111" => rgb <= "000000";
					when "01110000001111000" => rgb <= "000000";
					when "01110000001111001" => rgb <= "000000";
					when "01110000001111010" => rgb <= "000000";
					when "01110000001111011" => rgb <= "000000";
					when "01110000001111100" => rgb <= "000000";
					when "01110000001111101" => rgb <= "000000";
					when "01110000001111110" => rgb <= "000000";
					when "01110000001111111" => rgb <= "000000";
					when "01110000010000000" => rgb <= "000000";
					when "01110000010000001" => rgb <= "000000";
					when "01110000010000010" => rgb <= "000000";
					when "01110000010000011" => rgb <= "000000";
					when "01110000010000100" => rgb <= "000000";
					when "01110000010000101" => rgb <= "000000";
					when "01110000010000110" => rgb <= "000000";
					when "01110000010000111" => rgb <= "000000";
					when "01110000010001000" => rgb <= "010100";
					when "01110000010001001" => rgb <= "101000";
					when "01110000010001010" => rgb <= "101000";
					when "01110000010001011" => rgb <= "101000";
					when "01110000010001100" => rgb <= "101000";
					when "01110000010001101" => rgb <= "101000";
					when "01110000010001110" => rgb <= "101000";
					when "01110000010001111" => rgb <= "101000";
					when "01110000010010000" => rgb <= "101000";
					when "01110000010010001" => rgb <= "101000";
					when "01110000010010010" => rgb <= "101000";
					when "01110000010010011" => rgb <= "101000";
					when "01110000010010100" => rgb <= "101000";
					when "01110000010010101" => rgb <= "101000";
					when "01110000010010110" => rgb <= "101000";
					when "01110000010010111" => rgb <= "101000";
					when "01110000010011000" => rgb <= "101000";
					when "01110000010011001" => rgb <= "101000";
					when "01110000010011010" => rgb <= "101000";
					when "01110000010011011" => rgb <= "101000";
					when "01110000010011100" => rgb <= "101000";
					when "01110000010011101" => rgb <= "101000";
					when "01110000010011110" => rgb <= "101000";
					when "01110000010011111" => rgb <= "101000";
					when "01110000010100000" => rgb <= "101000";
					when "01110000010100001" => rgb <= "101000";
					when "01110000010100010" => rgb <= "101000";
					when "01110000010100011" => rgb <= "101000";
					when "01110000010100100" => rgb <= "101000";
					when "01110000010100101" => rgb <= "101000";
					when "01110000010100110" => rgb <= "101000";
					when "01110000010100111" => rgb <= "101000";
					when "01110000010101000" => rgb <= "101000";
					when "01110000010101001" => rgb <= "101000";
					when "01110000010101010" => rgb <= "101000";
					when "01110000010101011" => rgb <= "101000";
					when "01110000010101100" => rgb <= "101000";
					when "01110000010101101" => rgb <= "101000";
					when "01110000010101110" => rgb <= "101000";
					when "01110000010101111" => rgb <= "101000";
					when "01110000010110000" => rgb <= "101000";
					when "01110000010110001" => rgb <= "101000";
					when "01110000010110010" => rgb <= "101000";
					when "01110000010110011" => rgb <= "101000";
					when "01110000010110100" => rgb <= "101000";
					when "01110000010110101" => rgb <= "010100";
					when "01110000010110110" => rgb <= "000000";
					when "01110000010110111" => rgb <= "000000";
					when "01110000010111000" => rgb <= "000000";
					when "01110000010111001" => rgb <= "000000";
					when "01110000010111010" => rgb <= "000000";
					when "01110000010111011" => rgb <= "000000";
					when "01110000010111100" => rgb <= "000000";
					when "01110000010111101" => rgb <= "000000";
					when "01110000010111110" => rgb <= "000000";
					when "01110000010111111" => rgb <= "000000";
					when "01110000011000000" => rgb <= "000000";
					when "01110000011000001" => rgb <= "000000";
					when "01110000011000010" => rgb <= "000000";
					when "01110000011000011" => rgb <= "000000";
					when "01110000011000100" => rgb <= "000000";
					when "01110000011000101" => rgb <= "000000";
					when "01110000011000110" => rgb <= "000000";
					when "01110000011000111" => rgb <= "000000";
					when "01110000011001000" => rgb <= "000000";
					when "01110000011001001" => rgb <= "000000";
					when "01110000011001010" => rgb <= "000000";
					when "01110000011001011" => rgb <= "000000";
					when "01110000011001100" => rgb <= "000000";
					when "01110000011001101" => rgb <= "000000";
					when "01110000011001110" => rgb <= "000000";
					when "01110000011001111" => rgb <= "000000";
					when "01110000011010000" => rgb <= "000000";
					when "01110000011010001" => rgb <= "000000";
					when "01110000011010010" => rgb <= "000000";
					when "01110000011010011" => rgb <= "000000";
					when "01110000011010100" => rgb <= "000000";
					when "01110000011010101" => rgb <= "000000";
					when "01110000011010110" => rgb <= "000000";
					when "01110000011010111" => rgb <= "000000";
					when "01110000011011000" => rgb <= "000000";
					when "01110000011011001" => rgb <= "000000";
					when "01110000011011010" => rgb <= "000000";
					when "01110000011011011" => rgb <= "000000";
					when "01110000011011100" => rgb <= "000000";
					when "01110000011011101" => rgb <= "000000";
					when "01110000011011110" => rgb <= "000000";
					when "01110000011011111" => rgb <= "000000";
					when "01110000011100000" => rgb <= "000000";
					when "01110000011100001" => rgb <= "000000";
					when "01110000011100010" => rgb <= "000000";
					when "01110000011100011" => rgb <= "000000";
					when "01110000011100100" => rgb <= "000000";
					when "01110000011100101" => rgb <= "000000";
					when "01110000011100110" => rgb <= "000000";
					when "01110000011100111" => rgb <= "000000";
					when "01110000011101000" => rgb <= "000000";
					when "01110000011101001" => rgb <= "000000";
					when "01110000011101010" => rgb <= "000000";
					when "01110000011101011" => rgb <= "000000";
					when "01110000011101100" => rgb <= "000000";
					when "01110000011101101" => rgb <= "000000";
					when "01110000011101110" => rgb <= "000000";
					when "01110000011101111" => rgb <= "000000";
					when "01110000011110000" => rgb <= "000000";
					when "01110000011110001" => rgb <= "000000";
					when "01110000011110010" => rgb <= "000000";
					when "01110000011110011" => rgb <= "000000";
					when "01110000011110100" => rgb <= "000000";
					when "01110000011110101" => rgb <= "000000";
					when "01110000011110110" => rgb <= "000000";
					when "01110000011110111" => rgb <= "000000";
					when "01110000011111000" => rgb <= "000000";
					when "01110000011111001" => rgb <= "000000";
					when "01110000011111010" => rgb <= "000000";
					when "01110000011111011" => rgb <= "000000";
					when "01110000011111100" => rgb <= "000000";
					when "01110000011111101" => rgb <= "000000";
					when "01110000011111110" => rgb <= "000000";
					when "01110000011111111" => rgb <= "000000";
					when "01110000100000000" => rgb <= "000000";
					when "01110000100000001" => rgb <= "000000";
					when "01110000100000010" => rgb <= "000000";
					when "01110000100000011" => rgb <= "000000";
					when "01110000100000100" => rgb <= "000000";
					when "01110000100000101" => rgb <= "000000";
					when "01110000100000110" => rgb <= "000000";
					when "01110000100000111" => rgb <= "000000";
					when "01110000100001000" => rgb <= "000000";
					when "01110000100001001" => rgb <= "000000";
					when "01110000100001010" => rgb <= "000000";
					when "01110000100001011" => rgb <= "000000";
					when "01110000100001100" => rgb <= "000000";
					when "01110000100001101" => rgb <= "000000";
					when "01110000100001110" => rgb <= "000000";
					when "01110000100001111" => rgb <= "000000";
					when "01110000100010000" => rgb <= "000000";
					when "01110000100010001" => rgb <= "000000";
					when "01110000100010010" => rgb <= "000000";
					when "01110000100010011" => rgb <= "000000";
					when "01110000100010100" => rgb <= "000000";
					when "01110000100010101" => rgb <= "000000";
					when "01110000100010110" => rgb <= "000000";
					when "01110000100010111" => rgb <= "000000";
					when "01110000100011000" => rgb <= "000000";
					when "01110000100011001" => rgb <= "000000";
					when "01110000100011010" => rgb <= "000000";
					when "01110000100011011" => rgb <= "000000";
					when "01110000100011100" => rgb <= "000000";
					when "01110000100011101" => rgb <= "000000";
					when "01110000100011110" => rgb <= "000000";
					when "01110000100011111" => rgb <= "000000";
					when "01110000100100000" => rgb <= "000000";
					when "01110000100100001" => rgb <= "000000";
					when "01110000100100010" => rgb <= "000000";
					when "01110000100100011" => rgb <= "000000";
					when "01110000100100100" => rgb <= "000000";
					when "01110000100100101" => rgb <= "000000";
					when "01110000100100110" => rgb <= "000000";
					when "01110000100100111" => rgb <= "000000";
					when "01110000100101000" => rgb <= "000000";
					when "01110000100101001" => rgb <= "000000";
					when "01110000100101010" => rgb <= "000000";
					when "01110000100101011" => rgb <= "000000";
					when "01110000100101100" => rgb <= "000000";
					when "01110000100101101" => rgb <= "000000";
					when "01110000100101110" => rgb <= "000000";
					when "01110000100101111" => rgb <= "000000";
					when "01110000100110000" => rgb <= "000000";
					when "01110000100110001" => rgb <= "000000";
					when "01110000100110010" => rgb <= "000000";
					when "01110000100110011" => rgb <= "000000";
					when "01110000100110100" => rgb <= "000000";
					when "01110000100110101" => rgb <= "000000";
					when "01110000100110110" => rgb <= "000000";
					when "01110000100110111" => rgb <= "000000";
					when "01110000100111000" => rgb <= "000000";
					when "01110000100111001" => rgb <= "000000";
					when "01110000100111010" => rgb <= "000000";
					when "01110000100111011" => rgb <= "000000";
					when "01110000100111100" => rgb <= "000000";
					when "01110000100111101" => rgb <= "000000";
					when "01110000100111110" => rgb <= "000000";
					when "01110000100111111" => rgb <= "000000";
					when "01110001000000000" => rgb <= "000000";
					when "01110001000000001" => rgb <= "000000";
					when "01110001000000010" => rgb <= "000000";
					when "01110001000000011" => rgb <= "000000";
					when "01110001000000100" => rgb <= "000000";
					when "01110001000000101" => rgb <= "000000";
					when "01110001000000110" => rgb <= "000000";
					when "01110001000000111" => rgb <= "000000";
					when "01110001000001000" => rgb <= "000000";
					when "01110001000001001" => rgb <= "000000";
					when "01110001000001010" => rgb <= "000000";
					when "01110001000001011" => rgb <= "000000";
					when "01110001000001100" => rgb <= "000000";
					when "01110001000001101" => rgb <= "000000";
					when "01110001000001110" => rgb <= "000000";
					when "01110001000001111" => rgb <= "000000";
					when "01110001000010000" => rgb <= "000000";
					when "01110001000010001" => rgb <= "000000";
					when "01110001000010010" => rgb <= "000000";
					when "01110001000010011" => rgb <= "000000";
					when "01110001000010100" => rgb <= "000000";
					when "01110001000010101" => rgb <= "000000";
					when "01110001000010110" => rgb <= "000000";
					when "01110001000010111" => rgb <= "000000";
					when "01110001000011000" => rgb <= "000000";
					when "01110001000011001" => rgb <= "000000";
					when "01110001000011010" => rgb <= "000000";
					when "01110001000011011" => rgb <= "000000";
					when "01110001000011100" => rgb <= "000000";
					when "01110001000011101" => rgb <= "000000";
					when "01110001000011110" => rgb <= "000000";
					when "01110001000011111" => rgb <= "000000";
					when "01110001000100000" => rgb <= "000000";
					when "01110001000100001" => rgb <= "000000";
					when "01110001000100010" => rgb <= "000000";
					when "01110001000100011" => rgb <= "000000";
					when "01110001000100100" => rgb <= "000000";
					when "01110001000100101" => rgb <= "000000";
					when "01110001000100110" => rgb <= "000000";
					when "01110001000100111" => rgb <= "000000";
					when "01110001000101000" => rgb <= "000000";
					when "01110001000101001" => rgb <= "000000";
					when "01110001000101010" => rgb <= "000000";
					when "01110001000101011" => rgb <= "000000";
					when "01110001000101100" => rgb <= "000000";
					when "01110001000101101" => rgb <= "000000";
					when "01110001000101110" => rgb <= "000000";
					when "01110001000101111" => rgb <= "000000";
					when "01110001000110000" => rgb <= "000000";
					when "01110001000110001" => rgb <= "000000";
					when "01110001000110010" => rgb <= "000000";
					when "01110001000110011" => rgb <= "000000";
					when "01110001000110100" => rgb <= "000000";
					when "01110001000110101" => rgb <= "000000";
					when "01110001000110110" => rgb <= "000000";
					when "01110001000110111" => rgb <= "000000";
					when "01110001000111000" => rgb <= "000000";
					when "01110001000111001" => rgb <= "000000";
					when "01110001000111010" => rgb <= "000000";
					when "01110001000111011" => rgb <= "000000";
					when "01110001000111100" => rgb <= "000000";
					when "01110001000111101" => rgb <= "000000";
					when "01110001000111110" => rgb <= "000000";
					when "01110001000111111" => rgb <= "000000";
					when "01110001001000000" => rgb <= "000000";
					when "01110001001000001" => rgb <= "000000";
					when "01110001001000010" => rgb <= "000000";
					when "01110001001000011" => rgb <= "000000";
					when "01110001001000100" => rgb <= "000000";
					when "01110001001000101" => rgb <= "000000";
					when "01110001001000110" => rgb <= "000000";
					when "01110001001000111" => rgb <= "000000";
					when "01110001001001000" => rgb <= "000000";
					when "01110001001001001" => rgb <= "000000";
					when "01110001001001010" => rgb <= "000000";
					when "01110001001001011" => rgb <= "000000";
					when "01110001001001100" => rgb <= "000000";
					when "01110001001001101" => rgb <= "000000";
					when "01110001001001110" => rgb <= "000000";
					when "01110001001001111" => rgb <= "000000";
					when "01110001001010000" => rgb <= "000000";
					when "01110001001010001" => rgb <= "000000";
					when "01110001001010010" => rgb <= "000000";
					when "01110001001010011" => rgb <= "000000";
					when "01110001001010100" => rgb <= "000000";
					when "01110001001010101" => rgb <= "000000";
					when "01110001001010110" => rgb <= "000000";
					when "01110001001010111" => rgb <= "000000";
					when "01110001001011000" => rgb <= "000000";
					when "01110001001011001" => rgb <= "000000";
					when "01110001001011010" => rgb <= "000000";
					when "01110001001011011" => rgb <= "000000";
					when "01110001001011100" => rgb <= "000000";
					when "01110001001011101" => rgb <= "000000";
					when "01110001001011110" => rgb <= "000000";
					when "01110001001011111" => rgb <= "000000";
					when "01110001001100000" => rgb <= "000000";
					when "01110001001100001" => rgb <= "000000";
					when "01110001001100010" => rgb <= "000000";
					when "01110001001100011" => rgb <= "000000";
					when "01110001001100100" => rgb <= "000000";
					when "01110001001100101" => rgb <= "000000";
					when "01110001001100110" => rgb <= "000000";
					when "01110001001100111" => rgb <= "000000";
					when "01110001001101000" => rgb <= "000000";
					when "01110001001101001" => rgb <= "000000";
					when "01110001001101010" => rgb <= "000000";
					when "01110001001101011" => rgb <= "000000";
					when "01110001001101100" => rgb <= "000000";
					when "01110001001101101" => rgb <= "000000";
					when "01110001001101110" => rgb <= "000000";
					when "01110001001101111" => rgb <= "000000";
					when "01110001001110000" => rgb <= "000000";
					when "01110001001110001" => rgb <= "000000";
					when "01110001001110010" => rgb <= "000000";
					when "01110001001110011" => rgb <= "000000";
					when "01110001001110100" => rgb <= "000000";
					when "01110001001110101" => rgb <= "000000";
					when "01110001001110110" => rgb <= "000000";
					when "01110001001110111" => rgb <= "000000";
					when "01110001001111000" => rgb <= "000000";
					when "01110001001111001" => rgb <= "000000";
					when "01110001001111010" => rgb <= "000000";
					when "01110001001111011" => rgb <= "000000";
					when "01110001001111100" => rgb <= "000000";
					when "01110001001111101" => rgb <= "000000";
					when "01110001001111110" => rgb <= "000000";
					when "01110001001111111" => rgb <= "000000";
					when "01110001010000000" => rgb <= "000000";
					when "01110001010000001" => rgb <= "000000";
					when "01110001010000010" => rgb <= "000000";
					when "01110001010000011" => rgb <= "000000";
					when "01110001010000100" => rgb <= "000000";
					when "01110001010000101" => rgb <= "000000";
					when "01110001010000110" => rgb <= "000000";
					when "01110001010000111" => rgb <= "000000";
					when "01110001010001000" => rgb <= "010100";
					when "01110001010001001" => rgb <= "101000";
					when "01110001010001010" => rgb <= "101000";
					when "01110001010001011" => rgb <= "101000";
					when "01110001010001100" => rgb <= "101000";
					when "01110001010001101" => rgb <= "101000";
					when "01110001010001110" => rgb <= "101000";
					when "01110001010001111" => rgb <= "101000";
					when "01110001010010000" => rgb <= "101000";
					when "01110001010010001" => rgb <= "101000";
					when "01110001010010010" => rgb <= "101000";
					when "01110001010010011" => rgb <= "101000";
					when "01110001010010100" => rgb <= "101000";
					when "01110001010010101" => rgb <= "101000";
					when "01110001010010110" => rgb <= "101000";
					when "01110001010010111" => rgb <= "101000";
					when "01110001010011000" => rgb <= "101000";
					when "01110001010011001" => rgb <= "101000";
					when "01110001010011010" => rgb <= "101000";
					when "01110001010011011" => rgb <= "101000";
					when "01110001010011100" => rgb <= "101000";
					when "01110001010011101" => rgb <= "101000";
					when "01110001010011110" => rgb <= "101000";
					when "01110001010011111" => rgb <= "101000";
					when "01110001010100000" => rgb <= "101000";
					when "01110001010100001" => rgb <= "101000";
					when "01110001010100010" => rgb <= "101000";
					when "01110001010100011" => rgb <= "101000";
					when "01110001010100100" => rgb <= "101000";
					when "01110001010100101" => rgb <= "101000";
					when "01110001010100110" => rgb <= "101000";
					when "01110001010100111" => rgb <= "101000";
					when "01110001010101000" => rgb <= "101000";
					when "01110001010101001" => rgb <= "101000";
					when "01110001010101010" => rgb <= "101000";
					when "01110001010101011" => rgb <= "101000";
					when "01110001010101100" => rgb <= "101000";
					when "01110001010101101" => rgb <= "101000";
					when "01110001010101110" => rgb <= "101000";
					when "01110001010101111" => rgb <= "101000";
					when "01110001010110000" => rgb <= "101000";
					when "01110001010110001" => rgb <= "101000";
					when "01110001010110010" => rgb <= "101000";
					when "01110001010110011" => rgb <= "101000";
					when "01110001010110100" => rgb <= "101000";
					when "01110001010110101" => rgb <= "010100";
					when "01110001010110110" => rgb <= "000000";
					when "01110001010110111" => rgb <= "000000";
					when "01110001010111000" => rgb <= "000000";
					when "01110001010111001" => rgb <= "000000";
					when "01110001010111010" => rgb <= "000000";
					when "01110001010111011" => rgb <= "000000";
					when "01110001010111100" => rgb <= "000000";
					when "01110001010111101" => rgb <= "000000";
					when "01110001010111110" => rgb <= "000000";
					when "01110001010111111" => rgb <= "000000";
					when "01110001011000000" => rgb <= "000000";
					when "01110001011000001" => rgb <= "000000";
					when "01110001011000010" => rgb <= "000000";
					when "01110001011000011" => rgb <= "000000";
					when "01110001011000100" => rgb <= "000000";
					when "01110001011000101" => rgb <= "000000";
					when "01110001011000110" => rgb <= "000000";
					when "01110001011000111" => rgb <= "000000";
					when "01110001011001000" => rgb <= "000000";
					when "01110001011001001" => rgb <= "000000";
					when "01110001011001010" => rgb <= "000000";
					when "01110001011001011" => rgb <= "000000";
					when "01110001011001100" => rgb <= "000000";
					when "01110001011001101" => rgb <= "000000";
					when "01110001011001110" => rgb <= "000000";
					when "01110001011001111" => rgb <= "000000";
					when "01110001011010000" => rgb <= "000000";
					when "01110001011010001" => rgb <= "000000";
					when "01110001011010010" => rgb <= "000000";
					when "01110001011010011" => rgb <= "000000";
					when "01110001011010100" => rgb <= "000000";
					when "01110001011010101" => rgb <= "000000";
					when "01110001011010110" => rgb <= "000000";
					when "01110001011010111" => rgb <= "000000";
					when "01110001011011000" => rgb <= "000000";
					when "01110001011011001" => rgb <= "000000";
					when "01110001011011010" => rgb <= "000000";
					when "01110001011011011" => rgb <= "000000";
					when "01110001011011100" => rgb <= "000000";
					when "01110001011011101" => rgb <= "000000";
					when "01110001011011110" => rgb <= "000000";
					when "01110001011011111" => rgb <= "000000";
					when "01110001011100000" => rgb <= "000000";
					when "01110001011100001" => rgb <= "000000";
					when "01110001011100010" => rgb <= "000000";
					when "01110001011100011" => rgb <= "000000";
					when "01110001011100100" => rgb <= "000000";
					when "01110001011100101" => rgb <= "000000";
					when "01110001011100110" => rgb <= "000000";
					when "01110001011100111" => rgb <= "000000";
					when "01110001011101000" => rgb <= "000000";
					when "01110001011101001" => rgb <= "000000";
					when "01110001011101010" => rgb <= "000000";
					when "01110001011101011" => rgb <= "000000";
					when "01110001011101100" => rgb <= "000000";
					when "01110001011101101" => rgb <= "000000";
					when "01110001011101110" => rgb <= "000000";
					when "01110001011101111" => rgb <= "000000";
					when "01110001011110000" => rgb <= "000000";
					when "01110001011110001" => rgb <= "000000";
					when "01110001011110010" => rgb <= "000000";
					when "01110001011110011" => rgb <= "000000";
					when "01110001011110100" => rgb <= "000000";
					when "01110001011110101" => rgb <= "000000";
					when "01110001011110110" => rgb <= "000000";
					when "01110001011110111" => rgb <= "000000";
					when "01110001011111000" => rgb <= "000000";
					when "01110001011111001" => rgb <= "000000";
					when "01110001011111010" => rgb <= "000000";
					when "01110001011111011" => rgb <= "000000";
					when "01110001011111100" => rgb <= "000000";
					when "01110001011111101" => rgb <= "000000";
					when "01110001011111110" => rgb <= "000000";
					when "01110001011111111" => rgb <= "000000";
					when "01110001100000000" => rgb <= "000000";
					when "01110001100000001" => rgb <= "000000";
					when "01110001100000010" => rgb <= "000000";
					when "01110001100000011" => rgb <= "000000";
					when "01110001100000100" => rgb <= "000000";
					when "01110001100000101" => rgb <= "000000";
					when "01110001100000110" => rgb <= "000000";
					when "01110001100000111" => rgb <= "000000";
					when "01110001100001000" => rgb <= "000000";
					when "01110001100001001" => rgb <= "000000";
					when "01110001100001010" => rgb <= "000000";
					when "01110001100001011" => rgb <= "000000";
					when "01110001100001100" => rgb <= "000000";
					when "01110001100001101" => rgb <= "000000";
					when "01110001100001110" => rgb <= "000000";
					when "01110001100001111" => rgb <= "000000";
					when "01110001100010000" => rgb <= "000000";
					when "01110001100010001" => rgb <= "000000";
					when "01110001100010010" => rgb <= "000000";
					when "01110001100010011" => rgb <= "000000";
					when "01110001100010100" => rgb <= "000000";
					when "01110001100010101" => rgb <= "000000";
					when "01110001100010110" => rgb <= "000000";
					when "01110001100010111" => rgb <= "000000";
					when "01110001100011000" => rgb <= "000000";
					when "01110001100011001" => rgb <= "000000";
					when "01110001100011010" => rgb <= "000000";
					when "01110001100011011" => rgb <= "000000";
					when "01110001100011100" => rgb <= "000000";
					when "01110001100011101" => rgb <= "000000";
					when "01110001100011110" => rgb <= "000000";
					when "01110001100011111" => rgb <= "000000";
					when "01110001100100000" => rgb <= "000000";
					when "01110001100100001" => rgb <= "000000";
					when "01110001100100010" => rgb <= "000000";
					when "01110001100100011" => rgb <= "000000";
					when "01110001100100100" => rgb <= "000000";
					when "01110001100100101" => rgb <= "000000";
					when "01110001100100110" => rgb <= "000000";
					when "01110001100100111" => rgb <= "000000";
					when "01110001100101000" => rgb <= "000000";
					when "01110001100101001" => rgb <= "000000";
					when "01110001100101010" => rgb <= "000000";
					when "01110001100101011" => rgb <= "000000";
					when "01110001100101100" => rgb <= "000000";
					when "01110001100101101" => rgb <= "000000";
					when "01110001100101110" => rgb <= "000000";
					when "01110001100101111" => rgb <= "000000";
					when "01110001100110000" => rgb <= "000000";
					when "01110001100110001" => rgb <= "000000";
					when "01110001100110010" => rgb <= "000000";
					when "01110001100110011" => rgb <= "000000";
					when "01110001100110100" => rgb <= "000000";
					when "01110001100110101" => rgb <= "000000";
					when "01110001100110110" => rgb <= "000000";
					when "01110001100110111" => rgb <= "000000";
					when "01110001100111000" => rgb <= "000000";
					when "01110001100111001" => rgb <= "000000";
					when "01110001100111010" => rgb <= "000000";
					when "01110001100111011" => rgb <= "000000";
					when "01110001100111100" => rgb <= "000000";
					when "01110001100111101" => rgb <= "000000";
					when "01110001100111110" => rgb <= "000000";
					when "01110001100111111" => rgb <= "000000";
					when "01110010000000000" => rgb <= "000000";
					when "01110010000000001" => rgb <= "000000";
					when "01110010000000010" => rgb <= "000000";
					when "01110010000000011" => rgb <= "000000";
					when "01110010000000100" => rgb <= "000000";
					when "01110010000000101" => rgb <= "000000";
					when "01110010000000110" => rgb <= "000000";
					when "01110010000000111" => rgb <= "000000";
					when "01110010000001000" => rgb <= "000000";
					when "01110010000001001" => rgb <= "000000";
					when "01110010000001010" => rgb <= "000000";
					when "01110010000001011" => rgb <= "000000";
					when "01110010000001100" => rgb <= "000000";
					when "01110010000001101" => rgb <= "000000";
					when "01110010000001110" => rgb <= "000000";
					when "01110010000001111" => rgb <= "000000";
					when "01110010000010000" => rgb <= "000000";
					when "01110010000010001" => rgb <= "000000";
					when "01110010000010010" => rgb <= "000000";
					when "01110010000010011" => rgb <= "000000";
					when "01110010000010100" => rgb <= "000000";
					when "01110010000010101" => rgb <= "000000";
					when "01110010000010110" => rgb <= "000000";
					when "01110010000010111" => rgb <= "000000";
					when "01110010000011000" => rgb <= "000000";
					when "01110010000011001" => rgb <= "000000";
					when "01110010000011010" => rgb <= "000000";
					when "01110010000011011" => rgb <= "000000";
					when "01110010000011100" => rgb <= "000000";
					when "01110010000011101" => rgb <= "000000";
					when "01110010000011110" => rgb <= "000000";
					when "01110010000011111" => rgb <= "000000";
					when "01110010000100000" => rgb <= "000000";
					when "01110010000100001" => rgb <= "000000";
					when "01110010000100010" => rgb <= "000000";
					when "01110010000100011" => rgb <= "000000";
					when "01110010000100100" => rgb <= "000000";
					when "01110010000100101" => rgb <= "000000";
					when "01110010000100110" => rgb <= "000000";
					when "01110010000100111" => rgb <= "000000";
					when "01110010000101000" => rgb <= "000000";
					when "01110010000101001" => rgb <= "000000";
					when "01110010000101010" => rgb <= "000000";
					when "01110010000101011" => rgb <= "000000";
					when "01110010000101100" => rgb <= "000000";
					when "01110010000101101" => rgb <= "000000";
					when "01110010000101110" => rgb <= "000000";
					when "01110010000101111" => rgb <= "000000";
					when "01110010000110000" => rgb <= "000000";
					when "01110010000110001" => rgb <= "000000";
					when "01110010000110010" => rgb <= "000000";
					when "01110010000110011" => rgb <= "000000";
					when "01110010000110100" => rgb <= "000000";
					when "01110010000110101" => rgb <= "000000";
					when "01110010000110110" => rgb <= "000000";
					when "01110010000110111" => rgb <= "000000";
					when "01110010000111000" => rgb <= "000000";
					when "01110010000111001" => rgb <= "000000";
					when "01110010000111010" => rgb <= "000000";
					when "01110010000111011" => rgb <= "000000";
					when "01110010000111100" => rgb <= "000000";
					when "01110010000111101" => rgb <= "000000";
					when "01110010000111110" => rgb <= "000000";
					when "01110010000111111" => rgb <= "000000";
					when "01110010001000000" => rgb <= "000000";
					when "01110010001000001" => rgb <= "000000";
					when "01110010001000010" => rgb <= "000000";
					when "01110010001000011" => rgb <= "000000";
					when "01110010001000100" => rgb <= "000000";
					when "01110010001000101" => rgb <= "000000";
					when "01110010001000110" => rgb <= "000000";
					when "01110010001000111" => rgb <= "000000";
					when "01110010001001000" => rgb <= "000000";
					when "01110010001001001" => rgb <= "000000";
					when "01110010001001010" => rgb <= "000000";
					when "01110010001001011" => rgb <= "000000";
					when "01110010001001100" => rgb <= "000000";
					when "01110010001001101" => rgb <= "000000";
					when "01110010001001110" => rgb <= "000000";
					when "01110010001001111" => rgb <= "000000";
					when "01110010001010000" => rgb <= "000000";
					when "01110010001010001" => rgb <= "000000";
					when "01110010001010010" => rgb <= "000000";
					when "01110010001010011" => rgb <= "000000";
					when "01110010001010100" => rgb <= "000000";
					when "01110010001010101" => rgb <= "000000";
					when "01110010001010110" => rgb <= "000000";
					when "01110010001010111" => rgb <= "000000";
					when "01110010001011000" => rgb <= "000000";
					when "01110010001011001" => rgb <= "000000";
					when "01110010001011010" => rgb <= "000000";
					when "01110010001011011" => rgb <= "000000";
					when "01110010001011100" => rgb <= "000000";
					when "01110010001011101" => rgb <= "000000";
					when "01110010001011110" => rgb <= "000000";
					when "01110010001011111" => rgb <= "000000";
					when "01110010001100000" => rgb <= "000000";
					when "01110010001100001" => rgb <= "000000";
					when "01110010001100010" => rgb <= "000000";
					when "01110010001100011" => rgb <= "000000";
					when "01110010001100100" => rgb <= "000000";
					when "01110010001100101" => rgb <= "000000";
					when "01110010001100110" => rgb <= "000000";
					when "01110010001100111" => rgb <= "000000";
					when "01110010001101000" => rgb <= "000000";
					when "01110010001101001" => rgb <= "000000";
					when "01110010001101010" => rgb <= "000000";
					when "01110010001101011" => rgb <= "000000";
					when "01110010001101100" => rgb <= "000000";
					when "01110010001101101" => rgb <= "000000";
					when "01110010001101110" => rgb <= "000000";
					when "01110010001101111" => rgb <= "000000";
					when "01110010001110000" => rgb <= "000000";
					when "01110010001110001" => rgb <= "000000";
					when "01110010001110010" => rgb <= "000000";
					when "01110010001110011" => rgb <= "000000";
					when "01110010001110100" => rgb <= "000000";
					when "01110010001110101" => rgb <= "000000";
					when "01110010001110110" => rgb <= "000000";
					when "01110010001110111" => rgb <= "000000";
					when "01110010001111000" => rgb <= "000000";
					when "01110010001111001" => rgb <= "000000";
					when "01110010001111010" => rgb <= "000000";
					when "01110010001111011" => rgb <= "000000";
					when "01110010001111100" => rgb <= "000000";
					when "01110010001111101" => rgb <= "000000";
					when "01110010001111110" => rgb <= "000000";
					when "01110010001111111" => rgb <= "000000";
					when "01110010010000000" => rgb <= "000000";
					when "01110010010000001" => rgb <= "000000";
					when "01110010010000010" => rgb <= "000000";
					when "01110010010000011" => rgb <= "000000";
					when "01110010010000100" => rgb <= "000000";
					when "01110010010000101" => rgb <= "000000";
					when "01110010010000110" => rgb <= "000000";
					when "01110010010000111" => rgb <= "000000";
					when "01110010010001000" => rgb <= "010100";
					when "01110010010001001" => rgb <= "101000";
					when "01110010010001010" => rgb <= "101000";
					when "01110010010001011" => rgb <= "101000";
					when "01110010010001100" => rgb <= "101000";
					when "01110010010001101" => rgb <= "101000";
					when "01110010010001110" => rgb <= "101000";
					when "01110010010001111" => rgb <= "101000";
					when "01110010010010000" => rgb <= "101000";
					when "01110010010010001" => rgb <= "101000";
					when "01110010010010010" => rgb <= "101000";
					when "01110010010010011" => rgb <= "101000";
					when "01110010010010100" => rgb <= "101000";
					when "01110010010010101" => rgb <= "101000";
					when "01110010010010110" => rgb <= "101000";
					when "01110010010010111" => rgb <= "101000";
					when "01110010010011000" => rgb <= "101000";
					when "01110010010011001" => rgb <= "101000";
					when "01110010010011010" => rgb <= "101000";
					when "01110010010011011" => rgb <= "101000";
					when "01110010010011100" => rgb <= "101000";
					when "01110010010011101" => rgb <= "101000";
					when "01110010010011110" => rgb <= "101000";
					when "01110010010011111" => rgb <= "101000";
					when "01110010010100000" => rgb <= "101000";
					when "01110010010100001" => rgb <= "101000";
					when "01110010010100010" => rgb <= "101000";
					when "01110010010100011" => rgb <= "101000";
					when "01110010010100100" => rgb <= "101000";
					when "01110010010100101" => rgb <= "101000";
					when "01110010010100110" => rgb <= "101000";
					when "01110010010100111" => rgb <= "101000";
					when "01110010010101000" => rgb <= "101000";
					when "01110010010101001" => rgb <= "101000";
					when "01110010010101010" => rgb <= "101000";
					when "01110010010101011" => rgb <= "101000";
					when "01110010010101100" => rgb <= "101000";
					when "01110010010101101" => rgb <= "101000";
					when "01110010010101110" => rgb <= "101000";
					when "01110010010101111" => rgb <= "101000";
					when "01110010010110000" => rgb <= "101000";
					when "01110010010110001" => rgb <= "101000";
					when "01110010010110010" => rgb <= "101000";
					when "01110010010110011" => rgb <= "101000";
					when "01110010010110100" => rgb <= "101000";
					when "01110010010110101" => rgb <= "010100";
					when "01110010010110110" => rgb <= "000000";
					when "01110010010110111" => rgb <= "000000";
					when "01110010010111000" => rgb <= "000000";
					when "01110010010111001" => rgb <= "000000";
					when "01110010010111010" => rgb <= "000000";
					when "01110010010111011" => rgb <= "000000";
					when "01110010010111100" => rgb <= "000000";
					when "01110010010111101" => rgb <= "000000";
					when "01110010010111110" => rgb <= "000000";
					when "01110010010111111" => rgb <= "000000";
					when "01110010011000000" => rgb <= "000000";
					when "01110010011000001" => rgb <= "000000";
					when "01110010011000010" => rgb <= "000000";
					when "01110010011000011" => rgb <= "000000";
					when "01110010011000100" => rgb <= "000000";
					when "01110010011000101" => rgb <= "000000";
					when "01110010011000110" => rgb <= "000000";
					when "01110010011000111" => rgb <= "000000";
					when "01110010011001000" => rgb <= "000000";
					when "01110010011001001" => rgb <= "000000";
					when "01110010011001010" => rgb <= "000000";
					when "01110010011001011" => rgb <= "000000";
					when "01110010011001100" => rgb <= "000000";
					when "01110010011001101" => rgb <= "000000";
					when "01110010011001110" => rgb <= "000000";
					when "01110010011001111" => rgb <= "000000";
					when "01110010011010000" => rgb <= "000000";
					when "01110010011010001" => rgb <= "000000";
					when "01110010011010010" => rgb <= "000000";
					when "01110010011010011" => rgb <= "000000";
					when "01110010011010100" => rgb <= "000000";
					when "01110010011010101" => rgb <= "000000";
					when "01110010011010110" => rgb <= "000000";
					when "01110010011010111" => rgb <= "000000";
					when "01110010011011000" => rgb <= "000000";
					when "01110010011011001" => rgb <= "000000";
					when "01110010011011010" => rgb <= "000000";
					when "01110010011011011" => rgb <= "000000";
					when "01110010011011100" => rgb <= "000000";
					when "01110010011011101" => rgb <= "000000";
					when "01110010011011110" => rgb <= "000000";
					when "01110010011011111" => rgb <= "000000";
					when "01110010011100000" => rgb <= "000000";
					when "01110010011100001" => rgb <= "000000";
					when "01110010011100010" => rgb <= "000000";
					when "01110010011100011" => rgb <= "000000";
					when "01110010011100100" => rgb <= "000000";
					when "01110010011100101" => rgb <= "000000";
					when "01110010011100110" => rgb <= "000000";
					when "01110010011100111" => rgb <= "000000";
					when "01110010011101000" => rgb <= "000000";
					when "01110010011101001" => rgb <= "000000";
					when "01110010011101010" => rgb <= "000000";
					when "01110010011101011" => rgb <= "000000";
					when "01110010011101100" => rgb <= "000000";
					when "01110010011101101" => rgb <= "000000";
					when "01110010011101110" => rgb <= "000000";
					when "01110010011101111" => rgb <= "000000";
					when "01110010011110000" => rgb <= "000000";
					when "01110010011110001" => rgb <= "000000";
					when "01110010011110010" => rgb <= "000000";
					when "01110010011110011" => rgb <= "000000";
					when "01110010011110100" => rgb <= "000000";
					when "01110010011110101" => rgb <= "000000";
					when "01110010011110110" => rgb <= "000000";
					when "01110010011110111" => rgb <= "000000";
					when "01110010011111000" => rgb <= "000000";
					when "01110010011111001" => rgb <= "000000";
					when "01110010011111010" => rgb <= "000000";
					when "01110010011111011" => rgb <= "000000";
					when "01110010011111100" => rgb <= "000000";
					when "01110010011111101" => rgb <= "000000";
					when "01110010011111110" => rgb <= "000000";
					when "01110010011111111" => rgb <= "000000";
					when "01110010100000000" => rgb <= "000000";
					when "01110010100000001" => rgb <= "000000";
					when "01110010100000010" => rgb <= "000000";
					when "01110010100000011" => rgb <= "000000";
					when "01110010100000100" => rgb <= "000000";
					when "01110010100000101" => rgb <= "000000";
					when "01110010100000110" => rgb <= "000000";
					when "01110010100000111" => rgb <= "000000";
					when "01110010100001000" => rgb <= "000000";
					when "01110010100001001" => rgb <= "000000";
					when "01110010100001010" => rgb <= "000000";
					when "01110010100001011" => rgb <= "000000";
					when "01110010100001100" => rgb <= "000000";
					when "01110010100001101" => rgb <= "000000";
					when "01110010100001110" => rgb <= "000000";
					when "01110010100001111" => rgb <= "000000";
					when "01110010100010000" => rgb <= "000000";
					when "01110010100010001" => rgb <= "000000";
					when "01110010100010010" => rgb <= "000000";
					when "01110010100010011" => rgb <= "000000";
					when "01110010100010100" => rgb <= "000000";
					when "01110010100010101" => rgb <= "000000";
					when "01110010100010110" => rgb <= "000000";
					when "01110010100010111" => rgb <= "000000";
					when "01110010100011000" => rgb <= "000000";
					when "01110010100011001" => rgb <= "000000";
					when "01110010100011010" => rgb <= "000000";
					when "01110010100011011" => rgb <= "000000";
					when "01110010100011100" => rgb <= "000000";
					when "01110010100011101" => rgb <= "000000";
					when "01110010100011110" => rgb <= "000000";
					when "01110010100011111" => rgb <= "000000";
					when "01110010100100000" => rgb <= "000000";
					when "01110010100100001" => rgb <= "000000";
					when "01110010100100010" => rgb <= "000000";
					when "01110010100100011" => rgb <= "000000";
					when "01110010100100100" => rgb <= "000000";
					when "01110010100100101" => rgb <= "000000";
					when "01110010100100110" => rgb <= "000000";
					when "01110010100100111" => rgb <= "000000";
					when "01110010100101000" => rgb <= "000000";
					when "01110010100101001" => rgb <= "000000";
					when "01110010100101010" => rgb <= "000000";
					when "01110010100101011" => rgb <= "000000";
					when "01110010100101100" => rgb <= "000000";
					when "01110010100101101" => rgb <= "000000";
					when "01110010100101110" => rgb <= "000000";
					when "01110010100101111" => rgb <= "000000";
					when "01110010100110000" => rgb <= "000000";
					when "01110010100110001" => rgb <= "000000";
					when "01110010100110010" => rgb <= "000000";
					when "01110010100110011" => rgb <= "000000";
					when "01110010100110100" => rgb <= "000000";
					when "01110010100110101" => rgb <= "000000";
					when "01110010100110110" => rgb <= "000000";
					when "01110010100110111" => rgb <= "000000";
					when "01110010100111000" => rgb <= "000000";
					when "01110010100111001" => rgb <= "000000";
					when "01110010100111010" => rgb <= "000000";
					when "01110010100111011" => rgb <= "000000";
					when "01110010100111100" => rgb <= "000000";
					when "01110010100111101" => rgb <= "000000";
					when "01110010100111110" => rgb <= "000000";
					when "01110010100111111" => rgb <= "000000";
					when "01110011000000000" => rgb <= "000000";
					when "01110011000000001" => rgb <= "000000";
					when "01110011000000010" => rgb <= "000000";
					when "01110011000000011" => rgb <= "000000";
					when "01110011000000100" => rgb <= "000000";
					when "01110011000000101" => rgb <= "000000";
					when "01110011000000110" => rgb <= "000000";
					when "01110011000000111" => rgb <= "000000";
					when "01110011000001000" => rgb <= "000000";
					when "01110011000001001" => rgb <= "000000";
					when "01110011000001010" => rgb <= "000000";
					when "01110011000001011" => rgb <= "000000";
					when "01110011000001100" => rgb <= "000000";
					when "01110011000001101" => rgb <= "000000";
					when "01110011000001110" => rgb <= "000000";
					when "01110011000001111" => rgb <= "000000";
					when "01110011000010000" => rgb <= "000000";
					when "01110011000010001" => rgb <= "000000";
					when "01110011000010010" => rgb <= "000000";
					when "01110011000010011" => rgb <= "000000";
					when "01110011000010100" => rgb <= "000000";
					when "01110011000010101" => rgb <= "000000";
					when "01110011000010110" => rgb <= "000000";
					when "01110011000010111" => rgb <= "000000";
					when "01110011000011000" => rgb <= "000000";
					when "01110011000011001" => rgb <= "000000";
					when "01110011000011010" => rgb <= "000000";
					when "01110011000011011" => rgb <= "000000";
					when "01110011000011100" => rgb <= "000000";
					when "01110011000011101" => rgb <= "000000";
					when "01110011000011110" => rgb <= "000000";
					when "01110011000011111" => rgb <= "000000";
					when "01110011000100000" => rgb <= "000000";
					when "01110011000100001" => rgb <= "000000";
					when "01110011000100010" => rgb <= "000000";
					when "01110011000100011" => rgb <= "000000";
					when "01110011000100100" => rgb <= "000000";
					when "01110011000100101" => rgb <= "000000";
					when "01110011000100110" => rgb <= "000000";
					when "01110011000100111" => rgb <= "000000";
					when "01110011000101000" => rgb <= "000000";
					when "01110011000101001" => rgb <= "000000";
					when "01110011000101010" => rgb <= "000000";
					when "01110011000101011" => rgb <= "000000";
					when "01110011000101100" => rgb <= "000000";
					when "01110011000101101" => rgb <= "000000";
					when "01110011000101110" => rgb <= "000000";
					when "01110011000101111" => rgb <= "000000";
					when "01110011000110000" => rgb <= "000000";
					when "01110011000110001" => rgb <= "000000";
					when "01110011000110010" => rgb <= "000000";
					when "01110011000110011" => rgb <= "000000";
					when "01110011000110100" => rgb <= "000000";
					when "01110011000110101" => rgb <= "000000";
					when "01110011000110110" => rgb <= "000000";
					when "01110011000110111" => rgb <= "000000";
					when "01110011000111000" => rgb <= "000000";
					when "01110011000111001" => rgb <= "000000";
					when "01110011000111010" => rgb <= "000000";
					when "01110011000111011" => rgb <= "000000";
					when "01110011000111100" => rgb <= "000000";
					when "01110011000111101" => rgb <= "000000";
					when "01110011000111110" => rgb <= "000000";
					when "01110011000111111" => rgb <= "000000";
					when "01110011001000000" => rgb <= "000000";
					when "01110011001000001" => rgb <= "000000";
					when "01110011001000010" => rgb <= "000000";
					when "01110011001000011" => rgb <= "000000";
					when "01110011001000100" => rgb <= "000000";
					when "01110011001000101" => rgb <= "000000";
					when "01110011001000110" => rgb <= "000000";
					when "01110011001000111" => rgb <= "000000";
					when "01110011001001000" => rgb <= "000000";
					when "01110011001001001" => rgb <= "000000";
					when "01110011001001010" => rgb <= "000000";
					when "01110011001001011" => rgb <= "000000";
					when "01110011001001100" => rgb <= "000000";
					when "01110011001001101" => rgb <= "000000";
					when "01110011001001110" => rgb <= "000000";
					when "01110011001001111" => rgb <= "000000";
					when "01110011001010000" => rgb <= "000000";
					when "01110011001010001" => rgb <= "000000";
					when "01110011001010010" => rgb <= "000000";
					when "01110011001010011" => rgb <= "000000";
					when "01110011001010100" => rgb <= "000000";
					when "01110011001010101" => rgb <= "000000";
					when "01110011001010110" => rgb <= "000000";
					when "01110011001010111" => rgb <= "000000";
					when "01110011001011000" => rgb <= "000000";
					when "01110011001011001" => rgb <= "000000";
					when "01110011001011010" => rgb <= "000000";
					when "01110011001011011" => rgb <= "000000";
					when "01110011001011100" => rgb <= "000000";
					when "01110011001011101" => rgb <= "000000";
					when "01110011001011110" => rgb <= "000000";
					when "01110011001011111" => rgb <= "000000";
					when "01110011001100000" => rgb <= "000000";
					when "01110011001100001" => rgb <= "000000";
					when "01110011001100010" => rgb <= "000000";
					when "01110011001100011" => rgb <= "000000";
					when "01110011001100100" => rgb <= "000000";
					when "01110011001100101" => rgb <= "000000";
					when "01110011001100110" => rgb <= "000000";
					when "01110011001100111" => rgb <= "000000";
					when "01110011001101000" => rgb <= "000000";
					when "01110011001101001" => rgb <= "000000";
					when "01110011001101010" => rgb <= "000000";
					when "01110011001101011" => rgb <= "000000";
					when "01110011001101100" => rgb <= "000000";
					when "01110011001101101" => rgb <= "000000";
					when "01110011001101110" => rgb <= "000000";
					when "01110011001101111" => rgb <= "000000";
					when "01110011001110000" => rgb <= "000000";
					when "01110011001110001" => rgb <= "000000";
					when "01110011001110010" => rgb <= "000000";
					when "01110011001110011" => rgb <= "000000";
					when "01110011001110100" => rgb <= "000000";
					when "01110011001110101" => rgb <= "000000";
					when "01110011001110110" => rgb <= "000000";
					when "01110011001110111" => rgb <= "000000";
					when "01110011001111000" => rgb <= "000000";
					when "01110011001111001" => rgb <= "000000";
					when "01110011001111010" => rgb <= "000000";
					when "01110011001111011" => rgb <= "000000";
					when "01110011001111100" => rgb <= "000000";
					when "01110011001111101" => rgb <= "000000";
					when "01110011001111110" => rgb <= "000000";
					when "01110011001111111" => rgb <= "000000";
					when "01110011010000000" => rgb <= "000000";
					when "01110011010000001" => rgb <= "000000";
					when "01110011010000010" => rgb <= "000000";
					when "01110011010000011" => rgb <= "000000";
					when "01110011010000100" => rgb <= "000000";
					when "01110011010000101" => rgb <= "000000";
					when "01110011010000110" => rgb <= "000000";
					when "01110011010000111" => rgb <= "000000";
					when "01110011010001000" => rgb <= "010100";
					when "01110011010001001" => rgb <= "101000";
					when "01110011010001010" => rgb <= "101000";
					when "01110011010001011" => rgb <= "101000";
					when "01110011010001100" => rgb <= "101000";
					when "01110011010001101" => rgb <= "101000";
					when "01110011010001110" => rgb <= "101000";
					when "01110011010001111" => rgb <= "101000";
					when "01110011010010000" => rgb <= "101000";
					when "01110011010010001" => rgb <= "101000";
					when "01110011010010010" => rgb <= "101000";
					when "01110011010010011" => rgb <= "101000";
					when "01110011010010100" => rgb <= "101000";
					when "01110011010010101" => rgb <= "101000";
					when "01110011010010110" => rgb <= "101000";
					when "01110011010010111" => rgb <= "101000";
					when "01110011010011000" => rgb <= "101000";
					when "01110011010011001" => rgb <= "101000";
					when "01110011010011010" => rgb <= "101000";
					when "01110011010011011" => rgb <= "101000";
					when "01110011010011100" => rgb <= "101000";
					when "01110011010011101" => rgb <= "101000";
					when "01110011010011110" => rgb <= "101000";
					when "01110011010011111" => rgb <= "101000";
					when "01110011010100000" => rgb <= "101000";
					when "01110011010100001" => rgb <= "101000";
					when "01110011010100010" => rgb <= "101000";
					when "01110011010100011" => rgb <= "101000";
					when "01110011010100100" => rgb <= "101000";
					when "01110011010100101" => rgb <= "101000";
					when "01110011010100110" => rgb <= "101000";
					when "01110011010100111" => rgb <= "101000";
					when "01110011010101000" => rgb <= "101000";
					when "01110011010101001" => rgb <= "101000";
					when "01110011010101010" => rgb <= "101000";
					when "01110011010101011" => rgb <= "101000";
					when "01110011010101100" => rgb <= "101000";
					when "01110011010101101" => rgb <= "101000";
					when "01110011010101110" => rgb <= "101000";
					when "01110011010101111" => rgb <= "101000";
					when "01110011010110000" => rgb <= "101000";
					when "01110011010110001" => rgb <= "101000";
					when "01110011010110010" => rgb <= "101000";
					when "01110011010110011" => rgb <= "101000";
					when "01110011010110100" => rgb <= "101000";
					when "01110011010110101" => rgb <= "010100";
					when "01110011010110110" => rgb <= "000000";
					when "01110011010110111" => rgb <= "000000";
					when "01110011010111000" => rgb <= "000000";
					when "01110011010111001" => rgb <= "000000";
					when "01110011010111010" => rgb <= "000000";
					when "01110011010111011" => rgb <= "000000";
					when "01110011010111100" => rgb <= "000000";
					when "01110011010111101" => rgb <= "000000";
					when "01110011010111110" => rgb <= "000000";
					when "01110011010111111" => rgb <= "000000";
					when "01110011011000000" => rgb <= "000000";
					when "01110011011000001" => rgb <= "000000";
					when "01110011011000010" => rgb <= "000000";
					when "01110011011000011" => rgb <= "000000";
					when "01110011011000100" => rgb <= "000000";
					when "01110011011000101" => rgb <= "000000";
					when "01110011011000110" => rgb <= "000000";
					when "01110011011000111" => rgb <= "000000";
					when "01110011011001000" => rgb <= "000000";
					when "01110011011001001" => rgb <= "000000";
					when "01110011011001010" => rgb <= "000000";
					when "01110011011001011" => rgb <= "000000";
					when "01110011011001100" => rgb <= "000000";
					when "01110011011001101" => rgb <= "000000";
					when "01110011011001110" => rgb <= "000000";
					when "01110011011001111" => rgb <= "000000";
					when "01110011011010000" => rgb <= "000000";
					when "01110011011010001" => rgb <= "000000";
					when "01110011011010010" => rgb <= "000000";
					when "01110011011010011" => rgb <= "000000";
					when "01110011011010100" => rgb <= "000000";
					when "01110011011010101" => rgb <= "000000";
					when "01110011011010110" => rgb <= "000000";
					when "01110011011010111" => rgb <= "000000";
					when "01110011011011000" => rgb <= "000000";
					when "01110011011011001" => rgb <= "000000";
					when "01110011011011010" => rgb <= "000000";
					when "01110011011011011" => rgb <= "000000";
					when "01110011011011100" => rgb <= "000000";
					when "01110011011011101" => rgb <= "000000";
					when "01110011011011110" => rgb <= "000000";
					when "01110011011011111" => rgb <= "000000";
					when "01110011011100000" => rgb <= "000000";
					when "01110011011100001" => rgb <= "000000";
					when "01110011011100010" => rgb <= "000000";
					when "01110011011100011" => rgb <= "000000";
					when "01110011011100100" => rgb <= "000000";
					when "01110011011100101" => rgb <= "000000";
					when "01110011011100110" => rgb <= "000000";
					when "01110011011100111" => rgb <= "000000";
					when "01110011011101000" => rgb <= "000000";
					when "01110011011101001" => rgb <= "000000";
					when "01110011011101010" => rgb <= "000000";
					when "01110011011101011" => rgb <= "000000";
					when "01110011011101100" => rgb <= "000000";
					when "01110011011101101" => rgb <= "000000";
					when "01110011011101110" => rgb <= "000000";
					when "01110011011101111" => rgb <= "000000";
					when "01110011011110000" => rgb <= "000000";
					when "01110011011110001" => rgb <= "000000";
					when "01110011011110010" => rgb <= "000000";
					when "01110011011110011" => rgb <= "000000";
					when "01110011011110100" => rgb <= "000000";
					when "01110011011110101" => rgb <= "000000";
					when "01110011011110110" => rgb <= "000000";
					when "01110011011110111" => rgb <= "000000";
					when "01110011011111000" => rgb <= "000000";
					when "01110011011111001" => rgb <= "000000";
					when "01110011011111010" => rgb <= "000000";
					when "01110011011111011" => rgb <= "000000";
					when "01110011011111100" => rgb <= "000000";
					when "01110011011111101" => rgb <= "000000";
					when "01110011011111110" => rgb <= "000000";
					when "01110011011111111" => rgb <= "000000";
					when "01110011100000000" => rgb <= "000000";
					when "01110011100000001" => rgb <= "000000";
					when "01110011100000010" => rgb <= "000000";
					when "01110011100000011" => rgb <= "000000";
					when "01110011100000100" => rgb <= "000000";
					when "01110011100000101" => rgb <= "000000";
					when "01110011100000110" => rgb <= "000000";
					when "01110011100000111" => rgb <= "000000";
					when "01110011100001000" => rgb <= "000000";
					when "01110011100001001" => rgb <= "000000";
					when "01110011100001010" => rgb <= "000000";
					when "01110011100001011" => rgb <= "000000";
					when "01110011100001100" => rgb <= "000000";
					when "01110011100001101" => rgb <= "000000";
					when "01110011100001110" => rgb <= "000000";
					when "01110011100001111" => rgb <= "000000";
					when "01110011100010000" => rgb <= "000000";
					when "01110011100010001" => rgb <= "000000";
					when "01110011100010010" => rgb <= "000000";
					when "01110011100010011" => rgb <= "000000";
					when "01110011100010100" => rgb <= "000000";
					when "01110011100010101" => rgb <= "000000";
					when "01110011100010110" => rgb <= "000000";
					when "01110011100010111" => rgb <= "000000";
					when "01110011100011000" => rgb <= "000000";
					when "01110011100011001" => rgb <= "000000";
					when "01110011100011010" => rgb <= "000000";
					when "01110011100011011" => rgb <= "000000";
					when "01110011100011100" => rgb <= "000000";
					when "01110011100011101" => rgb <= "000000";
					when "01110011100011110" => rgb <= "000000";
					when "01110011100011111" => rgb <= "000000";
					when "01110011100100000" => rgb <= "000000";
					when "01110011100100001" => rgb <= "000000";
					when "01110011100100010" => rgb <= "000000";
					when "01110011100100011" => rgb <= "000000";
					when "01110011100100100" => rgb <= "000000";
					when "01110011100100101" => rgb <= "000000";
					when "01110011100100110" => rgb <= "000000";
					when "01110011100100111" => rgb <= "000000";
					when "01110011100101000" => rgb <= "000000";
					when "01110011100101001" => rgb <= "000000";
					when "01110011100101010" => rgb <= "000000";
					when "01110011100101011" => rgb <= "000000";
					when "01110011100101100" => rgb <= "000000";
					when "01110011100101101" => rgb <= "000000";
					when "01110011100101110" => rgb <= "000000";
					when "01110011100101111" => rgb <= "000000";
					when "01110011100110000" => rgb <= "000000";
					when "01110011100110001" => rgb <= "000000";
					when "01110011100110010" => rgb <= "000000";
					when "01110011100110011" => rgb <= "000000";
					when "01110011100110100" => rgb <= "000000";
					when "01110011100110101" => rgb <= "000000";
					when "01110011100110110" => rgb <= "000000";
					when "01110011100110111" => rgb <= "000000";
					when "01110011100111000" => rgb <= "000000";
					when "01110011100111001" => rgb <= "000000";
					when "01110011100111010" => rgb <= "000000";
					when "01110011100111011" => rgb <= "000000";
					when "01110011100111100" => rgb <= "000000";
					when "01110011100111101" => rgb <= "000000";
					when "01110011100111110" => rgb <= "000000";
					when "01110011100111111" => rgb <= "000000";
					when "01110100000000000" => rgb <= "000000";
					when "01110100000000001" => rgb <= "000000";
					when "01110100000000010" => rgb <= "000000";
					when "01110100000000011" => rgb <= "000000";
					when "01110100000000100" => rgb <= "000000";
					when "01110100000000101" => rgb <= "000000";
					when "01110100000000110" => rgb <= "000000";
					when "01110100000000111" => rgb <= "000000";
					when "01110100000001000" => rgb <= "000000";
					when "01110100000001001" => rgb <= "000000";
					when "01110100000001010" => rgb <= "000000";
					when "01110100000001011" => rgb <= "000000";
					when "01110100000001100" => rgb <= "000000";
					when "01110100000001101" => rgb <= "000000";
					when "01110100000001110" => rgb <= "000000";
					when "01110100000001111" => rgb <= "000000";
					when "01110100000010000" => rgb <= "000000";
					when "01110100000010001" => rgb <= "000000";
					when "01110100000010010" => rgb <= "000000";
					when "01110100000010011" => rgb <= "000000";
					when "01110100000010100" => rgb <= "000000";
					when "01110100000010101" => rgb <= "000000";
					when "01110100000010110" => rgb <= "000000";
					when "01110100000010111" => rgb <= "000000";
					when "01110100000011000" => rgb <= "000000";
					when "01110100000011001" => rgb <= "000000";
					when "01110100000011010" => rgb <= "000000";
					when "01110100000011011" => rgb <= "000000";
					when "01110100000011100" => rgb <= "000000";
					when "01110100000011101" => rgb <= "000000";
					when "01110100000011110" => rgb <= "000000";
					when "01110100000011111" => rgb <= "000000";
					when "01110100000100000" => rgb <= "000000";
					when "01110100000100001" => rgb <= "000000";
					when "01110100000100010" => rgb <= "000000";
					when "01110100000100011" => rgb <= "000000";
					when "01110100000100100" => rgb <= "000000";
					when "01110100000100101" => rgb <= "000000";
					when "01110100000100110" => rgb <= "000000";
					when "01110100000100111" => rgb <= "000000";
					when "01110100000101000" => rgb <= "000000";
					when "01110100000101001" => rgb <= "000000";
					when "01110100000101010" => rgb <= "000000";
					when "01110100000101011" => rgb <= "000000";
					when "01110100000101100" => rgb <= "000000";
					when "01110100000101101" => rgb <= "000000";
					when "01110100000101110" => rgb <= "000000";
					when "01110100000101111" => rgb <= "000000";
					when "01110100000110000" => rgb <= "000000";
					when "01110100000110001" => rgb <= "000000";
					when "01110100000110010" => rgb <= "000000";
					when "01110100000110011" => rgb <= "000000";
					when "01110100000110100" => rgb <= "000000";
					when "01110100000110101" => rgb <= "000000";
					when "01110100000110110" => rgb <= "000000";
					when "01110100000110111" => rgb <= "000000";
					when "01110100000111000" => rgb <= "000000";
					when "01110100000111001" => rgb <= "000000";
					when "01110100000111010" => rgb <= "000000";
					when "01110100000111011" => rgb <= "000000";
					when "01110100000111100" => rgb <= "000000";
					when "01110100000111101" => rgb <= "000000";
					when "01110100000111110" => rgb <= "000000";
					when "01110100000111111" => rgb <= "000000";
					when "01110100001000000" => rgb <= "000000";
					when "01110100001000001" => rgb <= "000000";
					when "01110100001000010" => rgb <= "000000";
					when "01110100001000011" => rgb <= "000000";
					when "01110100001000100" => rgb <= "000000";
					when "01110100001000101" => rgb <= "000000";
					when "01110100001000110" => rgb <= "000000";
					when "01110100001000111" => rgb <= "000000";
					when "01110100001001000" => rgb <= "000000";
					when "01110100001001001" => rgb <= "000000";
					when "01110100001001010" => rgb <= "000000";
					when "01110100001001011" => rgb <= "000000";
					when "01110100001001100" => rgb <= "000000";
					when "01110100001001101" => rgb <= "000000";
					when "01110100001001110" => rgb <= "000000";
					when "01110100001001111" => rgb <= "000000";
					when "01110100001010000" => rgb <= "000000";
					when "01110100001010001" => rgb <= "000000";
					when "01110100001010010" => rgb <= "000000";
					when "01110100001010011" => rgb <= "000000";
					when "01110100001010100" => rgb <= "000000";
					when "01110100001010101" => rgb <= "000000";
					when "01110100001010110" => rgb <= "000000";
					when "01110100001010111" => rgb <= "000000";
					when "01110100001011000" => rgb <= "000000";
					when "01110100001011001" => rgb <= "000000";
					when "01110100001011010" => rgb <= "000000";
					when "01110100001011011" => rgb <= "000000";
					when "01110100001011100" => rgb <= "000000";
					when "01110100001011101" => rgb <= "000000";
					when "01110100001011110" => rgb <= "000000";
					when "01110100001011111" => rgb <= "000000";
					when "01110100001100000" => rgb <= "000000";
					when "01110100001100001" => rgb <= "000000";
					when "01110100001100010" => rgb <= "000000";
					when "01110100001100011" => rgb <= "000000";
					when "01110100001100100" => rgb <= "000000";
					when "01110100001100101" => rgb <= "000000";
					when "01110100001100110" => rgb <= "000000";
					when "01110100001100111" => rgb <= "000000";
					when "01110100001101000" => rgb <= "000000";
					when "01110100001101001" => rgb <= "000000";
					when "01110100001101010" => rgb <= "000000";
					when "01110100001101011" => rgb <= "000000";
					when "01110100001101100" => rgb <= "000000";
					when "01110100001101101" => rgb <= "000000";
					when "01110100001101110" => rgb <= "000000";
					when "01110100001101111" => rgb <= "000000";
					when "01110100001110000" => rgb <= "000000";
					when "01110100001110001" => rgb <= "000000";
					when "01110100001110010" => rgb <= "000000";
					when "01110100001110011" => rgb <= "000000";
					when "01110100001110100" => rgb <= "000000";
					when "01110100001110101" => rgb <= "000000";
					when "01110100001110110" => rgb <= "000000";
					when "01110100001110111" => rgb <= "000000";
					when "01110100001111000" => rgb <= "000000";
					when "01110100001111001" => rgb <= "000000";
					when "01110100001111010" => rgb <= "000000";
					when "01110100001111011" => rgb <= "000000";
					when "01110100001111100" => rgb <= "000000";
					when "01110100001111101" => rgb <= "000000";
					when "01110100001111110" => rgb <= "000000";
					when "01110100001111111" => rgb <= "000000";
					when "01110100010000000" => rgb <= "000000";
					when "01110100010000001" => rgb <= "000000";
					when "01110100010000010" => rgb <= "000000";
					when "01110100010000011" => rgb <= "000000";
					when "01110100010000100" => rgb <= "000000";
					when "01110100010000101" => rgb <= "000000";
					when "01110100010000110" => rgb <= "000000";
					when "01110100010000111" => rgb <= "000000";
					when "01110100010001000" => rgb <= "010100";
					when "01110100010001001" => rgb <= "101000";
					when "01110100010001010" => rgb <= "101000";
					when "01110100010001011" => rgb <= "101000";
					when "01110100010001100" => rgb <= "101000";
					when "01110100010001101" => rgb <= "101000";
					when "01110100010001110" => rgb <= "101000";
					when "01110100010001111" => rgb <= "101000";
					when "01110100010010000" => rgb <= "101000";
					when "01110100010010001" => rgb <= "101000";
					when "01110100010010010" => rgb <= "101000";
					when "01110100010010011" => rgb <= "101000";
					when "01110100010010100" => rgb <= "101000";
					when "01110100010010101" => rgb <= "101000";
					when "01110100010010110" => rgb <= "101000";
					when "01110100010010111" => rgb <= "101000";
					when "01110100010011000" => rgb <= "101000";
					when "01110100010011001" => rgb <= "101000";
					when "01110100010011010" => rgb <= "101000";
					when "01110100010011011" => rgb <= "101000";
					when "01110100010011100" => rgb <= "101000";
					when "01110100010011101" => rgb <= "101000";
					when "01110100010011110" => rgb <= "101000";
					when "01110100010011111" => rgb <= "101000";
					when "01110100010100000" => rgb <= "101000";
					when "01110100010100001" => rgb <= "101000";
					when "01110100010100010" => rgb <= "101000";
					when "01110100010100011" => rgb <= "101000";
					when "01110100010100100" => rgb <= "101000";
					when "01110100010100101" => rgb <= "101000";
					when "01110100010100110" => rgb <= "101000";
					when "01110100010100111" => rgb <= "101000";
					when "01110100010101000" => rgb <= "101000";
					when "01110100010101001" => rgb <= "101000";
					when "01110100010101010" => rgb <= "101000";
					when "01110100010101011" => rgb <= "101000";
					when "01110100010101100" => rgb <= "101000";
					when "01110100010101101" => rgb <= "101000";
					when "01110100010101110" => rgb <= "101000";
					when "01110100010101111" => rgb <= "101000";
					when "01110100010110000" => rgb <= "101000";
					when "01110100010110001" => rgb <= "101000";
					when "01110100010110010" => rgb <= "101000";
					when "01110100010110011" => rgb <= "101000";
					when "01110100010110100" => rgb <= "101000";
					when "01110100010110101" => rgb <= "010100";
					when "01110100010110110" => rgb <= "000000";
					when "01110100010110111" => rgb <= "000000";
					when "01110100010111000" => rgb <= "000000";
					when "01110100010111001" => rgb <= "000000";
					when "01110100010111010" => rgb <= "000000";
					when "01110100010111011" => rgb <= "000000";
					when "01110100010111100" => rgb <= "000000";
					when "01110100010111101" => rgb <= "000000";
					when "01110100010111110" => rgb <= "000000";
					when "01110100010111111" => rgb <= "000000";
					when "01110100011000000" => rgb <= "000000";
					when "01110100011000001" => rgb <= "000000";
					when "01110100011000010" => rgb <= "000000";
					when "01110100011000011" => rgb <= "000000";
					when "01110100011000100" => rgb <= "000000";
					when "01110100011000101" => rgb <= "000000";
					when "01110100011000110" => rgb <= "000000";
					when "01110100011000111" => rgb <= "000000";
					when "01110100011001000" => rgb <= "000000";
					when "01110100011001001" => rgb <= "000000";
					when "01110100011001010" => rgb <= "000000";
					when "01110100011001011" => rgb <= "000000";
					when "01110100011001100" => rgb <= "000000";
					when "01110100011001101" => rgb <= "000000";
					when "01110100011001110" => rgb <= "000000";
					when "01110100011001111" => rgb <= "000000";
					when "01110100011010000" => rgb <= "000000";
					when "01110100011010001" => rgb <= "000000";
					when "01110100011010010" => rgb <= "000000";
					when "01110100011010011" => rgb <= "000000";
					when "01110100011010100" => rgb <= "000000";
					when "01110100011010101" => rgb <= "000000";
					when "01110100011010110" => rgb <= "000000";
					when "01110100011010111" => rgb <= "000000";
					when "01110100011011000" => rgb <= "000000";
					when "01110100011011001" => rgb <= "000000";
					when "01110100011011010" => rgb <= "000000";
					when "01110100011011011" => rgb <= "000000";
					when "01110100011011100" => rgb <= "000000";
					when "01110100011011101" => rgb <= "000000";
					when "01110100011011110" => rgb <= "000000";
					when "01110100011011111" => rgb <= "000000";
					when "01110100011100000" => rgb <= "000000";
					when "01110100011100001" => rgb <= "000000";
					when "01110100011100010" => rgb <= "000000";
					when "01110100011100011" => rgb <= "000000";
					when "01110100011100100" => rgb <= "000000";
					when "01110100011100101" => rgb <= "000000";
					when "01110100011100110" => rgb <= "000000";
					when "01110100011100111" => rgb <= "000000";
					when "01110100011101000" => rgb <= "000000";
					when "01110100011101001" => rgb <= "000000";
					when "01110100011101010" => rgb <= "000000";
					when "01110100011101011" => rgb <= "000000";
					when "01110100011101100" => rgb <= "000000";
					when "01110100011101101" => rgb <= "000000";
					when "01110100011101110" => rgb <= "000000";
					when "01110100011101111" => rgb <= "000000";
					when "01110100011110000" => rgb <= "000000";
					when "01110100011110001" => rgb <= "000000";
					when "01110100011110010" => rgb <= "000000";
					when "01110100011110011" => rgb <= "000000";
					when "01110100011110100" => rgb <= "000000";
					when "01110100011110101" => rgb <= "000000";
					when "01110100011110110" => rgb <= "000000";
					when "01110100011110111" => rgb <= "000000";
					when "01110100011111000" => rgb <= "000000";
					when "01110100011111001" => rgb <= "000000";
					when "01110100011111010" => rgb <= "000000";
					when "01110100011111011" => rgb <= "000000";
					when "01110100011111100" => rgb <= "000000";
					when "01110100011111101" => rgb <= "000000";
					when "01110100011111110" => rgb <= "000000";
					when "01110100011111111" => rgb <= "000000";
					when "01110100100000000" => rgb <= "000000";
					when "01110100100000001" => rgb <= "000000";
					when "01110100100000010" => rgb <= "000000";
					when "01110100100000011" => rgb <= "000000";
					when "01110100100000100" => rgb <= "000000";
					when "01110100100000101" => rgb <= "000000";
					when "01110100100000110" => rgb <= "000000";
					when "01110100100000111" => rgb <= "000000";
					when "01110100100001000" => rgb <= "000000";
					when "01110100100001001" => rgb <= "000000";
					when "01110100100001010" => rgb <= "000000";
					when "01110100100001011" => rgb <= "000000";
					when "01110100100001100" => rgb <= "000000";
					when "01110100100001101" => rgb <= "000000";
					when "01110100100001110" => rgb <= "000000";
					when "01110100100001111" => rgb <= "000000";
					when "01110100100010000" => rgb <= "000000";
					when "01110100100010001" => rgb <= "000000";
					when "01110100100010010" => rgb <= "000000";
					when "01110100100010011" => rgb <= "000000";
					when "01110100100010100" => rgb <= "000000";
					when "01110100100010101" => rgb <= "000000";
					when "01110100100010110" => rgb <= "000000";
					when "01110100100010111" => rgb <= "000000";
					when "01110100100011000" => rgb <= "000000";
					when "01110100100011001" => rgb <= "000000";
					when "01110100100011010" => rgb <= "000000";
					when "01110100100011011" => rgb <= "000000";
					when "01110100100011100" => rgb <= "000000";
					when "01110100100011101" => rgb <= "000000";
					when "01110100100011110" => rgb <= "000000";
					when "01110100100011111" => rgb <= "000000";
					when "01110100100100000" => rgb <= "000000";
					when "01110100100100001" => rgb <= "000000";
					when "01110100100100010" => rgb <= "000000";
					when "01110100100100011" => rgb <= "000000";
					when "01110100100100100" => rgb <= "000000";
					when "01110100100100101" => rgb <= "000000";
					when "01110100100100110" => rgb <= "000000";
					when "01110100100100111" => rgb <= "000000";
					when "01110100100101000" => rgb <= "000000";
					when "01110100100101001" => rgb <= "000000";
					when "01110100100101010" => rgb <= "000000";
					when "01110100100101011" => rgb <= "000000";
					when "01110100100101100" => rgb <= "000000";
					when "01110100100101101" => rgb <= "000000";
					when "01110100100101110" => rgb <= "000000";
					when "01110100100101111" => rgb <= "000000";
					when "01110100100110000" => rgb <= "000000";
					when "01110100100110001" => rgb <= "000000";
					when "01110100100110010" => rgb <= "000000";
					when "01110100100110011" => rgb <= "000000";
					when "01110100100110100" => rgb <= "000000";
					when "01110100100110101" => rgb <= "000000";
					when "01110100100110110" => rgb <= "000000";
					when "01110100100110111" => rgb <= "000000";
					when "01110100100111000" => rgb <= "000000";
					when "01110100100111001" => rgb <= "000000";
					when "01110100100111010" => rgb <= "000000";
					when "01110100100111011" => rgb <= "000000";
					when "01110100100111100" => rgb <= "000000";
					when "01110100100111101" => rgb <= "000000";
					when "01110100100111110" => rgb <= "000000";
					when "01110100100111111" => rgb <= "000000";
					when "01110101000000000" => rgb <= "000000";
					when "01110101000000001" => rgb <= "000000";
					when "01110101000000010" => rgb <= "000000";
					when "01110101000000011" => rgb <= "000000";
					when "01110101000000100" => rgb <= "000000";
					when "01110101000000101" => rgb <= "000000";
					when "01110101000000110" => rgb <= "000000";
					when "01110101000000111" => rgb <= "000000";
					when "01110101000001000" => rgb <= "000000";
					when "01110101000001001" => rgb <= "000000";
					when "01110101000001010" => rgb <= "000000";
					when "01110101000001011" => rgb <= "000000";
					when "01110101000001100" => rgb <= "000000";
					when "01110101000001101" => rgb <= "000000";
					when "01110101000001110" => rgb <= "000000";
					when "01110101000001111" => rgb <= "000000";
					when "01110101000010000" => rgb <= "000000";
					when "01110101000010001" => rgb <= "000000";
					when "01110101000010010" => rgb <= "000000";
					when "01110101000010011" => rgb <= "000000";
					when "01110101000010100" => rgb <= "000000";
					when "01110101000010101" => rgb <= "000000";
					when "01110101000010110" => rgb <= "000000";
					when "01110101000010111" => rgb <= "000000";
					when "01110101000011000" => rgb <= "000000";
					when "01110101000011001" => rgb <= "000000";
					when "01110101000011010" => rgb <= "000000";
					when "01110101000011011" => rgb <= "000000";
					when "01110101000011100" => rgb <= "000000";
					when "01110101000011101" => rgb <= "000000";
					when "01110101000011110" => rgb <= "000000";
					when "01110101000011111" => rgb <= "000000";
					when "01110101000100000" => rgb <= "000000";
					when "01110101000100001" => rgb <= "000000";
					when "01110101000100010" => rgb <= "000000";
					when "01110101000100011" => rgb <= "000000";
					when "01110101000100100" => rgb <= "000000";
					when "01110101000100101" => rgb <= "000000";
					when "01110101000100110" => rgb <= "000000";
					when "01110101000100111" => rgb <= "000000";
					when "01110101000101000" => rgb <= "000000";
					when "01110101000101001" => rgb <= "000000";
					when "01110101000101010" => rgb <= "000000";
					when "01110101000101011" => rgb <= "000000";
					when "01110101000101100" => rgb <= "000000";
					when "01110101000101101" => rgb <= "000000";
					when "01110101000101110" => rgb <= "000000";
					when "01110101000101111" => rgb <= "000000";
					when "01110101000110000" => rgb <= "000000";
					when "01110101000110001" => rgb <= "000000";
					when "01110101000110010" => rgb <= "000000";
					when "01110101000110011" => rgb <= "000000";
					when "01110101000110100" => rgb <= "000000";
					when "01110101000110101" => rgb <= "000000";
					when "01110101000110110" => rgb <= "000000";
					when "01110101000110111" => rgb <= "000000";
					when "01110101000111000" => rgb <= "000000";
					when "01110101000111001" => rgb <= "000000";
					when "01110101000111010" => rgb <= "000000";
					when "01110101000111011" => rgb <= "000000";
					when "01110101000111100" => rgb <= "000000";
					when "01110101000111101" => rgb <= "000000";
					when "01110101000111110" => rgb <= "000000";
					when "01110101000111111" => rgb <= "000000";
					when "01110101001000000" => rgb <= "000000";
					when "01110101001000001" => rgb <= "000000";
					when "01110101001000010" => rgb <= "000000";
					when "01110101001000011" => rgb <= "000000";
					when "01110101001000100" => rgb <= "000000";
					when "01110101001000101" => rgb <= "000000";
					when "01110101001000110" => rgb <= "000000";
					when "01110101001000111" => rgb <= "000000";
					when "01110101001001000" => rgb <= "000000";
					when "01110101001001001" => rgb <= "000000";
					when "01110101001001010" => rgb <= "000000";
					when "01110101001001011" => rgb <= "000000";
					when "01110101001001100" => rgb <= "000000";
					when "01110101001001101" => rgb <= "000000";
					when "01110101001001110" => rgb <= "000000";
					when "01110101001001111" => rgb <= "000000";
					when "01110101001010000" => rgb <= "000000";
					when "01110101001010001" => rgb <= "000000";
					when "01110101001010010" => rgb <= "000000";
					when "01110101001010011" => rgb <= "000000";
					when "01110101001010100" => rgb <= "000000";
					when "01110101001010101" => rgb <= "000000";
					when "01110101001010110" => rgb <= "000000";
					when "01110101001010111" => rgb <= "000000";
					when "01110101001011000" => rgb <= "000000";
					when "01110101001011001" => rgb <= "000000";
					when "01110101001011010" => rgb <= "000000";
					when "01110101001011011" => rgb <= "000000";
					when "01110101001011100" => rgb <= "000000";
					when "01110101001011101" => rgb <= "000000";
					when "01110101001011110" => rgb <= "000000";
					when "01110101001011111" => rgb <= "000000";
					when "01110101001100000" => rgb <= "000000";
					when "01110101001100001" => rgb <= "000000";
					when "01110101001100010" => rgb <= "000000";
					when "01110101001100011" => rgb <= "000000";
					when "01110101001100100" => rgb <= "000000";
					when "01110101001100101" => rgb <= "000000";
					when "01110101001100110" => rgb <= "000000";
					when "01110101001100111" => rgb <= "000000";
					when "01110101001101000" => rgb <= "000000";
					when "01110101001101001" => rgb <= "000000";
					when "01110101001101010" => rgb <= "000000";
					when "01110101001101011" => rgb <= "000000";
					when "01110101001101100" => rgb <= "000000";
					when "01110101001101101" => rgb <= "000000";
					when "01110101001101110" => rgb <= "000000";
					when "01110101001101111" => rgb <= "000000";
					when "01110101001110000" => rgb <= "000000";
					when "01110101001110001" => rgb <= "000000";
					when "01110101001110010" => rgb <= "000000";
					when "01110101001110011" => rgb <= "000000";
					when "01110101001110100" => rgb <= "000000";
					when "01110101001110101" => rgb <= "000000";
					when "01110101001110110" => rgb <= "000000";
					when "01110101001110111" => rgb <= "000000";
					when "01110101001111000" => rgb <= "000000";
					when "01110101001111001" => rgb <= "000000";
					when "01110101001111010" => rgb <= "000000";
					when "01110101001111011" => rgb <= "000000";
					when "01110101001111100" => rgb <= "000000";
					when "01110101001111101" => rgb <= "000000";
					when "01110101001111110" => rgb <= "000000";
					when "01110101001111111" => rgb <= "000000";
					when "01110101010000000" => rgb <= "000000";
					when "01110101010000001" => rgb <= "000000";
					when "01110101010000010" => rgb <= "000000";
					when "01110101010000011" => rgb <= "000000";
					when "01110101010000100" => rgb <= "000000";
					when "01110101010000101" => rgb <= "000000";
					when "01110101010000110" => rgb <= "000000";
					when "01110101010000111" => rgb <= "000000";
					when "01110101010001000" => rgb <= "010100";
					when "01110101010001001" => rgb <= "101000";
					when "01110101010001010" => rgb <= "101000";
					when "01110101010001011" => rgb <= "101000";
					when "01110101010001100" => rgb <= "101000";
					when "01110101010001101" => rgb <= "101000";
					when "01110101010001110" => rgb <= "101000";
					when "01110101010001111" => rgb <= "101000";
					when "01110101010010000" => rgb <= "101000";
					when "01110101010010001" => rgb <= "101000";
					when "01110101010010010" => rgb <= "101000";
					when "01110101010010011" => rgb <= "101000";
					when "01110101010010100" => rgb <= "101000";
					when "01110101010010101" => rgb <= "101000";
					when "01110101010010110" => rgb <= "101000";
					when "01110101010010111" => rgb <= "101000";
					when "01110101010011000" => rgb <= "101000";
					when "01110101010011001" => rgb <= "101000";
					when "01110101010011010" => rgb <= "101000";
					when "01110101010011011" => rgb <= "101000";
					when "01110101010011100" => rgb <= "101000";
					when "01110101010011101" => rgb <= "101000";
					when "01110101010011110" => rgb <= "101000";
					when "01110101010011111" => rgb <= "101000";
					when "01110101010100000" => rgb <= "101000";
					when "01110101010100001" => rgb <= "101000";
					when "01110101010100010" => rgb <= "101000";
					when "01110101010100011" => rgb <= "101000";
					when "01110101010100100" => rgb <= "101000";
					when "01110101010100101" => rgb <= "101000";
					when "01110101010100110" => rgb <= "101000";
					when "01110101010100111" => rgb <= "101000";
					when "01110101010101000" => rgb <= "101000";
					when "01110101010101001" => rgb <= "101000";
					when "01110101010101010" => rgb <= "101000";
					when "01110101010101011" => rgb <= "101000";
					when "01110101010101100" => rgb <= "101000";
					when "01110101010101101" => rgb <= "101000";
					when "01110101010101110" => rgb <= "101000";
					when "01110101010101111" => rgb <= "101000";
					when "01110101010110000" => rgb <= "101000";
					when "01110101010110001" => rgb <= "101000";
					when "01110101010110010" => rgb <= "101000";
					when "01110101010110011" => rgb <= "101000";
					when "01110101010110100" => rgb <= "101000";
					when "01110101010110101" => rgb <= "010100";
					when "01110101010110110" => rgb <= "000000";
					when "01110101010110111" => rgb <= "000000";
					when "01110101010111000" => rgb <= "000000";
					when "01110101010111001" => rgb <= "000000";
					when "01110101010111010" => rgb <= "000000";
					when "01110101010111011" => rgb <= "000000";
					when "01110101010111100" => rgb <= "000000";
					when "01110101010111101" => rgb <= "000000";
					when "01110101010111110" => rgb <= "000000";
					when "01110101010111111" => rgb <= "000000";
					when "01110101011000000" => rgb <= "000000";
					when "01110101011000001" => rgb <= "000000";
					when "01110101011000010" => rgb <= "000000";
					when "01110101011000011" => rgb <= "000000";
					when "01110101011000100" => rgb <= "000000";
					when "01110101011000101" => rgb <= "000000";
					when "01110101011000110" => rgb <= "000000";
					when "01110101011000111" => rgb <= "000000";
					when "01110101011001000" => rgb <= "000000";
					when "01110101011001001" => rgb <= "000000";
					when "01110101011001010" => rgb <= "000000";
					when "01110101011001011" => rgb <= "000000";
					when "01110101011001100" => rgb <= "000000";
					when "01110101011001101" => rgb <= "000000";
					when "01110101011001110" => rgb <= "000000";
					when "01110101011001111" => rgb <= "000000";
					when "01110101011010000" => rgb <= "000000";
					when "01110101011010001" => rgb <= "000000";
					when "01110101011010010" => rgb <= "000000";
					when "01110101011010011" => rgb <= "000000";
					when "01110101011010100" => rgb <= "000000";
					when "01110101011010101" => rgb <= "000000";
					when "01110101011010110" => rgb <= "000000";
					when "01110101011010111" => rgb <= "000000";
					when "01110101011011000" => rgb <= "000000";
					when "01110101011011001" => rgb <= "000000";
					when "01110101011011010" => rgb <= "000000";
					when "01110101011011011" => rgb <= "000000";
					when "01110101011011100" => rgb <= "000000";
					when "01110101011011101" => rgb <= "000000";
					when "01110101011011110" => rgb <= "000000";
					when "01110101011011111" => rgb <= "000000";
					when "01110101011100000" => rgb <= "000000";
					when "01110101011100001" => rgb <= "000000";
					when "01110101011100010" => rgb <= "000000";
					when "01110101011100011" => rgb <= "000000";
					when "01110101011100100" => rgb <= "000000";
					when "01110101011100101" => rgb <= "000000";
					when "01110101011100110" => rgb <= "000000";
					when "01110101011100111" => rgb <= "000000";
					when "01110101011101000" => rgb <= "000000";
					when "01110101011101001" => rgb <= "000000";
					when "01110101011101010" => rgb <= "000000";
					when "01110101011101011" => rgb <= "000000";
					when "01110101011101100" => rgb <= "000000";
					when "01110101011101101" => rgb <= "000000";
					when "01110101011101110" => rgb <= "000000";
					when "01110101011101111" => rgb <= "000000";
					when "01110101011110000" => rgb <= "000000";
					when "01110101011110001" => rgb <= "000000";
					when "01110101011110010" => rgb <= "000000";
					when "01110101011110011" => rgb <= "000000";
					when "01110101011110100" => rgb <= "000000";
					when "01110101011110101" => rgb <= "000000";
					when "01110101011110110" => rgb <= "000000";
					when "01110101011110111" => rgb <= "000000";
					when "01110101011111000" => rgb <= "000000";
					when "01110101011111001" => rgb <= "000000";
					when "01110101011111010" => rgb <= "000000";
					when "01110101011111011" => rgb <= "000000";
					when "01110101011111100" => rgb <= "000000";
					when "01110101011111101" => rgb <= "000000";
					when "01110101011111110" => rgb <= "000000";
					when "01110101011111111" => rgb <= "000000";
					when "01110101100000000" => rgb <= "000000";
					when "01110101100000001" => rgb <= "000000";
					when "01110101100000010" => rgb <= "000000";
					when "01110101100000011" => rgb <= "000000";
					when "01110101100000100" => rgb <= "000000";
					when "01110101100000101" => rgb <= "000000";
					when "01110101100000110" => rgb <= "000000";
					when "01110101100000111" => rgb <= "000000";
					when "01110101100001000" => rgb <= "000000";
					when "01110101100001001" => rgb <= "000000";
					when "01110101100001010" => rgb <= "000000";
					when "01110101100001011" => rgb <= "000000";
					when "01110101100001100" => rgb <= "000000";
					when "01110101100001101" => rgb <= "000000";
					when "01110101100001110" => rgb <= "000000";
					when "01110101100001111" => rgb <= "000000";
					when "01110101100010000" => rgb <= "000000";
					when "01110101100010001" => rgb <= "000000";
					when "01110101100010010" => rgb <= "000000";
					when "01110101100010011" => rgb <= "000000";
					when "01110101100010100" => rgb <= "000000";
					when "01110101100010101" => rgb <= "000000";
					when "01110101100010110" => rgb <= "000000";
					when "01110101100010111" => rgb <= "000000";
					when "01110101100011000" => rgb <= "000000";
					when "01110101100011001" => rgb <= "000000";
					when "01110101100011010" => rgb <= "000000";
					when "01110101100011011" => rgb <= "000000";
					when "01110101100011100" => rgb <= "000000";
					when "01110101100011101" => rgb <= "000000";
					when "01110101100011110" => rgb <= "000000";
					when "01110101100011111" => rgb <= "000000";
					when "01110101100100000" => rgb <= "000000";
					when "01110101100100001" => rgb <= "000000";
					when "01110101100100010" => rgb <= "000000";
					when "01110101100100011" => rgb <= "000000";
					when "01110101100100100" => rgb <= "000000";
					when "01110101100100101" => rgb <= "000000";
					when "01110101100100110" => rgb <= "000000";
					when "01110101100100111" => rgb <= "000000";
					when "01110101100101000" => rgb <= "000000";
					when "01110101100101001" => rgb <= "000000";
					when "01110101100101010" => rgb <= "000000";
					when "01110101100101011" => rgb <= "000000";
					when "01110101100101100" => rgb <= "000000";
					when "01110101100101101" => rgb <= "000000";
					when "01110101100101110" => rgb <= "000000";
					when "01110101100101111" => rgb <= "000000";
					when "01110101100110000" => rgb <= "000000";
					when "01110101100110001" => rgb <= "000000";
					when "01110101100110010" => rgb <= "000000";
					when "01110101100110011" => rgb <= "000000";
					when "01110101100110100" => rgb <= "000000";
					when "01110101100110101" => rgb <= "000000";
					when "01110101100110110" => rgb <= "000000";
					when "01110101100110111" => rgb <= "000000";
					when "01110101100111000" => rgb <= "000000";
					when "01110101100111001" => rgb <= "000000";
					when "01110101100111010" => rgb <= "000000";
					when "01110101100111011" => rgb <= "000000";
					when "01110101100111100" => rgb <= "000000";
					when "01110101100111101" => rgb <= "000000";
					when "01110101100111110" => rgb <= "000000";
					when "01110101100111111" => rgb <= "000000";
					when "01110110000000000" => rgb <= "000000";
					when "01110110000000001" => rgb <= "000000";
					when "01110110000000010" => rgb <= "000000";
					when "01110110000000011" => rgb <= "000000";
					when "01110110000000100" => rgb <= "000000";
					when "01110110000000101" => rgb <= "000000";
					when "01110110000000110" => rgb <= "000000";
					when "01110110000000111" => rgb <= "000000";
					when "01110110000001000" => rgb <= "000000";
					when "01110110000001001" => rgb <= "000000";
					when "01110110000001010" => rgb <= "000000";
					when "01110110000001011" => rgb <= "000000";
					when "01110110000001100" => rgb <= "000000";
					when "01110110000001101" => rgb <= "000000";
					when "01110110000001110" => rgb <= "000000";
					when "01110110000001111" => rgb <= "000000";
					when "01110110000010000" => rgb <= "000000";
					when "01110110000010001" => rgb <= "000000";
					when "01110110000010010" => rgb <= "000000";
					when "01110110000010011" => rgb <= "000000";
					when "01110110000010100" => rgb <= "000000";
					when "01110110000010101" => rgb <= "000000";
					when "01110110000010110" => rgb <= "000000";
					when "01110110000010111" => rgb <= "000000";
					when "01110110000011000" => rgb <= "000000";
					when "01110110000011001" => rgb <= "000000";
					when "01110110000011010" => rgb <= "000000";
					when "01110110000011011" => rgb <= "000000";
					when "01110110000011100" => rgb <= "000000";
					when "01110110000011101" => rgb <= "000000";
					when "01110110000011110" => rgb <= "000000";
					when "01110110000011111" => rgb <= "000000";
					when "01110110000100000" => rgb <= "000000";
					when "01110110000100001" => rgb <= "000000";
					when "01110110000100010" => rgb <= "000000";
					when "01110110000100011" => rgb <= "000000";
					when "01110110000100100" => rgb <= "000000";
					when "01110110000100101" => rgb <= "000000";
					when "01110110000100110" => rgb <= "000000";
					when "01110110000100111" => rgb <= "000000";
					when "01110110000101000" => rgb <= "000000";
					when "01110110000101001" => rgb <= "000000";
					when "01110110000101010" => rgb <= "000000";
					when "01110110000101011" => rgb <= "000000";
					when "01110110000101100" => rgb <= "000000";
					when "01110110000101101" => rgb <= "000000";
					when "01110110000101110" => rgb <= "000000";
					when "01110110000101111" => rgb <= "000000";
					when "01110110000110000" => rgb <= "000000";
					when "01110110000110001" => rgb <= "000000";
					when "01110110000110010" => rgb <= "000000";
					when "01110110000110011" => rgb <= "000000";
					when "01110110000110100" => rgb <= "000000";
					when "01110110000110101" => rgb <= "000000";
					when "01110110000110110" => rgb <= "000000";
					when "01110110000110111" => rgb <= "000000";
					when "01110110000111000" => rgb <= "000000";
					when "01110110000111001" => rgb <= "000000";
					when "01110110000111010" => rgb <= "000000";
					when "01110110000111011" => rgb <= "000000";
					when "01110110000111100" => rgb <= "000000";
					when "01110110000111101" => rgb <= "000000";
					when "01110110000111110" => rgb <= "000000";
					when "01110110000111111" => rgb <= "000000";
					when "01110110001000000" => rgb <= "000000";
					when "01110110001000001" => rgb <= "000000";
					when "01110110001000010" => rgb <= "000000";
					when "01110110001000011" => rgb <= "000000";
					when "01110110001000100" => rgb <= "000000";
					when "01110110001000101" => rgb <= "000000";
					when "01110110001000110" => rgb <= "000000";
					when "01110110001000111" => rgb <= "000000";
					when "01110110001001000" => rgb <= "000000";
					when "01110110001001001" => rgb <= "000000";
					when "01110110001001010" => rgb <= "000000";
					when "01110110001001011" => rgb <= "000000";
					when "01110110001001100" => rgb <= "000000";
					when "01110110001001101" => rgb <= "000000";
					when "01110110001001110" => rgb <= "000000";
					when "01110110001001111" => rgb <= "000000";
					when "01110110001010000" => rgb <= "000000";
					when "01110110001010001" => rgb <= "000000";
					when "01110110001010010" => rgb <= "000000";
					when "01110110001010011" => rgb <= "000000";
					when "01110110001010100" => rgb <= "000000";
					when "01110110001010101" => rgb <= "000000";
					when "01110110001010110" => rgb <= "000000";
					when "01110110001010111" => rgb <= "000000";
					when "01110110001011000" => rgb <= "000000";
					when "01110110001011001" => rgb <= "000000";
					when "01110110001011010" => rgb <= "000000";
					when "01110110001011011" => rgb <= "000000";
					when "01110110001011100" => rgb <= "000000";
					when "01110110001011101" => rgb <= "000000";
					when "01110110001011110" => rgb <= "000000";
					when "01110110001011111" => rgb <= "000000";
					when "01110110001100000" => rgb <= "000000";
					when "01110110001100001" => rgb <= "000000";
					when "01110110001100010" => rgb <= "000000";
					when "01110110001100011" => rgb <= "000000";
					when "01110110001100100" => rgb <= "000000";
					when "01110110001100101" => rgb <= "000000";
					when "01110110001100110" => rgb <= "000000";
					when "01110110001100111" => rgb <= "000000";
					when "01110110001101000" => rgb <= "000000";
					when "01110110001101001" => rgb <= "000000";
					when "01110110001101010" => rgb <= "000000";
					when "01110110001101011" => rgb <= "000000";
					when "01110110001101100" => rgb <= "000000";
					when "01110110001101101" => rgb <= "000000";
					when "01110110001101110" => rgb <= "000000";
					when "01110110001101111" => rgb <= "000000";
					when "01110110001110000" => rgb <= "000000";
					when "01110110001110001" => rgb <= "000000";
					when "01110110001110010" => rgb <= "000000";
					when "01110110001110011" => rgb <= "000000";
					when "01110110001110100" => rgb <= "000000";
					when "01110110001110101" => rgb <= "000000";
					when "01110110001110110" => rgb <= "000000";
					when "01110110001110111" => rgb <= "000000";
					when "01110110001111000" => rgb <= "000000";
					when "01110110001111001" => rgb <= "000000";
					when "01110110001111010" => rgb <= "000000";
					when "01110110001111011" => rgb <= "000000";
					when "01110110001111100" => rgb <= "000000";
					when "01110110001111101" => rgb <= "000000";
					when "01110110001111110" => rgb <= "000000";
					when "01110110001111111" => rgb <= "000000";
					when "01110110010000000" => rgb <= "000000";
					when "01110110010000001" => rgb <= "000000";
					when "01110110010000010" => rgb <= "000000";
					when "01110110010000011" => rgb <= "000000";
					when "01110110010000100" => rgb <= "000000";
					when "01110110010000101" => rgb <= "000000";
					when "01110110010000110" => rgb <= "000000";
					when "01110110010000111" => rgb <= "000000";
					when "01110110010001000" => rgb <= "010100";
					when "01110110010001001" => rgb <= "101000";
					when "01110110010001010" => rgb <= "101000";
					when "01110110010001011" => rgb <= "101000";
					when "01110110010001100" => rgb <= "101000";
					when "01110110010001101" => rgb <= "101000";
					when "01110110010001110" => rgb <= "101000";
					when "01110110010001111" => rgb <= "101000";
					when "01110110010010000" => rgb <= "101000";
					when "01110110010010001" => rgb <= "101000";
					when "01110110010010010" => rgb <= "101000";
					when "01110110010010011" => rgb <= "101000";
					when "01110110010010100" => rgb <= "101000";
					when "01110110010010101" => rgb <= "101000";
					when "01110110010010110" => rgb <= "101000";
					when "01110110010010111" => rgb <= "101000";
					when "01110110010011000" => rgb <= "101000";
					when "01110110010011001" => rgb <= "101000";
					when "01110110010011010" => rgb <= "101000";
					when "01110110010011011" => rgb <= "101000";
					when "01110110010011100" => rgb <= "101000";
					when "01110110010011101" => rgb <= "101000";
					when "01110110010011110" => rgb <= "101000";
					when "01110110010011111" => rgb <= "101000";
					when "01110110010100000" => rgb <= "101000";
					when "01110110010100001" => rgb <= "101000";
					when "01110110010100010" => rgb <= "101000";
					when "01110110010100011" => rgb <= "101000";
					when "01110110010100100" => rgb <= "101000";
					when "01110110010100101" => rgb <= "101000";
					when "01110110010100110" => rgb <= "101000";
					when "01110110010100111" => rgb <= "101000";
					when "01110110010101000" => rgb <= "101000";
					when "01110110010101001" => rgb <= "101000";
					when "01110110010101010" => rgb <= "101000";
					when "01110110010101011" => rgb <= "101000";
					when "01110110010101100" => rgb <= "101000";
					when "01110110010101101" => rgb <= "101000";
					when "01110110010101110" => rgb <= "101000";
					when "01110110010101111" => rgb <= "101000";
					when "01110110010110000" => rgb <= "101000";
					when "01110110010110001" => rgb <= "101000";
					when "01110110010110010" => rgb <= "101000";
					when "01110110010110011" => rgb <= "101000";
					when "01110110010110100" => rgb <= "101000";
					when "01110110010110101" => rgb <= "010100";
					when "01110110010110110" => rgb <= "000000";
					when "01110110010110111" => rgb <= "000000";
					when "01110110010111000" => rgb <= "000000";
					when "01110110010111001" => rgb <= "000000";
					when "01110110010111010" => rgb <= "000000";
					when "01110110010111011" => rgb <= "000000";
					when "01110110010111100" => rgb <= "000000";
					when "01110110010111101" => rgb <= "000000";
					when "01110110010111110" => rgb <= "000000";
					when "01110110010111111" => rgb <= "000000";
					when "01110110011000000" => rgb <= "000000";
					when "01110110011000001" => rgb <= "000000";
					when "01110110011000010" => rgb <= "000000";
					when "01110110011000011" => rgb <= "000000";
					when "01110110011000100" => rgb <= "000000";
					when "01110110011000101" => rgb <= "000000";
					when "01110110011000110" => rgb <= "000000";
					when "01110110011000111" => rgb <= "000000";
					when "01110110011001000" => rgb <= "000000";
					when "01110110011001001" => rgb <= "000000";
					when "01110110011001010" => rgb <= "000000";
					when "01110110011001011" => rgb <= "000000";
					when "01110110011001100" => rgb <= "000000";
					when "01110110011001101" => rgb <= "000000";
					when "01110110011001110" => rgb <= "000000";
					when "01110110011001111" => rgb <= "000000";
					when "01110110011010000" => rgb <= "000000";
					when "01110110011010001" => rgb <= "000000";
					when "01110110011010010" => rgb <= "000000";
					when "01110110011010011" => rgb <= "000000";
					when "01110110011010100" => rgb <= "000000";
					when "01110110011010101" => rgb <= "000000";
					when "01110110011010110" => rgb <= "000000";
					when "01110110011010111" => rgb <= "000000";
					when "01110110011011000" => rgb <= "000000";
					when "01110110011011001" => rgb <= "000000";
					when "01110110011011010" => rgb <= "000000";
					when "01110110011011011" => rgb <= "000000";
					when "01110110011011100" => rgb <= "000000";
					when "01110110011011101" => rgb <= "000000";
					when "01110110011011110" => rgb <= "000000";
					when "01110110011011111" => rgb <= "000000";
					when "01110110011100000" => rgb <= "000000";
					when "01110110011100001" => rgb <= "000000";
					when "01110110011100010" => rgb <= "000000";
					when "01110110011100011" => rgb <= "000000";
					when "01110110011100100" => rgb <= "000000";
					when "01110110011100101" => rgb <= "000000";
					when "01110110011100110" => rgb <= "000000";
					when "01110110011100111" => rgb <= "000000";
					when "01110110011101000" => rgb <= "000000";
					when "01110110011101001" => rgb <= "000000";
					when "01110110011101010" => rgb <= "000000";
					when "01110110011101011" => rgb <= "000000";
					when "01110110011101100" => rgb <= "000000";
					when "01110110011101101" => rgb <= "000000";
					when "01110110011101110" => rgb <= "000000";
					when "01110110011101111" => rgb <= "000000";
					when "01110110011110000" => rgb <= "000000";
					when "01110110011110001" => rgb <= "000000";
					when "01110110011110010" => rgb <= "000000";
					when "01110110011110011" => rgb <= "000000";
					when "01110110011110100" => rgb <= "000000";
					when "01110110011110101" => rgb <= "000000";
					when "01110110011110110" => rgb <= "000000";
					when "01110110011110111" => rgb <= "000000";
					when "01110110011111000" => rgb <= "000000";
					when "01110110011111001" => rgb <= "000000";
					when "01110110011111010" => rgb <= "000000";
					when "01110110011111011" => rgb <= "000000";
					when "01110110011111100" => rgb <= "000000";
					when "01110110011111101" => rgb <= "000000";
					when "01110110011111110" => rgb <= "000000";
					when "01110110011111111" => rgb <= "000000";
					when "01110110100000000" => rgb <= "000000";
					when "01110110100000001" => rgb <= "000000";
					when "01110110100000010" => rgb <= "000000";
					when "01110110100000011" => rgb <= "000000";
					when "01110110100000100" => rgb <= "000000";
					when "01110110100000101" => rgb <= "000000";
					when "01110110100000110" => rgb <= "000000";
					when "01110110100000111" => rgb <= "000000";
					when "01110110100001000" => rgb <= "000000";
					when "01110110100001001" => rgb <= "000000";
					when "01110110100001010" => rgb <= "000000";
					when "01110110100001011" => rgb <= "000000";
					when "01110110100001100" => rgb <= "000000";
					when "01110110100001101" => rgb <= "000000";
					when "01110110100001110" => rgb <= "000000";
					when "01110110100001111" => rgb <= "000000";
					when "01110110100010000" => rgb <= "000000";
					when "01110110100010001" => rgb <= "000000";
					when "01110110100010010" => rgb <= "000000";
					when "01110110100010011" => rgb <= "000000";
					when "01110110100010100" => rgb <= "000000";
					when "01110110100010101" => rgb <= "000000";
					when "01110110100010110" => rgb <= "000000";
					when "01110110100010111" => rgb <= "000000";
					when "01110110100011000" => rgb <= "000000";
					when "01110110100011001" => rgb <= "000000";
					when "01110110100011010" => rgb <= "000000";
					when "01110110100011011" => rgb <= "000000";
					when "01110110100011100" => rgb <= "000000";
					when "01110110100011101" => rgb <= "000000";
					when "01110110100011110" => rgb <= "000000";
					when "01110110100011111" => rgb <= "000000";
					when "01110110100100000" => rgb <= "000000";
					when "01110110100100001" => rgb <= "000000";
					when "01110110100100010" => rgb <= "000000";
					when "01110110100100011" => rgb <= "000000";
					when "01110110100100100" => rgb <= "000000";
					when "01110110100100101" => rgb <= "000000";
					when "01110110100100110" => rgb <= "000000";
					when "01110110100100111" => rgb <= "000000";
					when "01110110100101000" => rgb <= "000000";
					when "01110110100101001" => rgb <= "000000";
					when "01110110100101010" => rgb <= "000000";
					when "01110110100101011" => rgb <= "000000";
					when "01110110100101100" => rgb <= "000000";
					when "01110110100101101" => rgb <= "000000";
					when "01110110100101110" => rgb <= "000000";
					when "01110110100101111" => rgb <= "000000";
					when "01110110100110000" => rgb <= "000000";
					when "01110110100110001" => rgb <= "000000";
					when "01110110100110010" => rgb <= "000000";
					when "01110110100110011" => rgb <= "000000";
					when "01110110100110100" => rgb <= "000000";
					when "01110110100110101" => rgb <= "000000";
					when "01110110100110110" => rgb <= "000000";
					when "01110110100110111" => rgb <= "000000";
					when "01110110100111000" => rgb <= "000000";
					when "01110110100111001" => rgb <= "000000";
					when "01110110100111010" => rgb <= "000000";
					when "01110110100111011" => rgb <= "000000";
					when "01110110100111100" => rgb <= "000000";
					when "01110110100111101" => rgb <= "000000";
					when "01110110100111110" => rgb <= "000000";
					when "01110110100111111" => rgb <= "000000";
					when "01110111000000000" => rgb <= "000000";
					when "01110111000000001" => rgb <= "000000";
					when "01110111000000010" => rgb <= "000000";
					when "01110111000000011" => rgb <= "000000";
					when "01110111000000100" => rgb <= "000000";
					when "01110111000000101" => rgb <= "000000";
					when "01110111000000110" => rgb <= "000000";
					when "01110111000000111" => rgb <= "000000";
					when "01110111000001000" => rgb <= "000000";
					when "01110111000001001" => rgb <= "000000";
					when "01110111000001010" => rgb <= "000000";
					when "01110111000001011" => rgb <= "000000";
					when "01110111000001100" => rgb <= "000000";
					when "01110111000001101" => rgb <= "000000";
					when "01110111000001110" => rgb <= "000000";
					when "01110111000001111" => rgb <= "000000";
					when "01110111000010000" => rgb <= "000000";
					when "01110111000010001" => rgb <= "000000";
					when "01110111000010010" => rgb <= "000000";
					when "01110111000010011" => rgb <= "000000";
					when "01110111000010100" => rgb <= "000000";
					when "01110111000010101" => rgb <= "000000";
					when "01110111000010110" => rgb <= "000000";
					when "01110111000010111" => rgb <= "000000";
					when "01110111000011000" => rgb <= "000000";
					when "01110111000011001" => rgb <= "000000";
					when "01110111000011010" => rgb <= "000000";
					when "01110111000011011" => rgb <= "000000";
					when "01110111000011100" => rgb <= "000000";
					when "01110111000011101" => rgb <= "000000";
					when "01110111000011110" => rgb <= "000000";
					when "01110111000011111" => rgb <= "000000";
					when "01110111000100000" => rgb <= "000000";
					when "01110111000100001" => rgb <= "000000";
					when "01110111000100010" => rgb <= "000000";
					when "01110111000100011" => rgb <= "000000";
					when "01110111000100100" => rgb <= "000000";
					when "01110111000100101" => rgb <= "000000";
					when "01110111000100110" => rgb <= "000000";
					when "01110111000100111" => rgb <= "000000";
					when "01110111000101000" => rgb <= "000000";
					when "01110111000101001" => rgb <= "000000";
					when "01110111000101010" => rgb <= "000000";
					when "01110111000101011" => rgb <= "000000";
					when "01110111000101100" => rgb <= "000000";
					when "01110111000101101" => rgb <= "000000";
					when "01110111000101110" => rgb <= "000000";
					when "01110111000101111" => rgb <= "000000";
					when "01110111000110000" => rgb <= "000000";
					when "01110111000110001" => rgb <= "000000";
					when "01110111000110010" => rgb <= "000000";
					when "01110111000110011" => rgb <= "000000";
					when "01110111000110100" => rgb <= "000000";
					when "01110111000110101" => rgb <= "000000";
					when "01110111000110110" => rgb <= "000000";
					when "01110111000110111" => rgb <= "000000";
					when "01110111000111000" => rgb <= "000000";
					when "01110111000111001" => rgb <= "000000";
					when "01110111000111010" => rgb <= "000000";
					when "01110111000111011" => rgb <= "000000";
					when "01110111000111100" => rgb <= "000000";
					when "01110111000111101" => rgb <= "000000";
					when "01110111000111110" => rgb <= "000000";
					when "01110111000111111" => rgb <= "000000";
					when "01110111001000000" => rgb <= "000000";
					when "01110111001000001" => rgb <= "000000";
					when "01110111001000010" => rgb <= "000000";
					when "01110111001000011" => rgb <= "000000";
					when "01110111001000100" => rgb <= "000000";
					when "01110111001000101" => rgb <= "000000";
					when "01110111001000110" => rgb <= "000000";
					when "01110111001000111" => rgb <= "000000";
					when "01110111001001000" => rgb <= "000000";
					when "01110111001001001" => rgb <= "000000";
					when "01110111001001010" => rgb <= "000000";
					when "01110111001001011" => rgb <= "000000";
					when "01110111001001100" => rgb <= "000000";
					when "01110111001001101" => rgb <= "000000";
					when "01110111001001110" => rgb <= "000000";
					when "01110111001001111" => rgb <= "000000";
					when "01110111001010000" => rgb <= "000000";
					when "01110111001010001" => rgb <= "000000";
					when "01110111001010010" => rgb <= "000000";
					when "01110111001010011" => rgb <= "000000";
					when "01110111001010100" => rgb <= "000000";
					when "01110111001010101" => rgb <= "000000";
					when "01110111001010110" => rgb <= "000000";
					when "01110111001010111" => rgb <= "000000";
					when "01110111001011000" => rgb <= "000000";
					when "01110111001011001" => rgb <= "000000";
					when "01110111001011010" => rgb <= "000000";
					when "01110111001011011" => rgb <= "000000";
					when "01110111001011100" => rgb <= "000000";
					when "01110111001011101" => rgb <= "000000";
					when "01110111001011110" => rgb <= "000000";
					when "01110111001011111" => rgb <= "000000";
					when "01110111001100000" => rgb <= "000000";
					when "01110111001100001" => rgb <= "000000";
					when "01110111001100010" => rgb <= "000000";
					when "01110111001100011" => rgb <= "000000";
					when "01110111001100100" => rgb <= "000000";
					when "01110111001100101" => rgb <= "000000";
					when "01110111001100110" => rgb <= "000000";
					when "01110111001100111" => rgb <= "000000";
					when "01110111001101000" => rgb <= "000000";
					when "01110111001101001" => rgb <= "000000";
					when "01110111001101010" => rgb <= "000000";
					when "01110111001101011" => rgb <= "000000";
					when "01110111001101100" => rgb <= "000000";
					when "01110111001101101" => rgb <= "000000";
					when "01110111001101110" => rgb <= "000000";
					when "01110111001101111" => rgb <= "000000";
					when "01110111001110000" => rgb <= "000000";
					when "01110111001110001" => rgb <= "000000";
					when "01110111001110010" => rgb <= "000000";
					when "01110111001110011" => rgb <= "000000";
					when "01110111001110100" => rgb <= "000000";
					when "01110111001110101" => rgb <= "000000";
					when "01110111001110110" => rgb <= "000000";
					when "01110111001110111" => rgb <= "000000";
					when "01110111001111000" => rgb <= "000000";
					when "01110111001111001" => rgb <= "000000";
					when "01110111001111010" => rgb <= "000000";
					when "01110111001111011" => rgb <= "000000";
					when "01110111001111100" => rgb <= "000000";
					when "01110111001111101" => rgb <= "000000";
					when "01110111001111110" => rgb <= "000000";
					when "01110111001111111" => rgb <= "000000";
					when "01110111010000000" => rgb <= "000000";
					when "01110111010000001" => rgb <= "000000";
					when "01110111010000010" => rgb <= "000000";
					when "01110111010000011" => rgb <= "000000";
					when "01110111010000100" => rgb <= "000000";
					when "01110111010000101" => rgb <= "000000";
					when "01110111010000110" => rgb <= "000000";
					when "01110111010000111" => rgb <= "000000";
					when "01110111010001000" => rgb <= "000000";
					when "01110111010001001" => rgb <= "000000";
					when "01110111010001010" => rgb <= "000000";
					when "01110111010001011" => rgb <= "000000";
					when "01110111010001100" => rgb <= "000000";
					when "01110111010001101" => rgb <= "000000";
					when "01110111010001110" => rgb <= "000000";
					when "01110111010001111" => rgb <= "000000";
					when "01110111010010000" => rgb <= "000000";
					when "01110111010010001" => rgb <= "000000";
					when "01110111010010010" => rgb <= "000000";
					when "01110111010010011" => rgb <= "000000";
					when "01110111010010100" => rgb <= "000000";
					when "01110111010010101" => rgb <= "000000";
					when "01110111010010110" => rgb <= "000000";
					when "01110111010010111" => rgb <= "000000";
					when "01110111010011000" => rgb <= "000000";
					when "01110111010011001" => rgb <= "000000";
					when "01110111010011010" => rgb <= "000000";
					when "01110111010011011" => rgb <= "000000";
					when "01110111010011100" => rgb <= "000000";
					when "01110111010011101" => rgb <= "000000";
					when "01110111010011110" => rgb <= "000000";
					when "01110111010011111" => rgb <= "000000";
					when "01110111010100000" => rgb <= "000000";
					when "01110111010100001" => rgb <= "000000";
					when "01110111010100010" => rgb <= "000000";
					when "01110111010100011" => rgb <= "000000";
					when "01110111010100100" => rgb <= "000000";
					when "01110111010100101" => rgb <= "000000";
					when "01110111010100110" => rgb <= "000000";
					when "01110111010100111" => rgb <= "000000";
					when "01110111010101000" => rgb <= "000000";
					when "01110111010101001" => rgb <= "000000";
					when "01110111010101010" => rgb <= "000000";
					when "01110111010101011" => rgb <= "000000";
					when "01110111010101100" => rgb <= "000000";
					when "01110111010101101" => rgb <= "000000";
					when "01110111010101110" => rgb <= "000000";
					when "01110111010101111" => rgb <= "000000";
					when "01110111010110000" => rgb <= "000000";
					when "01110111010110001" => rgb <= "000000";
					when "01110111010110010" => rgb <= "000000";
					when "01110111010110011" => rgb <= "000000";
					when "01110111010110100" => rgb <= "000000";
					when "01110111010110101" => rgb <= "000000";
					when "01110111010110110" => rgb <= "000000";
					when "01110111010110111" => rgb <= "000000";
					when "01110111010111000" => rgb <= "000000";
					when "01110111010111001" => rgb <= "000000";
					when "01110111010111010" => rgb <= "000000";
					when "01110111010111011" => rgb <= "000000";
					when "01110111010111100" => rgb <= "000000";
					when "01110111010111101" => rgb <= "000000";
					when "01110111010111110" => rgb <= "000000";
					when "01110111010111111" => rgb <= "000000";
					when "01110111011000000" => rgb <= "000000";
					when "01110111011000001" => rgb <= "000000";
					when "01110111011000010" => rgb <= "000000";
					when "01110111011000011" => rgb <= "000000";
					when "01110111011000100" => rgb <= "000000";
					when "01110111011000101" => rgb <= "000000";
					when "01110111011000110" => rgb <= "000000";
					when "01110111011000111" => rgb <= "000000";
					when "01110111011001000" => rgb <= "000000";
					when "01110111011001001" => rgb <= "000000";
					when "01110111011001010" => rgb <= "000000";
					when "01110111011001011" => rgb <= "000000";
					when "01110111011001100" => rgb <= "000000";
					when "01110111011001101" => rgb <= "000000";
					when "01110111011001110" => rgb <= "000000";
					when "01110111011001111" => rgb <= "000000";
					when "01110111011010000" => rgb <= "000000";
					when "01110111011010001" => rgb <= "000000";
					when "01110111011010010" => rgb <= "000000";
					when "01110111011010011" => rgb <= "000000";
					when "01110111011010100" => rgb <= "000000";
					when "01110111011010101" => rgb <= "000000";
					when "01110111011010110" => rgb <= "000000";
					when "01110111011010111" => rgb <= "000000";
					when "01110111011011000" => rgb <= "000000";
					when "01110111011011001" => rgb <= "000000";
					when "01110111011011010" => rgb <= "000000";
					when "01110111011011011" => rgb <= "000000";
					when "01110111011011100" => rgb <= "000000";
					when "01110111011011101" => rgb <= "000000";
					when "01110111011011110" => rgb <= "000000";
					when "01110111011011111" => rgb <= "000000";
					when "01110111011100000" => rgb <= "000000";
					when "01110111011100001" => rgb <= "000000";
					when "01110111011100010" => rgb <= "000000";
					when "01110111011100011" => rgb <= "000000";
					when "01110111011100100" => rgb <= "000000";
					when "01110111011100101" => rgb <= "000000";
					when "01110111011100110" => rgb <= "000000";
					when "01110111011100111" => rgb <= "000000";
					when "01110111011101000" => rgb <= "000000";
					when "01110111011101001" => rgb <= "000000";
					when "01110111011101010" => rgb <= "000000";
					when "01110111011101011" => rgb <= "000000";
					when "01110111011101100" => rgb <= "000000";
					when "01110111011101101" => rgb <= "000000";
					when "01110111011101110" => rgb <= "000000";
					when "01110111011101111" => rgb <= "000000";
					when "01110111011110000" => rgb <= "000000";
					when "01110111011110001" => rgb <= "000000";
					when "01110111011110010" => rgb <= "000000";
					when "01110111011110011" => rgb <= "000000";
					when "01110111011110100" => rgb <= "000000";
					when "01110111011110101" => rgb <= "000000";
					when "01110111011110110" => rgb <= "000000";
					when "01110111011110111" => rgb <= "000000";
					when "01110111011111000" => rgb <= "000000";
					when "01110111011111001" => rgb <= "000000";
					when "01110111011111010" => rgb <= "000000";
					when "01110111011111011" => rgb <= "000000";
					when "01110111011111100" => rgb <= "000000";
					when "01110111011111101" => rgb <= "000000";
					when "01110111011111110" => rgb <= "000000";
					when "01110111011111111" => rgb <= "000000";
					when "01110111100000000" => rgb <= "000000";
					when "01110111100000001" => rgb <= "000000";
					when "01110111100000010" => rgb <= "000000";
					when "01110111100000011" => rgb <= "000000";
					when "01110111100000100" => rgb <= "000000";
					when "01110111100000101" => rgb <= "000000";
					when "01110111100000110" => rgb <= "000000";
					when "01110111100000111" => rgb <= "000000";
					when "01110111100001000" => rgb <= "000000";
					when "01110111100001001" => rgb <= "000000";
					when "01110111100001010" => rgb <= "000000";
					when "01110111100001011" => rgb <= "000000";
					when "01110111100001100" => rgb <= "000000";
					when "01110111100001101" => rgb <= "000000";
					when "01110111100001110" => rgb <= "000000";
					when "01110111100001111" => rgb <= "000000";
					when "01110111100010000" => rgb <= "000000";
					when "01110111100010001" => rgb <= "000000";
					when "01110111100010010" => rgb <= "000000";
					when "01110111100010011" => rgb <= "000000";
					when "01110111100010100" => rgb <= "000000";
					when "01110111100010101" => rgb <= "000000";
					when "01110111100010110" => rgb <= "000000";
					when "01110111100010111" => rgb <= "000000";
					when "01110111100011000" => rgb <= "000000";
					when "01110111100011001" => rgb <= "000000";
					when "01110111100011010" => rgb <= "000000";
					when "01110111100011011" => rgb <= "000000";
					when "01110111100011100" => rgb <= "000000";
					when "01110111100011101" => rgb <= "000000";
					when "01110111100011110" => rgb <= "000000";
					when "01110111100011111" => rgb <= "000000";
					when "01110111100100000" => rgb <= "000000";
					when "01110111100100001" => rgb <= "000000";
					when "01110111100100010" => rgb <= "000000";
					when "01110111100100011" => rgb <= "000000";
					when "01110111100100100" => rgb <= "000000";
					when "01110111100100101" => rgb <= "000000";
					when "01110111100100110" => rgb <= "000000";
					when "01110111100100111" => rgb <= "000000";
					when "01110111100101000" => rgb <= "000000";
					when "01110111100101001" => rgb <= "000000";
					when "01110111100101010" => rgb <= "000000";
					when "01110111100101011" => rgb <= "000000";
					when "01110111100101100" => rgb <= "000000";
					when "01110111100101101" => rgb <= "000000";
					when "01110111100101110" => rgb <= "000000";
					when "01110111100101111" => rgb <= "000000";
					when "01110111100110000" => rgb <= "000000";
					when "01110111100110001" => rgb <= "000000";
					when "01110111100110010" => rgb <= "000000";
					when "01110111100110011" => rgb <= "000000";
					when "01110111100110100" => rgb <= "000000";
					when "01110111100110101" => rgb <= "000000";
					when "01110111100110110" => rgb <= "000000";
					when "01110111100110111" => rgb <= "000000";
					when "01110111100111000" => rgb <= "000000";
					when "01110111100111001" => rgb <= "000000";
					when "01110111100111010" => rgb <= "000000";
					when "01110111100111011" => rgb <= "000000";
					when "01110111100111100" => rgb <= "000000";
					when "01110111100111101" => rgb <= "000000";
					when "01110111100111110" => rgb <= "000000";
					when "01110111100111111" => rgb <= "000000";
					when "01111000000000000" => rgb <= "000000";
					when "01111000000000001" => rgb <= "000000";
					when "01111000000000010" => rgb <= "000000";
					when "01111000000000011" => rgb <= "000000";
					when "01111000000000100" => rgb <= "000000";
					when "01111000000000101" => rgb <= "000000";
					when "01111000000000110" => rgb <= "000000";
					when "01111000000000111" => rgb <= "000000";
					when "01111000000001000" => rgb <= "000000";
					when "01111000000001001" => rgb <= "000000";
					when "01111000000001010" => rgb <= "000000";
					when "01111000000001011" => rgb <= "000000";
					when "01111000000001100" => rgb <= "000000";
					when "01111000000001101" => rgb <= "000000";
					when "01111000000001110" => rgb <= "000000";
					when "01111000000001111" => rgb <= "000000";
					when "01111000000010000" => rgb <= "000000";
					when "01111000000010001" => rgb <= "000000";
					when "01111000000010010" => rgb <= "000000";
					when "01111000000010011" => rgb <= "000000";
					when "01111000000010100" => rgb <= "000000";
					when "01111000000010101" => rgb <= "000000";
					when "01111000000010110" => rgb <= "000000";
					when "01111000000010111" => rgb <= "000000";
					when "01111000000011000" => rgb <= "000000";
					when "01111000000011001" => rgb <= "000000";
					when "01111000000011010" => rgb <= "000000";
					when "01111000000011011" => rgb <= "000000";
					when "01111000000011100" => rgb <= "000000";
					when "01111000000011101" => rgb <= "000000";
					when "01111000000011110" => rgb <= "000000";
					when "01111000000011111" => rgb <= "000000";
					when "01111000000100000" => rgb <= "000000";
					when "01111000000100001" => rgb <= "000000";
					when "01111000000100010" => rgb <= "000000";
					when "01111000000100011" => rgb <= "000000";
					when "01111000000100100" => rgb <= "000000";
					when "01111000000100101" => rgb <= "000000";
					when "01111000000100110" => rgb <= "000000";
					when "01111000000100111" => rgb <= "000000";
					when "01111000000101000" => rgb <= "000000";
					when "01111000000101001" => rgb <= "000000";
					when "01111000000101010" => rgb <= "000000";
					when "01111000000101011" => rgb <= "000000";
					when "01111000000101100" => rgb <= "000000";
					when "01111000000101101" => rgb <= "000000";
					when "01111000000101110" => rgb <= "000000";
					when "01111000000101111" => rgb <= "000000";
					when "01111000000110000" => rgb <= "000000";
					when "01111000000110001" => rgb <= "000000";
					when "01111000000110010" => rgb <= "000000";
					when "01111000000110011" => rgb <= "000000";
					when "01111000000110100" => rgb <= "000000";
					when "01111000000110101" => rgb <= "000000";
					when "01111000000110110" => rgb <= "000000";
					when "01111000000110111" => rgb <= "000000";
					when "01111000000111000" => rgb <= "000000";
					when "01111000000111001" => rgb <= "000000";
					when "01111000000111010" => rgb <= "000000";
					when "01111000000111011" => rgb <= "000000";
					when "01111000000111100" => rgb <= "000000";
					when "01111000000111101" => rgb <= "000000";
					when "01111000000111110" => rgb <= "000000";
					when "01111000000111111" => rgb <= "000000";
					when "01111000001000000" => rgb <= "000000";
					when "01111000001000001" => rgb <= "000000";
					when "01111000001000010" => rgb <= "000000";
					when "01111000001000011" => rgb <= "000000";
					when "01111000001000100" => rgb <= "000000";
					when "01111000001000101" => rgb <= "000000";
					when "01111000001000110" => rgb <= "000000";
					when "01111000001000111" => rgb <= "000000";
					when "01111000001001000" => rgb <= "000000";
					when "01111000001001001" => rgb <= "000000";
					when "01111000001001010" => rgb <= "000000";
					when "01111000001001011" => rgb <= "000000";
					when "01111000001001100" => rgb <= "000000";
					when "01111000001001101" => rgb <= "000000";
					when "01111000001001110" => rgb <= "000000";
					when "01111000001001111" => rgb <= "000000";
					when "01111000001010000" => rgb <= "000000";
					when "01111000001010001" => rgb <= "000000";
					when "01111000001010010" => rgb <= "000000";
					when "01111000001010011" => rgb <= "000000";
					when "01111000001010100" => rgb <= "000000";
					when "01111000001010101" => rgb <= "000000";
					when "01111000001010110" => rgb <= "000000";
					when "01111000001010111" => rgb <= "000000";
					when "01111000001011000" => rgb <= "000000";
					when "01111000001011001" => rgb <= "000000";
					when "01111000001011010" => rgb <= "000000";
					when "01111000001011011" => rgb <= "000000";
					when "01111000001011100" => rgb <= "000000";
					when "01111000001011101" => rgb <= "000000";
					when "01111000001011110" => rgb <= "000000";
					when "01111000001011111" => rgb <= "000000";
					when "01111000001100000" => rgb <= "000000";
					when "01111000001100001" => rgb <= "000000";
					when "01111000001100010" => rgb <= "000000";
					when "01111000001100011" => rgb <= "000000";
					when "01111000001100100" => rgb <= "000000";
					when "01111000001100101" => rgb <= "000000";
					when "01111000001100110" => rgb <= "000000";
					when "01111000001100111" => rgb <= "000000";
					when "01111000001101000" => rgb <= "000000";
					when "01111000001101001" => rgb <= "000000";
					when "01111000001101010" => rgb <= "000000";
					when "01111000001101011" => rgb <= "000000";
					when "01111000001101100" => rgb <= "000000";
					when "01111000001101101" => rgb <= "000000";
					when "01111000001101110" => rgb <= "000000";
					when "01111000001101111" => rgb <= "000000";
					when "01111000001110000" => rgb <= "000000";
					when "01111000001110001" => rgb <= "000000";
					when "01111000001110010" => rgb <= "000000";
					when "01111000001110011" => rgb <= "000000";
					when "01111000001110100" => rgb <= "000000";
					when "01111000001110101" => rgb <= "000000";
					when "01111000001110110" => rgb <= "000000";
					when "01111000001110111" => rgb <= "000000";
					when "01111000001111000" => rgb <= "000000";
					when "01111000001111001" => rgb <= "000000";
					when "01111000001111010" => rgb <= "000000";
					when "01111000001111011" => rgb <= "000000";
					when "01111000001111100" => rgb <= "000000";
					when "01111000001111101" => rgb <= "000000";
					when "01111000001111110" => rgb <= "000000";
					when "01111000001111111" => rgb <= "000000";
					when "01111000010000000" => rgb <= "000000";
					when "01111000010000001" => rgb <= "000000";
					when "01111000010000010" => rgb <= "000000";
					when "01111000010000011" => rgb <= "000000";
					when "01111000010000100" => rgb <= "000000";
					when "01111000010000101" => rgb <= "000000";
					when "01111000010000110" => rgb <= "000000";
					when "01111000010000111" => rgb <= "000000";
					when "01111000010001000" => rgb <= "000000";
					when "01111000010001001" => rgb <= "000000";
					when "01111000010001010" => rgb <= "000000";
					when "01111000010001011" => rgb <= "000000";
					when "01111000010001100" => rgb <= "000000";
					when "01111000010001101" => rgb <= "000000";
					when "01111000010001110" => rgb <= "000000";
					when "01111000010001111" => rgb <= "000000";
					when "01111000010010000" => rgb <= "000000";
					when "01111000010010001" => rgb <= "000000";
					when "01111000010010010" => rgb <= "000000";
					when "01111000010010011" => rgb <= "000000";
					when "01111000010010100" => rgb <= "000000";
					when "01111000010010101" => rgb <= "000000";
					when "01111000010010110" => rgb <= "000000";
					when "01111000010010111" => rgb <= "000000";
					when "01111000010011000" => rgb <= "000000";
					when "01111000010011001" => rgb <= "000000";
					when "01111000010011010" => rgb <= "000000";
					when "01111000010011011" => rgb <= "000000";
					when "01111000010011100" => rgb <= "000000";
					when "01111000010011101" => rgb <= "000000";
					when "01111000010011110" => rgb <= "000000";
					when "01111000010011111" => rgb <= "000000";
					when "01111000010100000" => rgb <= "000000";
					when "01111000010100001" => rgb <= "000000";
					when "01111000010100010" => rgb <= "000000";
					when "01111000010100011" => rgb <= "000000";
					when "01111000010100100" => rgb <= "000000";
					when "01111000010100101" => rgb <= "000000";
					when "01111000010100110" => rgb <= "000000";
					when "01111000010100111" => rgb <= "000000";
					when "01111000010101000" => rgb <= "000000";
					when "01111000010101001" => rgb <= "000000";
					when "01111000010101010" => rgb <= "000000";
					when "01111000010101011" => rgb <= "000000";
					when "01111000010101100" => rgb <= "000000";
					when "01111000010101101" => rgb <= "000000";
					when "01111000010101110" => rgb <= "000000";
					when "01111000010101111" => rgb <= "000000";
					when "01111000010110000" => rgb <= "000000";
					when "01111000010110001" => rgb <= "000000";
					when "01111000010110010" => rgb <= "000000";
					when "01111000010110011" => rgb <= "000000";
					when "01111000010110100" => rgb <= "000000";
					when "01111000010110101" => rgb <= "000000";
					when "01111000010110110" => rgb <= "000000";
					when "01111000010110111" => rgb <= "000000";
					when "01111000010111000" => rgb <= "000000";
					when "01111000010111001" => rgb <= "000000";
					when "01111000010111010" => rgb <= "000000";
					when "01111000010111011" => rgb <= "000000";
					when "01111000010111100" => rgb <= "000000";
					when "01111000010111101" => rgb <= "000000";
					when "01111000010111110" => rgb <= "000000";
					when "01111000010111111" => rgb <= "000000";
					when "01111000011000000" => rgb <= "000000";
					when "01111000011000001" => rgb <= "000000";
					when "01111000011000010" => rgb <= "000000";
					when "01111000011000011" => rgb <= "000000";
					when "01111000011000100" => rgb <= "000000";
					when "01111000011000101" => rgb <= "000000";
					when "01111000011000110" => rgb <= "000000";
					when "01111000011000111" => rgb <= "000000";
					when "01111000011001000" => rgb <= "000000";
					when "01111000011001001" => rgb <= "000000";
					when "01111000011001010" => rgb <= "000000";
					when "01111000011001011" => rgb <= "000000";
					when "01111000011001100" => rgb <= "000000";
					when "01111000011001101" => rgb <= "000000";
					when "01111000011001110" => rgb <= "000000";
					when "01111000011001111" => rgb <= "000000";
					when "01111000011010000" => rgb <= "000000";
					when "01111000011010001" => rgb <= "000000";
					when "01111000011010010" => rgb <= "000000";
					when "01111000011010011" => rgb <= "000000";
					when "01111000011010100" => rgb <= "000000";
					when "01111000011010101" => rgb <= "000000";
					when "01111000011010110" => rgb <= "000000";
					when "01111000011010111" => rgb <= "000000";
					when "01111000011011000" => rgb <= "000000";
					when "01111000011011001" => rgb <= "000000";
					when "01111000011011010" => rgb <= "000000";
					when "01111000011011011" => rgb <= "000000";
					when "01111000011011100" => rgb <= "000000";
					when "01111000011011101" => rgb <= "000000";
					when "01111000011011110" => rgb <= "000000";
					when "01111000011011111" => rgb <= "000000";
					when "01111000011100000" => rgb <= "000000";
					when "01111000011100001" => rgb <= "000000";
					when "01111000011100010" => rgb <= "000000";
					when "01111000011100011" => rgb <= "000000";
					when "01111000011100100" => rgb <= "000000";
					when "01111000011100101" => rgb <= "000000";
					when "01111000011100110" => rgb <= "000000";
					when "01111000011100111" => rgb <= "000000";
					when "01111000011101000" => rgb <= "000000";
					when "01111000011101001" => rgb <= "000000";
					when "01111000011101010" => rgb <= "000000";
					when "01111000011101011" => rgb <= "000000";
					when "01111000011101100" => rgb <= "000000";
					when "01111000011101101" => rgb <= "000000";
					when "01111000011101110" => rgb <= "000000";
					when "01111000011101111" => rgb <= "000000";
					when "01111000011110000" => rgb <= "000000";
					when "01111000011110001" => rgb <= "000000";
					when "01111000011110010" => rgb <= "000000";
					when "01111000011110011" => rgb <= "000000";
					when "01111000011110100" => rgb <= "000000";
					when "01111000011110101" => rgb <= "000000";
					when "01111000011110110" => rgb <= "000000";
					when "01111000011110111" => rgb <= "000000";
					when "01111000011111000" => rgb <= "000000";
					when "01111000011111001" => rgb <= "000000";
					when "01111000011111010" => rgb <= "000000";
					when "01111000011111011" => rgb <= "000000";
					when "01111000011111100" => rgb <= "000000";
					when "01111000011111101" => rgb <= "000000";
					when "01111000011111110" => rgb <= "000000";
					when "01111000011111111" => rgb <= "000000";
					when "01111000100000000" => rgb <= "000000";
					when "01111000100000001" => rgb <= "000000";
					when "01111000100000010" => rgb <= "000000";
					when "01111000100000011" => rgb <= "000000";
					when "01111000100000100" => rgb <= "000000";
					when "01111000100000101" => rgb <= "000000";
					when "01111000100000110" => rgb <= "000000";
					when "01111000100000111" => rgb <= "000000";
					when "01111000100001000" => rgb <= "000000";
					when "01111000100001001" => rgb <= "000000";
					when "01111000100001010" => rgb <= "000000";
					when "01111000100001011" => rgb <= "000000";
					when "01111000100001100" => rgb <= "000000";
					when "01111000100001101" => rgb <= "000000";
					when "01111000100001110" => rgb <= "000000";
					when "01111000100001111" => rgb <= "000000";
					when "01111000100010000" => rgb <= "000000";
					when "01111000100010001" => rgb <= "000000";
					when "01111000100010010" => rgb <= "000000";
					when "01111000100010011" => rgb <= "000000";
					when "01111000100010100" => rgb <= "000000";
					when "01111000100010101" => rgb <= "000000";
					when "01111000100010110" => rgb <= "000000";
					when "01111000100010111" => rgb <= "000000";
					when "01111000100011000" => rgb <= "000000";
					when "01111000100011001" => rgb <= "000000";
					when "01111000100011010" => rgb <= "000000";
					when "01111000100011011" => rgb <= "000000";
					when "01111000100011100" => rgb <= "000000";
					when "01111000100011101" => rgb <= "000000";
					when "01111000100011110" => rgb <= "000000";
					when "01111000100011111" => rgb <= "000000";
					when "01111000100100000" => rgb <= "000000";
					when "01111000100100001" => rgb <= "000000";
					when "01111000100100010" => rgb <= "000000";
					when "01111000100100011" => rgb <= "000000";
					when "01111000100100100" => rgb <= "000000";
					when "01111000100100101" => rgb <= "000000";
					when "01111000100100110" => rgb <= "000000";
					when "01111000100100111" => rgb <= "000000";
					when "01111000100101000" => rgb <= "000000";
					when "01111000100101001" => rgb <= "000000";
					when "01111000100101010" => rgb <= "000000";
					when "01111000100101011" => rgb <= "000000";
					when "01111000100101100" => rgb <= "000000";
					when "01111000100101101" => rgb <= "000000";
					when "01111000100101110" => rgb <= "000000";
					when "01111000100101111" => rgb <= "000000";
					when "01111000100110000" => rgb <= "000000";
					when "01111000100110001" => rgb <= "000000";
					when "01111000100110010" => rgb <= "000000";
					when "01111000100110011" => rgb <= "000000";
					when "01111000100110100" => rgb <= "000000";
					when "01111000100110101" => rgb <= "000000";
					when "01111000100110110" => rgb <= "000000";
					when "01111000100110111" => rgb <= "000000";
					when "01111000100111000" => rgb <= "000000";
					when "01111000100111001" => rgb <= "000000";
					when "01111000100111010" => rgb <= "000000";
					when "01111000100111011" => rgb <= "000000";
					when "01111000100111100" => rgb <= "000000";
					when "01111000100111101" => rgb <= "000000";
					when "01111000100111110" => rgb <= "000000";
					when "01111000100111111" => rgb <= "000000";
					when "01111001000000000" => rgb <= "000000";
					when "01111001000000001" => rgb <= "000000";
					when "01111001000000010" => rgb <= "000000";
					when "01111001000000011" => rgb <= "000000";
					when "01111001000000100" => rgb <= "000000";
					when "01111001000000101" => rgb <= "000000";
					when "01111001000000110" => rgb <= "000000";
					when "01111001000000111" => rgb <= "000000";
					when "01111001000001000" => rgb <= "000000";
					when "01111001000001001" => rgb <= "000000";
					when "01111001000001010" => rgb <= "000000";
					when "01111001000001011" => rgb <= "000000";
					when "01111001000001100" => rgb <= "000000";
					when "01111001000001101" => rgb <= "000000";
					when "01111001000001110" => rgb <= "000000";
					when "01111001000001111" => rgb <= "000000";
					when "01111001000010000" => rgb <= "000000";
					when "01111001000010001" => rgb <= "000000";
					when "01111001000010010" => rgb <= "000000";
					when "01111001000010011" => rgb <= "000000";
					when "01111001000010100" => rgb <= "000000";
					when "01111001000010101" => rgb <= "000000";
					when "01111001000010110" => rgb <= "000000";
					when "01111001000010111" => rgb <= "000000";
					when "01111001000011000" => rgb <= "000000";
					when "01111001000011001" => rgb <= "000000";
					when "01111001000011010" => rgb <= "000000";
					when "01111001000011011" => rgb <= "000000";
					when "01111001000011100" => rgb <= "000000";
					when "01111001000011101" => rgb <= "000000";
					when "01111001000011110" => rgb <= "000000";
					when "01111001000011111" => rgb <= "000000";
					when "01111001000100000" => rgb <= "000000";
					when "01111001000100001" => rgb <= "000000";
					when "01111001000100010" => rgb <= "000000";
					when "01111001000100011" => rgb <= "000000";
					when "01111001000100100" => rgb <= "000000";
					when "01111001000100101" => rgb <= "000000";
					when "01111001000100110" => rgb <= "000000";
					when "01111001000100111" => rgb <= "000000";
					when "01111001000101000" => rgb <= "000000";
					when "01111001000101001" => rgb <= "000000";
					when "01111001000101010" => rgb <= "000000";
					when "01111001000101011" => rgb <= "000000";
					when "01111001000101100" => rgb <= "000000";
					when "01111001000101101" => rgb <= "000000";
					when "01111001000101110" => rgb <= "000000";
					when "01111001000101111" => rgb <= "000000";
					when "01111001000110000" => rgb <= "000000";
					when "01111001000110001" => rgb <= "000000";
					when "01111001000110010" => rgb <= "000000";
					when "01111001000110011" => rgb <= "000000";
					when "01111001000110100" => rgb <= "000000";
					when "01111001000110101" => rgb <= "000000";
					when "01111001000110110" => rgb <= "000000";
					when "01111001000110111" => rgb <= "000000";
					when "01111001000111000" => rgb <= "000000";
					when "01111001000111001" => rgb <= "000000";
					when "01111001000111010" => rgb <= "000000";
					when "01111001000111011" => rgb <= "000000";
					when "01111001000111100" => rgb <= "000000";
					when "01111001000111101" => rgb <= "000000";
					when "01111001000111110" => rgb <= "000000";
					when "01111001000111111" => rgb <= "000000";
					when "01111001001000000" => rgb <= "000000";
					when "01111001001000001" => rgb <= "000000";
					when "01111001001000010" => rgb <= "000000";
					when "01111001001000011" => rgb <= "000000";
					when "01111001001000100" => rgb <= "000000";
					when "01111001001000101" => rgb <= "000000";
					when "01111001001000110" => rgb <= "000000";
					when "01111001001000111" => rgb <= "000000";
					when "01111001001001000" => rgb <= "000000";
					when "01111001001001001" => rgb <= "000000";
					when "01111001001001010" => rgb <= "000000";
					when "01111001001001011" => rgb <= "000000";
					when "01111001001001100" => rgb <= "000000";
					when "01111001001001101" => rgb <= "000000";
					when "01111001001001110" => rgb <= "000000";
					when "01111001001001111" => rgb <= "000000";
					when "01111001001010000" => rgb <= "000000";
					when "01111001001010001" => rgb <= "000000";
					when "01111001001010010" => rgb <= "000000";
					when "01111001001010011" => rgb <= "000000";
					when "01111001001010100" => rgb <= "000000";
					when "01111001001010101" => rgb <= "000000";
					when "01111001001010110" => rgb <= "000000";
					when "01111001001010111" => rgb <= "000000";
					when "01111001001011000" => rgb <= "000000";
					when "01111001001011001" => rgb <= "000000";
					when "01111001001011010" => rgb <= "000000";
					when "01111001001011011" => rgb <= "000000";
					when "01111001001011100" => rgb <= "000000";
					when "01111001001011101" => rgb <= "000000";
					when "01111001001011110" => rgb <= "000000";
					when "01111001001011111" => rgb <= "000000";
					when "01111001001100000" => rgb <= "000000";
					when "01111001001100001" => rgb <= "000000";
					when "01111001001100010" => rgb <= "000000";
					when "01111001001100011" => rgb <= "000000";
					when "01111001001100100" => rgb <= "000000";
					when "01111001001100101" => rgb <= "000000";
					when "01111001001100110" => rgb <= "000000";
					when "01111001001100111" => rgb <= "000000";
					when "01111001001101000" => rgb <= "000000";
					when "01111001001101001" => rgb <= "000000";
					when "01111001001101010" => rgb <= "000000";
					when "01111001001101011" => rgb <= "000000";
					when "01111001001101100" => rgb <= "000000";
					when "01111001001101101" => rgb <= "000000";
					when "01111001001101110" => rgb <= "000000";
					when "01111001001101111" => rgb <= "000000";
					when "01111001001110000" => rgb <= "000000";
					when "01111001001110001" => rgb <= "000000";
					when "01111001001110010" => rgb <= "000000";
					when "01111001001110011" => rgb <= "000000";
					when "01111001001110100" => rgb <= "000000";
					when "01111001001110101" => rgb <= "000000";
					when "01111001001110110" => rgb <= "000000";
					when "01111001001110111" => rgb <= "000000";
					when "01111001001111000" => rgb <= "000000";
					when "01111001001111001" => rgb <= "000000";
					when "01111001001111010" => rgb <= "000000";
					when "01111001001111011" => rgb <= "000000";
					when "01111001001111100" => rgb <= "000000";
					when "01111001001111101" => rgb <= "000000";
					when "01111001001111110" => rgb <= "000000";
					when "01111001001111111" => rgb <= "000000";
					when "01111001010000000" => rgb <= "000000";
					when "01111001010000001" => rgb <= "000000";
					when "01111001010000010" => rgb <= "000000";
					when "01111001010000011" => rgb <= "000000";
					when "01111001010000100" => rgb <= "000000";
					when "01111001010000101" => rgb <= "000000";
					when "01111001010000110" => rgb <= "000000";
					when "01111001010000111" => rgb <= "000000";
					when "01111001010001000" => rgb <= "000000";
					when "01111001010001001" => rgb <= "000000";
					when "01111001010001010" => rgb <= "000000";
					when "01111001010001011" => rgb <= "000000";
					when "01111001010001100" => rgb <= "000000";
					when "01111001010001101" => rgb <= "000000";
					when "01111001010001110" => rgb <= "000000";
					when "01111001010001111" => rgb <= "000000";
					when "01111001010010000" => rgb <= "000000";
					when "01111001010010001" => rgb <= "000000";
					when "01111001010010010" => rgb <= "000000";
					when "01111001010010011" => rgb <= "000000";
					when "01111001010010100" => rgb <= "000000";
					when "01111001010010101" => rgb <= "000000";
					when "01111001010010110" => rgb <= "000000";
					when "01111001010010111" => rgb <= "000000";
					when "01111001010011000" => rgb <= "000000";
					when "01111001010011001" => rgb <= "000000";
					when "01111001010011010" => rgb <= "000000";
					when "01111001010011011" => rgb <= "000000";
					when "01111001010011100" => rgb <= "000000";
					when "01111001010011101" => rgb <= "000000";
					when "01111001010011110" => rgb <= "000000";
					when "01111001010011111" => rgb <= "000000";
					when "01111001010100000" => rgb <= "000000";
					when "01111001010100001" => rgb <= "000000";
					when "01111001010100010" => rgb <= "000000";
					when "01111001010100011" => rgb <= "000000";
					when "01111001010100100" => rgb <= "000000";
					when "01111001010100101" => rgb <= "000000";
					when "01111001010100110" => rgb <= "000000";
					when "01111001010100111" => rgb <= "000000";
					when "01111001010101000" => rgb <= "000000";
					when "01111001010101001" => rgb <= "000000";
					when "01111001010101010" => rgb <= "000000";
					when "01111001010101011" => rgb <= "000000";
					when "01111001010101100" => rgb <= "000000";
					when "01111001010101101" => rgb <= "000000";
					when "01111001010101110" => rgb <= "000000";
					when "01111001010101111" => rgb <= "000000";
					when "01111001010110000" => rgb <= "000000";
					when "01111001010110001" => rgb <= "000000";
					when "01111001010110010" => rgb <= "000000";
					when "01111001010110011" => rgb <= "000000";
					when "01111001010110100" => rgb <= "000000";
					when "01111001010110101" => rgb <= "000000";
					when "01111001010110110" => rgb <= "000000";
					when "01111001010110111" => rgb <= "000000";
					when "01111001010111000" => rgb <= "000000";
					when "01111001010111001" => rgb <= "000000";
					when "01111001010111010" => rgb <= "000000";
					when "01111001010111011" => rgb <= "000000";
					when "01111001010111100" => rgb <= "000000";
					when "01111001010111101" => rgb <= "000000";
					when "01111001010111110" => rgb <= "000000";
					when "01111001010111111" => rgb <= "000000";
					when "01111001011000000" => rgb <= "000000";
					when "01111001011000001" => rgb <= "000000";
					when "01111001011000010" => rgb <= "000000";
					when "01111001011000011" => rgb <= "000000";
					when "01111001011000100" => rgb <= "000000";
					when "01111001011000101" => rgb <= "000000";
					when "01111001011000110" => rgb <= "000000";
					when "01111001011000111" => rgb <= "000000";
					when "01111001011001000" => rgb <= "000000";
					when "01111001011001001" => rgb <= "000000";
					when "01111001011001010" => rgb <= "000000";
					when "01111001011001011" => rgb <= "000000";
					when "01111001011001100" => rgb <= "000000";
					when "01111001011001101" => rgb <= "000000";
					when "01111001011001110" => rgb <= "000000";
					when "01111001011001111" => rgb <= "000000";
					when "01111001011010000" => rgb <= "000000";
					when "01111001011010001" => rgb <= "000000";
					when "01111001011010010" => rgb <= "000000";
					when "01111001011010011" => rgb <= "000000";
					when "01111001011010100" => rgb <= "000000";
					when "01111001011010101" => rgb <= "000000";
					when "01111001011010110" => rgb <= "000000";
					when "01111001011010111" => rgb <= "000000";
					when "01111001011011000" => rgb <= "000000";
					when "01111001011011001" => rgb <= "000000";
					when "01111001011011010" => rgb <= "000000";
					when "01111001011011011" => rgb <= "000000";
					when "01111001011011100" => rgb <= "000000";
					when "01111001011011101" => rgb <= "000000";
					when "01111001011011110" => rgb <= "000000";
					when "01111001011011111" => rgb <= "000000";
					when "01111001011100000" => rgb <= "000000";
					when "01111001011100001" => rgb <= "000000";
					when "01111001011100010" => rgb <= "000000";
					when "01111001011100011" => rgb <= "000000";
					when "01111001011100100" => rgb <= "000000";
					when "01111001011100101" => rgb <= "000000";
					when "01111001011100110" => rgb <= "000000";
					when "01111001011100111" => rgb <= "000000";
					when "01111001011101000" => rgb <= "000000";
					when "01111001011101001" => rgb <= "000000";
					when "01111001011101010" => rgb <= "000000";
					when "01111001011101011" => rgb <= "000000";
					when "01111001011101100" => rgb <= "000000";
					when "01111001011101101" => rgb <= "000000";
					when "01111001011101110" => rgb <= "000000";
					when "01111001011101111" => rgb <= "000000";
					when "01111001011110000" => rgb <= "000000";
					when "01111001011110001" => rgb <= "000000";
					when "01111001011110010" => rgb <= "000000";
					when "01111001011110011" => rgb <= "000000";
					when "01111001011110100" => rgb <= "000000";
					when "01111001011110101" => rgb <= "000000";
					when "01111001011110110" => rgb <= "000000";
					when "01111001011110111" => rgb <= "000000";
					when "01111001011111000" => rgb <= "000000";
					when "01111001011111001" => rgb <= "000000";
					when "01111001011111010" => rgb <= "000000";
					when "01111001011111011" => rgb <= "000000";
					when "01111001011111100" => rgb <= "000000";
					when "01111001011111101" => rgb <= "000000";
					when "01111001011111110" => rgb <= "000000";
					when "01111001011111111" => rgb <= "000000";
					when "01111001100000000" => rgb <= "000000";
					when "01111001100000001" => rgb <= "000000";
					when "01111001100000010" => rgb <= "000000";
					when "01111001100000011" => rgb <= "000000";
					when "01111001100000100" => rgb <= "000000";
					when "01111001100000101" => rgb <= "000000";
					when "01111001100000110" => rgb <= "000000";
					when "01111001100000111" => rgb <= "000000";
					when "01111001100001000" => rgb <= "000000";
					when "01111001100001001" => rgb <= "000000";
					when "01111001100001010" => rgb <= "000000";
					when "01111001100001011" => rgb <= "000000";
					when "01111001100001100" => rgb <= "000000";
					when "01111001100001101" => rgb <= "000000";
					when "01111001100001110" => rgb <= "000000";
					when "01111001100001111" => rgb <= "000000";
					when "01111001100010000" => rgb <= "000000";
					when "01111001100010001" => rgb <= "000000";
					when "01111001100010010" => rgb <= "000000";
					when "01111001100010011" => rgb <= "000000";
					when "01111001100010100" => rgb <= "000000";
					when "01111001100010101" => rgb <= "000000";
					when "01111001100010110" => rgb <= "000000";
					when "01111001100010111" => rgb <= "000000";
					when "01111001100011000" => rgb <= "000000";
					when "01111001100011001" => rgb <= "000000";
					when "01111001100011010" => rgb <= "000000";
					when "01111001100011011" => rgb <= "000000";
					when "01111001100011100" => rgb <= "000000";
					when "01111001100011101" => rgb <= "000000";
					when "01111001100011110" => rgb <= "000000";
					when "01111001100011111" => rgb <= "000000";
					when "01111001100100000" => rgb <= "000000";
					when "01111001100100001" => rgb <= "000000";
					when "01111001100100010" => rgb <= "000000";
					when "01111001100100011" => rgb <= "000000";
					when "01111001100100100" => rgb <= "000000";
					when "01111001100100101" => rgb <= "000000";
					when "01111001100100110" => rgb <= "000000";
					when "01111001100100111" => rgb <= "000000";
					when "01111001100101000" => rgb <= "000000";
					when "01111001100101001" => rgb <= "000000";
					when "01111001100101010" => rgb <= "000000";
					when "01111001100101011" => rgb <= "000000";
					when "01111001100101100" => rgb <= "000000";
					when "01111001100101101" => rgb <= "000000";
					when "01111001100101110" => rgb <= "000000";
					when "01111001100101111" => rgb <= "000000";
					when "01111001100110000" => rgb <= "000000";
					when "01111001100110001" => rgb <= "000000";
					when "01111001100110010" => rgb <= "000000";
					when "01111001100110011" => rgb <= "000000";
					when "01111001100110100" => rgb <= "000000";
					when "01111001100110101" => rgb <= "000000";
					when "01111001100110110" => rgb <= "000000";
					when "01111001100110111" => rgb <= "000000";
					when "01111001100111000" => rgb <= "000000";
					when "01111001100111001" => rgb <= "000000";
					when "01111001100111010" => rgb <= "000000";
					when "01111001100111011" => rgb <= "000000";
					when "01111001100111100" => rgb <= "000000";
					when "01111001100111101" => rgb <= "000000";
					when "01111001100111110" => rgb <= "000000";
					when "01111001100111111" => rgb <= "000000";
					when "01111010000000000" => rgb <= "000000";
					when "01111010000000001" => rgb <= "000000";
					when "01111010000000010" => rgb <= "000000";
					when "01111010000000011" => rgb <= "000000";
					when "01111010000000100" => rgb <= "000000";
					when "01111010000000101" => rgb <= "000000";
					when "01111010000000110" => rgb <= "000000";
					when "01111010000000111" => rgb <= "000000";
					when "01111010000001000" => rgb <= "000000";
					when "01111010000001001" => rgb <= "000000";
					when "01111010000001010" => rgb <= "000000";
					when "01111010000001011" => rgb <= "000000";
					when "01111010000001100" => rgb <= "000000";
					when "01111010000001101" => rgb <= "000000";
					when "01111010000001110" => rgb <= "000000";
					when "01111010000001111" => rgb <= "000000";
					when "01111010000010000" => rgb <= "000000";
					when "01111010000010001" => rgb <= "000000";
					when "01111010000010010" => rgb <= "000000";
					when "01111010000010011" => rgb <= "000000";
					when "01111010000010100" => rgb <= "000000";
					when "01111010000010101" => rgb <= "000000";
					when "01111010000010110" => rgb <= "000000";
					when "01111010000010111" => rgb <= "000000";
					when "01111010000011000" => rgb <= "000000";
					when "01111010000011001" => rgb <= "000000";
					when "01111010000011010" => rgb <= "000000";
					when "01111010000011011" => rgb <= "000000";
					when "01111010000011100" => rgb <= "000000";
					when "01111010000011101" => rgb <= "000000";
					when "01111010000011110" => rgb <= "000000";
					when "01111010000011111" => rgb <= "000000";
					when "01111010000100000" => rgb <= "000000";
					when "01111010000100001" => rgb <= "000000";
					when "01111010000100010" => rgb <= "000000";
					when "01111010000100011" => rgb <= "000000";
					when "01111010000100100" => rgb <= "000000";
					when "01111010000100101" => rgb <= "000000";
					when "01111010000100110" => rgb <= "000000";
					when "01111010000100111" => rgb <= "000000";
					when "01111010000101000" => rgb <= "000000";
					when "01111010000101001" => rgb <= "000000";
					when "01111010000101010" => rgb <= "000000";
					when "01111010000101011" => rgb <= "000000";
					when "01111010000101100" => rgb <= "000000";
					when "01111010000101101" => rgb <= "000000";
					when "01111010000101110" => rgb <= "000000";
					when "01111010000101111" => rgb <= "000000";
					when "01111010000110000" => rgb <= "000000";
					when "01111010000110001" => rgb <= "000000";
					when "01111010000110010" => rgb <= "000000";
					when "01111010000110011" => rgb <= "000000";
					when "01111010000110100" => rgb <= "000000";
					when "01111010000110101" => rgb <= "000000";
					when "01111010000110110" => rgb <= "000000";
					when "01111010000110111" => rgb <= "000000";
					when "01111010000111000" => rgb <= "000000";
					when "01111010000111001" => rgb <= "000000";
					when "01111010000111010" => rgb <= "000000";
					when "01111010000111011" => rgb <= "000000";
					when "01111010000111100" => rgb <= "000000";
					when "01111010000111101" => rgb <= "000000";
					when "01111010000111110" => rgb <= "000000";
					when "01111010000111111" => rgb <= "000000";
					when "01111010001000000" => rgb <= "000000";
					when "01111010001000001" => rgb <= "000000";
					when "01111010001000010" => rgb <= "000000";
					when "01111010001000011" => rgb <= "000000";
					when "01111010001000100" => rgb <= "000000";
					when "01111010001000101" => rgb <= "000000";
					when "01111010001000110" => rgb <= "000000";
					when "01111010001000111" => rgb <= "000000";
					when "01111010001001000" => rgb <= "000000";
					when "01111010001001001" => rgb <= "000000";
					when "01111010001001010" => rgb <= "000000";
					when "01111010001001011" => rgb <= "000000";
					when "01111010001001100" => rgb <= "000000";
					when "01111010001001101" => rgb <= "000000";
					when "01111010001001110" => rgb <= "000000";
					when "01111010001001111" => rgb <= "000000";
					when "01111010001010000" => rgb <= "000000";
					when "01111010001010001" => rgb <= "000000";
					when "01111010001010010" => rgb <= "000000";
					when "01111010001010011" => rgb <= "000000";
					when "01111010001010100" => rgb <= "000000";
					when "01111010001010101" => rgb <= "000000";
					when "01111010001010110" => rgb <= "000000";
					when "01111010001010111" => rgb <= "000000";
					when "01111010001011000" => rgb <= "000000";
					when "01111010001011001" => rgb <= "000000";
					when "01111010001011010" => rgb <= "000000";
					when "01111010001011011" => rgb <= "000000";
					when "01111010001011100" => rgb <= "000000";
					when "01111010001011101" => rgb <= "000000";
					when "01111010001011110" => rgb <= "000000";
					when "01111010001011111" => rgb <= "000000";
					when "01111010001100000" => rgb <= "000000";
					when "01111010001100001" => rgb <= "000000";
					when "01111010001100010" => rgb <= "000000";
					when "01111010001100011" => rgb <= "000000";
					when "01111010001100100" => rgb <= "000000";
					when "01111010001100101" => rgb <= "000000";
					when "01111010001100110" => rgb <= "000000";
					when "01111010001100111" => rgb <= "000000";
					when "01111010001101000" => rgb <= "000000";
					when "01111010001101001" => rgb <= "000000";
					when "01111010001101010" => rgb <= "000000";
					when "01111010001101011" => rgb <= "000000";
					when "01111010001101100" => rgb <= "000000";
					when "01111010001101101" => rgb <= "000000";
					when "01111010001101110" => rgb <= "000000";
					when "01111010001101111" => rgb <= "000000";
					when "01111010001110000" => rgb <= "000000";
					when "01111010001110001" => rgb <= "000000";
					when "01111010001110010" => rgb <= "000000";
					when "01111010001110011" => rgb <= "000000";
					when "01111010001110100" => rgb <= "000000";
					when "01111010001110101" => rgb <= "000000";
					when "01111010001110110" => rgb <= "000000";
					when "01111010001110111" => rgb <= "000000";
					when "01111010001111000" => rgb <= "000000";
					when "01111010001111001" => rgb <= "000000";
					when "01111010001111010" => rgb <= "000000";
					when "01111010001111011" => rgb <= "000000";
					when "01111010001111100" => rgb <= "000000";
					when "01111010001111101" => rgb <= "000000";
					when "01111010001111110" => rgb <= "000000";
					when "01111010001111111" => rgb <= "000000";
					when "01111010010000000" => rgb <= "000000";
					when "01111010010000001" => rgb <= "000000";
					when "01111010010000010" => rgb <= "000000";
					when "01111010010000011" => rgb <= "000000";
					when "01111010010000100" => rgb <= "000000";
					when "01111010010000101" => rgb <= "000000";
					when "01111010010000110" => rgb <= "000000";
					when "01111010010000111" => rgb <= "000000";
					when "01111010010001000" => rgb <= "000000";
					when "01111010010001001" => rgb <= "000000";
					when "01111010010001010" => rgb <= "000000";
					when "01111010010001011" => rgb <= "000000";
					when "01111010010001100" => rgb <= "000000";
					when "01111010010001101" => rgb <= "000000";
					when "01111010010001110" => rgb <= "000000";
					when "01111010010001111" => rgb <= "000000";
					when "01111010010010000" => rgb <= "000000";
					when "01111010010010001" => rgb <= "000000";
					when "01111010010010010" => rgb <= "000000";
					when "01111010010010011" => rgb <= "000000";
					when "01111010010010100" => rgb <= "000000";
					when "01111010010010101" => rgb <= "000000";
					when "01111010010010110" => rgb <= "000000";
					when "01111010010010111" => rgb <= "000000";
					when "01111010010011000" => rgb <= "000000";
					when "01111010010011001" => rgb <= "000000";
					when "01111010010011010" => rgb <= "000000";
					when "01111010010011011" => rgb <= "000000";
					when "01111010010011100" => rgb <= "000000";
					when "01111010010011101" => rgb <= "000000";
					when "01111010010011110" => rgb <= "000000";
					when "01111010010011111" => rgb <= "000000";
					when "01111010010100000" => rgb <= "000000";
					when "01111010010100001" => rgb <= "000000";
					when "01111010010100010" => rgb <= "000000";
					when "01111010010100011" => rgb <= "000000";
					when "01111010010100100" => rgb <= "000000";
					when "01111010010100101" => rgb <= "000000";
					when "01111010010100110" => rgb <= "000000";
					when "01111010010100111" => rgb <= "000000";
					when "01111010010101000" => rgb <= "000000";
					when "01111010010101001" => rgb <= "000000";
					when "01111010010101010" => rgb <= "000000";
					when "01111010010101011" => rgb <= "000000";
					when "01111010010101100" => rgb <= "000000";
					when "01111010010101101" => rgb <= "000000";
					when "01111010010101110" => rgb <= "000000";
					when "01111010010101111" => rgb <= "000000";
					when "01111010010110000" => rgb <= "000000";
					when "01111010010110001" => rgb <= "000000";
					when "01111010010110010" => rgb <= "000000";
					when "01111010010110011" => rgb <= "000000";
					when "01111010010110100" => rgb <= "000000";
					when "01111010010110101" => rgb <= "000000";
					when "01111010010110110" => rgb <= "000000";
					when "01111010010110111" => rgb <= "000000";
					when "01111010010111000" => rgb <= "000000";
					when "01111010010111001" => rgb <= "000000";
					when "01111010010111010" => rgb <= "000000";
					when "01111010010111011" => rgb <= "000000";
					when "01111010010111100" => rgb <= "000000";
					when "01111010010111101" => rgb <= "000000";
					when "01111010010111110" => rgb <= "000000";
					when "01111010010111111" => rgb <= "000000";
					when "01111010011000000" => rgb <= "000000";
					when "01111010011000001" => rgb <= "000000";
					when "01111010011000010" => rgb <= "000000";
					when "01111010011000011" => rgb <= "000000";
					when "01111010011000100" => rgb <= "000000";
					when "01111010011000101" => rgb <= "000000";
					when "01111010011000110" => rgb <= "000000";
					when "01111010011000111" => rgb <= "000000";
					when "01111010011001000" => rgb <= "000000";
					when "01111010011001001" => rgb <= "000000";
					when "01111010011001010" => rgb <= "000000";
					when "01111010011001011" => rgb <= "000000";
					when "01111010011001100" => rgb <= "000000";
					when "01111010011001101" => rgb <= "000000";
					when "01111010011001110" => rgb <= "000000";
					when "01111010011001111" => rgb <= "000000";
					when "01111010011010000" => rgb <= "000000";
					when "01111010011010001" => rgb <= "000000";
					when "01111010011010010" => rgb <= "000000";
					when "01111010011010011" => rgb <= "000000";
					when "01111010011010100" => rgb <= "000000";
					when "01111010011010101" => rgb <= "000000";
					when "01111010011010110" => rgb <= "000000";
					when "01111010011010111" => rgb <= "000000";
					when "01111010011011000" => rgb <= "000000";
					when "01111010011011001" => rgb <= "000000";
					when "01111010011011010" => rgb <= "000000";
					when "01111010011011011" => rgb <= "000000";
					when "01111010011011100" => rgb <= "000000";
					when "01111010011011101" => rgb <= "000000";
					when "01111010011011110" => rgb <= "000000";
					when "01111010011011111" => rgb <= "000000";
					when "01111010011100000" => rgb <= "000000";
					when "01111010011100001" => rgb <= "000000";
					when "01111010011100010" => rgb <= "000000";
					when "01111010011100011" => rgb <= "000000";
					when "01111010011100100" => rgb <= "000000";
					when "01111010011100101" => rgb <= "000000";
					when "01111010011100110" => rgb <= "000000";
					when "01111010011100111" => rgb <= "000000";
					when "01111010011101000" => rgb <= "000000";
					when "01111010011101001" => rgb <= "000000";
					when "01111010011101010" => rgb <= "000000";
					when "01111010011101011" => rgb <= "000000";
					when "01111010011101100" => rgb <= "000000";
					when "01111010011101101" => rgb <= "000000";
					when "01111010011101110" => rgb <= "000000";
					when "01111010011101111" => rgb <= "000000";
					when "01111010011110000" => rgb <= "000000";
					when "01111010011110001" => rgb <= "000000";
					when "01111010011110010" => rgb <= "000000";
					when "01111010011110011" => rgb <= "000000";
					when "01111010011110100" => rgb <= "000000";
					when "01111010011110101" => rgb <= "000000";
					when "01111010011110110" => rgb <= "000000";
					when "01111010011110111" => rgb <= "000000";
					when "01111010011111000" => rgb <= "000000";
					when "01111010011111001" => rgb <= "000000";
					when "01111010011111010" => rgb <= "000000";
					when "01111010011111011" => rgb <= "000000";
					when "01111010011111100" => rgb <= "000000";
					when "01111010011111101" => rgb <= "000000";
					when "01111010011111110" => rgb <= "000000";
					when "01111010011111111" => rgb <= "000000";
					when "01111010100000000" => rgb <= "000000";
					when "01111010100000001" => rgb <= "000000";
					when "01111010100000010" => rgb <= "000000";
					when "01111010100000011" => rgb <= "000000";
					when "01111010100000100" => rgb <= "000000";
					when "01111010100000101" => rgb <= "000000";
					when "01111010100000110" => rgb <= "000000";
					when "01111010100000111" => rgb <= "000000";
					when "01111010100001000" => rgb <= "000000";
					when "01111010100001001" => rgb <= "000000";
					when "01111010100001010" => rgb <= "000000";
					when "01111010100001011" => rgb <= "000000";
					when "01111010100001100" => rgb <= "000000";
					when "01111010100001101" => rgb <= "000000";
					when "01111010100001110" => rgb <= "000000";
					when "01111010100001111" => rgb <= "000000";
					when "01111010100010000" => rgb <= "000000";
					when "01111010100010001" => rgb <= "000000";
					when "01111010100010010" => rgb <= "000000";
					when "01111010100010011" => rgb <= "000000";
					when "01111010100010100" => rgb <= "000000";
					when "01111010100010101" => rgb <= "000000";
					when "01111010100010110" => rgb <= "000000";
					when "01111010100010111" => rgb <= "000000";
					when "01111010100011000" => rgb <= "000000";
					when "01111010100011001" => rgb <= "000000";
					when "01111010100011010" => rgb <= "000000";
					when "01111010100011011" => rgb <= "000000";
					when "01111010100011100" => rgb <= "000000";
					when "01111010100011101" => rgb <= "000000";
					when "01111010100011110" => rgb <= "000000";
					when "01111010100011111" => rgb <= "000000";
					when "01111010100100000" => rgb <= "000000";
					when "01111010100100001" => rgb <= "000000";
					when "01111010100100010" => rgb <= "000000";
					when "01111010100100011" => rgb <= "000000";
					when "01111010100100100" => rgb <= "000000";
					when "01111010100100101" => rgb <= "000000";
					when "01111010100100110" => rgb <= "000000";
					when "01111010100100111" => rgb <= "000000";
					when "01111010100101000" => rgb <= "000000";
					when "01111010100101001" => rgb <= "000000";
					when "01111010100101010" => rgb <= "000000";
					when "01111010100101011" => rgb <= "000000";
					when "01111010100101100" => rgb <= "000000";
					when "01111010100101101" => rgb <= "000000";
					when "01111010100101110" => rgb <= "000000";
					when "01111010100101111" => rgb <= "000000";
					when "01111010100110000" => rgb <= "000000";
					when "01111010100110001" => rgb <= "000000";
					when "01111010100110010" => rgb <= "000000";
					when "01111010100110011" => rgb <= "000000";
					when "01111010100110100" => rgb <= "000000";
					when "01111010100110101" => rgb <= "000000";
					when "01111010100110110" => rgb <= "000000";
					when "01111010100110111" => rgb <= "000000";
					when "01111010100111000" => rgb <= "000000";
					when "01111010100111001" => rgb <= "000000";
					when "01111010100111010" => rgb <= "000000";
					when "01111010100111011" => rgb <= "000000";
					when "01111010100111100" => rgb <= "000000";
					when "01111010100111101" => rgb <= "000000";
					when "01111010100111110" => rgb <= "000000";
					when "01111010100111111" => rgb <= "000000";
					when "01111011000000000" => rgb <= "000000";
					when "01111011000000001" => rgb <= "000000";
					when "01111011000000010" => rgb <= "000000";
					when "01111011000000011" => rgb <= "000000";
					when "01111011000000100" => rgb <= "000000";
					when "01111011000000101" => rgb <= "000000";
					when "01111011000000110" => rgb <= "000000";
					when "01111011000000111" => rgb <= "000000";
					when "01111011000001000" => rgb <= "000000";
					when "01111011000001001" => rgb <= "000000";
					when "01111011000001010" => rgb <= "000000";
					when "01111011000001011" => rgb <= "000000";
					when "01111011000001100" => rgb <= "000000";
					when "01111011000001101" => rgb <= "000000";
					when "01111011000001110" => rgb <= "000000";
					when "01111011000001111" => rgb <= "000000";
					when "01111011000010000" => rgb <= "000000";
					when "01111011000010001" => rgb <= "000000";
					when "01111011000010010" => rgb <= "000000";
					when "01111011000010011" => rgb <= "000000";
					when "01111011000010100" => rgb <= "000000";
					when "01111011000010101" => rgb <= "000000";
					when "01111011000010110" => rgb <= "000000";
					when "01111011000010111" => rgb <= "000000";
					when "01111011000011000" => rgb <= "000000";
					when "01111011000011001" => rgb <= "000000";
					when "01111011000011010" => rgb <= "000000";
					when "01111011000011011" => rgb <= "000000";
					when "01111011000011100" => rgb <= "000000";
					when "01111011000011101" => rgb <= "000000";
					when "01111011000011110" => rgb <= "000000";
					when "01111011000011111" => rgb <= "000000";
					when "01111011000100000" => rgb <= "000000";
					when "01111011000100001" => rgb <= "000000";
					when "01111011000100010" => rgb <= "000000";
					when "01111011000100011" => rgb <= "000000";
					when "01111011000100100" => rgb <= "000000";
					when "01111011000100101" => rgb <= "000000";
					when "01111011000100110" => rgb <= "000000";
					when "01111011000100111" => rgb <= "000000";
					when "01111011000101000" => rgb <= "000000";
					when "01111011000101001" => rgb <= "000000";
					when "01111011000101010" => rgb <= "000000";
					when "01111011000101011" => rgb <= "000000";
					when "01111011000101100" => rgb <= "000000";
					when "01111011000101101" => rgb <= "000000";
					when "01111011000101110" => rgb <= "000000";
					when "01111011000101111" => rgb <= "000000";
					when "01111011000110000" => rgb <= "000000";
					when "01111011000110001" => rgb <= "000000";
					when "01111011000110010" => rgb <= "000000";
					when "01111011000110011" => rgb <= "000000";
					when "01111011000110100" => rgb <= "000000";
					when "01111011000110101" => rgb <= "000000";
					when "01111011000110110" => rgb <= "000000";
					when "01111011000110111" => rgb <= "000000";
					when "01111011000111000" => rgb <= "000000";
					when "01111011000111001" => rgb <= "000000";
					when "01111011000111010" => rgb <= "000000";
					when "01111011000111011" => rgb <= "000000";
					when "01111011000111100" => rgb <= "000000";
					when "01111011000111101" => rgb <= "000000";
					when "01111011000111110" => rgb <= "000000";
					when "01111011000111111" => rgb <= "000000";
					when "01111011001000000" => rgb <= "000000";
					when "01111011001000001" => rgb <= "000000";
					when "01111011001000010" => rgb <= "000000";
					when "01111011001000011" => rgb <= "000000";
					when "01111011001000100" => rgb <= "000000";
					when "01111011001000101" => rgb <= "000000";
					when "01111011001000110" => rgb <= "000000";
					when "01111011001000111" => rgb <= "000000";
					when "01111011001001000" => rgb <= "000000";
					when "01111011001001001" => rgb <= "000000";
					when "01111011001001010" => rgb <= "000000";
					when "01111011001001011" => rgb <= "000000";
					when "01111011001001100" => rgb <= "000000";
					when "01111011001001101" => rgb <= "000000";
					when "01111011001001110" => rgb <= "000000";
					when "01111011001001111" => rgb <= "000000";
					when "01111011001010000" => rgb <= "000000";
					when "01111011001010001" => rgb <= "000000";
					when "01111011001010010" => rgb <= "000000";
					when "01111011001010011" => rgb <= "000000";
					when "01111011001010100" => rgb <= "000000";
					when "01111011001010101" => rgb <= "000000";
					when "01111011001010110" => rgb <= "000000";
					when "01111011001010111" => rgb <= "000000";
					when "01111011001011000" => rgb <= "000000";
					when "01111011001011001" => rgb <= "000000";
					when "01111011001011010" => rgb <= "000000";
					when "01111011001011011" => rgb <= "000000";
					when "01111011001011100" => rgb <= "000000";
					when "01111011001011101" => rgb <= "000000";
					when "01111011001011110" => rgb <= "000000";
					when "01111011001011111" => rgb <= "000000";
					when "01111011001100000" => rgb <= "000000";
					when "01111011001100001" => rgb <= "000000";
					when "01111011001100010" => rgb <= "000000";
					when "01111011001100011" => rgb <= "000000";
					when "01111011001100100" => rgb <= "000000";
					when "01111011001100101" => rgb <= "000000";
					when "01111011001100110" => rgb <= "000000";
					when "01111011001100111" => rgb <= "000000";
					when "01111011001101000" => rgb <= "000000";
					when "01111011001101001" => rgb <= "000000";
					when "01111011001101010" => rgb <= "000000";
					when "01111011001101011" => rgb <= "000000";
					when "01111011001101100" => rgb <= "000000";
					when "01111011001101101" => rgb <= "000000";
					when "01111011001101110" => rgb <= "000000";
					when "01111011001101111" => rgb <= "000000";
					when "01111011001110000" => rgb <= "000000";
					when "01111011001110001" => rgb <= "000000";
					when "01111011001110010" => rgb <= "000000";
					when "01111011001110011" => rgb <= "000000";
					when "01111011001110100" => rgb <= "000000";
					when "01111011001110101" => rgb <= "000000";
					when "01111011001110110" => rgb <= "000000";
					when "01111011001110111" => rgb <= "000000";
					when "01111011001111000" => rgb <= "000000";
					when "01111011001111001" => rgb <= "000000";
					when "01111011001111010" => rgb <= "000000";
					when "01111011001111011" => rgb <= "000000";
					when "01111011001111100" => rgb <= "000000";
					when "01111011001111101" => rgb <= "000000";
					when "01111011001111110" => rgb <= "000000";
					when "01111011001111111" => rgb <= "000000";
					when "01111011010000000" => rgb <= "000000";
					when "01111011010000001" => rgb <= "000000";
					when "01111011010000010" => rgb <= "000000";
					when "01111011010000011" => rgb <= "000000";
					when "01111011010000100" => rgb <= "000000";
					when "01111011010000101" => rgb <= "000000";
					when "01111011010000110" => rgb <= "000000";
					when "01111011010000111" => rgb <= "000000";
					when "01111011010001000" => rgb <= "000000";
					when "01111011010001001" => rgb <= "000000";
					when "01111011010001010" => rgb <= "000000";
					when "01111011010001011" => rgb <= "000000";
					when "01111011010001100" => rgb <= "000000";
					when "01111011010001101" => rgb <= "000000";
					when "01111011010001110" => rgb <= "000000";
					when "01111011010001111" => rgb <= "000000";
					when "01111011010010000" => rgb <= "000000";
					when "01111011010010001" => rgb <= "000000";
					when "01111011010010010" => rgb <= "000000";
					when "01111011010010011" => rgb <= "000000";
					when "01111011010010100" => rgb <= "000000";
					when "01111011010010101" => rgb <= "000000";
					when "01111011010010110" => rgb <= "000000";
					when "01111011010010111" => rgb <= "000000";
					when "01111011010011000" => rgb <= "000000";
					when "01111011010011001" => rgb <= "000000";
					when "01111011010011010" => rgb <= "000000";
					when "01111011010011011" => rgb <= "000000";
					when "01111011010011100" => rgb <= "000000";
					when "01111011010011101" => rgb <= "000000";
					when "01111011010011110" => rgb <= "000000";
					when "01111011010011111" => rgb <= "000000";
					when "01111011010100000" => rgb <= "000000";
					when "01111011010100001" => rgb <= "000000";
					when "01111011010100010" => rgb <= "000000";
					when "01111011010100011" => rgb <= "000000";
					when "01111011010100100" => rgb <= "000000";
					when "01111011010100101" => rgb <= "000000";
					when "01111011010100110" => rgb <= "000000";
					when "01111011010100111" => rgb <= "000000";
					when "01111011010101000" => rgb <= "000000";
					when "01111011010101001" => rgb <= "000000";
					when "01111011010101010" => rgb <= "000000";
					when "01111011010101011" => rgb <= "000000";
					when "01111011010101100" => rgb <= "000000";
					when "01111011010101101" => rgb <= "000000";
					when "01111011010101110" => rgb <= "000000";
					when "01111011010101111" => rgb <= "000000";
					when "01111011010110000" => rgb <= "000000";
					when "01111011010110001" => rgb <= "000000";
					when "01111011010110010" => rgb <= "000000";
					when "01111011010110011" => rgb <= "000000";
					when "01111011010110100" => rgb <= "000000";
					when "01111011010110101" => rgb <= "000000";
					when "01111011010110110" => rgb <= "000000";
					when "01111011010110111" => rgb <= "000000";
					when "01111011010111000" => rgb <= "000000";
					when "01111011010111001" => rgb <= "000000";
					when "01111011010111010" => rgb <= "000000";
					when "01111011010111011" => rgb <= "000000";
					when "01111011010111100" => rgb <= "000000";
					when "01111011010111101" => rgb <= "000000";
					when "01111011010111110" => rgb <= "000000";
					when "01111011010111111" => rgb <= "000000";
					when "01111011011000000" => rgb <= "000000";
					when "01111011011000001" => rgb <= "000000";
					when "01111011011000010" => rgb <= "000000";
					when "01111011011000011" => rgb <= "000000";
					when "01111011011000100" => rgb <= "000000";
					when "01111011011000101" => rgb <= "000000";
					when "01111011011000110" => rgb <= "000000";
					when "01111011011000111" => rgb <= "000000";
					when "01111011011001000" => rgb <= "000000";
					when "01111011011001001" => rgb <= "000000";
					when "01111011011001010" => rgb <= "000000";
					when "01111011011001011" => rgb <= "000000";
					when "01111011011001100" => rgb <= "000000";
					when "01111011011001101" => rgb <= "000000";
					when "01111011011001110" => rgb <= "000000";
					when "01111011011001111" => rgb <= "000000";
					when "01111011011010000" => rgb <= "000000";
					when "01111011011010001" => rgb <= "000000";
					when "01111011011010010" => rgb <= "000000";
					when "01111011011010011" => rgb <= "000000";
					when "01111011011010100" => rgb <= "000000";
					when "01111011011010101" => rgb <= "000000";
					when "01111011011010110" => rgb <= "000000";
					when "01111011011010111" => rgb <= "000000";
					when "01111011011011000" => rgb <= "000000";
					when "01111011011011001" => rgb <= "000000";
					when "01111011011011010" => rgb <= "000000";
					when "01111011011011011" => rgb <= "000000";
					when "01111011011011100" => rgb <= "000000";
					when "01111011011011101" => rgb <= "000000";
					when "01111011011011110" => rgb <= "000000";
					when "01111011011011111" => rgb <= "000000";
					when "01111011011100000" => rgb <= "000000";
					when "01111011011100001" => rgb <= "000000";
					when "01111011011100010" => rgb <= "000000";
					when "01111011011100011" => rgb <= "000000";
					when "01111011011100100" => rgb <= "000000";
					when "01111011011100101" => rgb <= "000000";
					when "01111011011100110" => rgb <= "000000";
					when "01111011011100111" => rgb <= "000000";
					when "01111011011101000" => rgb <= "000000";
					when "01111011011101001" => rgb <= "000000";
					when "01111011011101010" => rgb <= "000000";
					when "01111011011101011" => rgb <= "000000";
					when "01111011011101100" => rgb <= "000000";
					when "01111011011101101" => rgb <= "000000";
					when "01111011011101110" => rgb <= "000000";
					when "01111011011101111" => rgb <= "000000";
					when "01111011011110000" => rgb <= "000000";
					when "01111011011110001" => rgb <= "000000";
					when "01111011011110010" => rgb <= "000000";
					when "01111011011110011" => rgb <= "000000";
					when "01111011011110100" => rgb <= "000000";
					when "01111011011110101" => rgb <= "000000";
					when "01111011011110110" => rgb <= "000000";
					when "01111011011110111" => rgb <= "000000";
					when "01111011011111000" => rgb <= "000000";
					when "01111011011111001" => rgb <= "000000";
					when "01111011011111010" => rgb <= "000000";
					when "01111011011111011" => rgb <= "000000";
					when "01111011011111100" => rgb <= "000000";
					when "01111011011111101" => rgb <= "000000";
					when "01111011011111110" => rgb <= "000000";
					when "01111011011111111" => rgb <= "000000";
					when "01111011100000000" => rgb <= "000000";
					when "01111011100000001" => rgb <= "000000";
					when "01111011100000010" => rgb <= "000000";
					when "01111011100000011" => rgb <= "000000";
					when "01111011100000100" => rgb <= "000000";
					when "01111011100000101" => rgb <= "000000";
					when "01111011100000110" => rgb <= "000000";
					when "01111011100000111" => rgb <= "000000";
					when "01111011100001000" => rgb <= "000000";
					when "01111011100001001" => rgb <= "000000";
					when "01111011100001010" => rgb <= "000000";
					when "01111011100001011" => rgb <= "000000";
					when "01111011100001100" => rgb <= "000000";
					when "01111011100001101" => rgb <= "000000";
					when "01111011100001110" => rgb <= "000000";
					when "01111011100001111" => rgb <= "000000";
					when "01111011100010000" => rgb <= "000000";
					when "01111011100010001" => rgb <= "000000";
					when "01111011100010010" => rgb <= "000000";
					when "01111011100010011" => rgb <= "000000";
					when "01111011100010100" => rgb <= "000000";
					when "01111011100010101" => rgb <= "000000";
					when "01111011100010110" => rgb <= "000000";
					when "01111011100010111" => rgb <= "000000";
					when "01111011100011000" => rgb <= "000000";
					when "01111011100011001" => rgb <= "000000";
					when "01111011100011010" => rgb <= "000000";
					when "01111011100011011" => rgb <= "000000";
					when "01111011100011100" => rgb <= "000000";
					when "01111011100011101" => rgb <= "000000";
					when "01111011100011110" => rgb <= "000000";
					when "01111011100011111" => rgb <= "000000";
					when "01111011100100000" => rgb <= "000000";
					when "01111011100100001" => rgb <= "000000";
					when "01111011100100010" => rgb <= "000000";
					when "01111011100100011" => rgb <= "000000";
					when "01111011100100100" => rgb <= "000000";
					when "01111011100100101" => rgb <= "000000";
					when "01111011100100110" => rgb <= "000000";
					when "01111011100100111" => rgb <= "000000";
					when "01111011100101000" => rgb <= "000000";
					when "01111011100101001" => rgb <= "000000";
					when "01111011100101010" => rgb <= "000000";
					when "01111011100101011" => rgb <= "000000";
					when "01111011100101100" => rgb <= "000000";
					when "01111011100101101" => rgb <= "000000";
					when "01111011100101110" => rgb <= "000000";
					when "01111011100101111" => rgb <= "000000";
					when "01111011100110000" => rgb <= "000000";
					when "01111011100110001" => rgb <= "000000";
					when "01111011100110010" => rgb <= "000000";
					when "01111011100110011" => rgb <= "000000";
					when "01111011100110100" => rgb <= "000000";
					when "01111011100110101" => rgb <= "000000";
					when "01111011100110110" => rgb <= "000000";
					when "01111011100110111" => rgb <= "000000";
					when "01111011100111000" => rgb <= "000000";
					when "01111011100111001" => rgb <= "000000";
					when "01111011100111010" => rgb <= "000000";
					when "01111011100111011" => rgb <= "000000";
					when "01111011100111100" => rgb <= "000000";
					when "01111011100111101" => rgb <= "000000";
					when "01111011100111110" => rgb <= "000000";
					when "01111011100111111" => rgb <= "000000";
					when "01111100000000000" => rgb <= "000000";
					when "01111100000000001" => rgb <= "000000";
					when "01111100000000010" => rgb <= "000000";
					when "01111100000000011" => rgb <= "000000";
					when "01111100000000100" => rgb <= "000000";
					when "01111100000000101" => rgb <= "000000";
					when "01111100000000110" => rgb <= "000000";
					when "01111100000000111" => rgb <= "000000";
					when "01111100000001000" => rgb <= "000000";
					when "01111100000001001" => rgb <= "000000";
					when "01111100000001010" => rgb <= "000000";
					when "01111100000001011" => rgb <= "000000";
					when "01111100000001100" => rgb <= "000000";
					when "01111100000001101" => rgb <= "000000";
					when "01111100000001110" => rgb <= "000000";
					when "01111100000001111" => rgb <= "000000";
					when "01111100000010000" => rgb <= "000000";
					when "01111100000010001" => rgb <= "000000";
					when "01111100000010010" => rgb <= "000000";
					when "01111100000010011" => rgb <= "000000";
					when "01111100000010100" => rgb <= "000000";
					when "01111100000010101" => rgb <= "000000";
					when "01111100000010110" => rgb <= "000000";
					when "01111100000010111" => rgb <= "000000";
					when "01111100000011000" => rgb <= "000000";
					when "01111100000011001" => rgb <= "000000";
					when "01111100000011010" => rgb <= "000000";
					when "01111100000011011" => rgb <= "000000";
					when "01111100000011100" => rgb <= "000000";
					when "01111100000011101" => rgb <= "000000";
					when "01111100000011110" => rgb <= "000000";
					when "01111100000011111" => rgb <= "000000";
					when "01111100000100000" => rgb <= "000000";
					when "01111100000100001" => rgb <= "000000";
					when "01111100000100010" => rgb <= "000000";
					when "01111100000100011" => rgb <= "000000";
					when "01111100000100100" => rgb <= "000000";
					when "01111100000100101" => rgb <= "000000";
					when "01111100000100110" => rgb <= "000000";
					when "01111100000100111" => rgb <= "000000";
					when "01111100000101000" => rgb <= "000000";
					when "01111100000101001" => rgb <= "000000";
					when "01111100000101010" => rgb <= "000000";
					when "01111100000101011" => rgb <= "000000";
					when "01111100000101100" => rgb <= "000000";
					when "01111100000101101" => rgb <= "000000";
					when "01111100000101110" => rgb <= "000000";
					when "01111100000101111" => rgb <= "000000";
					when "01111100000110000" => rgb <= "000000";
					when "01111100000110001" => rgb <= "000000";
					when "01111100000110010" => rgb <= "000000";
					when "01111100000110011" => rgb <= "000000";
					when "01111100000110100" => rgb <= "000000";
					when "01111100000110101" => rgb <= "000000";
					when "01111100000110110" => rgb <= "000000";
					when "01111100000110111" => rgb <= "000000";
					when "01111100000111000" => rgb <= "000000";
					when "01111100000111001" => rgb <= "000000";
					when "01111100000111010" => rgb <= "000000";
					when "01111100000111011" => rgb <= "000000";
					when "01111100000111100" => rgb <= "000000";
					when "01111100000111101" => rgb <= "000000";
					when "01111100000111110" => rgb <= "000000";
					when "01111100000111111" => rgb <= "000000";
					when "01111100001000000" => rgb <= "000000";
					when "01111100001000001" => rgb <= "000000";
					when "01111100001000010" => rgb <= "000000";
					when "01111100001000011" => rgb <= "000000";
					when "01111100001000100" => rgb <= "000000";
					when "01111100001000101" => rgb <= "000000";
					when "01111100001000110" => rgb <= "000000";
					when "01111100001000111" => rgb <= "000000";
					when "01111100001001000" => rgb <= "000000";
					when "01111100001001001" => rgb <= "000000";
					when "01111100001001010" => rgb <= "000000";
					when "01111100001001011" => rgb <= "000000";
					when "01111100001001100" => rgb <= "000000";
					when "01111100001001101" => rgb <= "000000";
					when "01111100001001110" => rgb <= "000000";
					when "01111100001001111" => rgb <= "000000";
					when "01111100001010000" => rgb <= "000000";
					when "01111100001010001" => rgb <= "000000";
					when "01111100001010010" => rgb <= "000000";
					when "01111100001010011" => rgb <= "000000";
					when "01111100001010100" => rgb <= "000000";
					when "01111100001010101" => rgb <= "000000";
					when "01111100001010110" => rgb <= "000000";
					when "01111100001010111" => rgb <= "000000";
					when "01111100001011000" => rgb <= "000000";
					when "01111100001011001" => rgb <= "000000";
					when "01111100001011010" => rgb <= "000000";
					when "01111100001011011" => rgb <= "000000";
					when "01111100001011100" => rgb <= "000000";
					when "01111100001011101" => rgb <= "000000";
					when "01111100001011110" => rgb <= "000000";
					when "01111100001011111" => rgb <= "000000";
					when "01111100001100000" => rgb <= "000000";
					when "01111100001100001" => rgb <= "000000";
					when "01111100001100010" => rgb <= "000000";
					when "01111100001100011" => rgb <= "000000";
					when "01111100001100100" => rgb <= "000000";
					when "01111100001100101" => rgb <= "000000";
					when "01111100001100110" => rgb <= "000000";
					when "01111100001100111" => rgb <= "000000";
					when "01111100001101000" => rgb <= "000000";
					when "01111100001101001" => rgb <= "000000";
					when "01111100001101010" => rgb <= "000000";
					when "01111100001101011" => rgb <= "000000";
					when "01111100001101100" => rgb <= "000000";
					when "01111100001101101" => rgb <= "000000";
					when "01111100001101110" => rgb <= "000000";
					when "01111100001101111" => rgb <= "000000";
					when "01111100001110000" => rgb <= "000000";
					when "01111100001110001" => rgb <= "000000";
					when "01111100001110010" => rgb <= "000000";
					when "01111100001110011" => rgb <= "000000";
					when "01111100001110100" => rgb <= "000000";
					when "01111100001110101" => rgb <= "000000";
					when "01111100001110110" => rgb <= "000000";
					when "01111100001110111" => rgb <= "000000";
					when "01111100001111000" => rgb <= "000000";
					when "01111100001111001" => rgb <= "000000";
					when "01111100001111010" => rgb <= "000000";
					when "01111100001111011" => rgb <= "000000";
					when "01111100001111100" => rgb <= "000000";
					when "01111100001111101" => rgb <= "000000";
					when "01111100001111110" => rgb <= "000000";
					when "01111100001111111" => rgb <= "000000";
					when "01111100010000000" => rgb <= "000000";
					when "01111100010000001" => rgb <= "000000";
					when "01111100010000010" => rgb <= "000000";
					when "01111100010000011" => rgb <= "000000";
					when "01111100010000100" => rgb <= "000000";
					when "01111100010000101" => rgb <= "000000";
					when "01111100010000110" => rgb <= "000000";
					when "01111100010000111" => rgb <= "000000";
					when "01111100010001000" => rgb <= "000000";
					when "01111100010001001" => rgb <= "000000";
					when "01111100010001010" => rgb <= "000000";
					when "01111100010001011" => rgb <= "000000";
					when "01111100010001100" => rgb <= "000000";
					when "01111100010001101" => rgb <= "000000";
					when "01111100010001110" => rgb <= "000000";
					when "01111100010001111" => rgb <= "000000";
					when "01111100010010000" => rgb <= "000000";
					when "01111100010010001" => rgb <= "000000";
					when "01111100010010010" => rgb <= "000000";
					when "01111100010010011" => rgb <= "000000";
					when "01111100010010100" => rgb <= "000000";
					when "01111100010010101" => rgb <= "000000";
					when "01111100010010110" => rgb <= "000000";
					when "01111100010010111" => rgb <= "000000";
					when "01111100010011000" => rgb <= "000000";
					when "01111100010011001" => rgb <= "000000";
					when "01111100010011010" => rgb <= "000000";
					when "01111100010011011" => rgb <= "000000";
					when "01111100010011100" => rgb <= "000000";
					when "01111100010011101" => rgb <= "000000";
					when "01111100010011110" => rgb <= "000000";
					when "01111100010011111" => rgb <= "000000";
					when "01111100010100000" => rgb <= "000000";
					when "01111100010100001" => rgb <= "000000";
					when "01111100010100010" => rgb <= "000000";
					when "01111100010100011" => rgb <= "000000";
					when "01111100010100100" => rgb <= "000000";
					when "01111100010100101" => rgb <= "000000";
					when "01111100010100110" => rgb <= "000000";
					when "01111100010100111" => rgb <= "000000";
					when "01111100010101000" => rgb <= "000000";
					when "01111100010101001" => rgb <= "000000";
					when "01111100010101010" => rgb <= "000000";
					when "01111100010101011" => rgb <= "000000";
					when "01111100010101100" => rgb <= "000000";
					when "01111100010101101" => rgb <= "000000";
					when "01111100010101110" => rgb <= "000000";
					when "01111100010101111" => rgb <= "000000";
					when "01111100010110000" => rgb <= "000000";
					when "01111100010110001" => rgb <= "000000";
					when "01111100010110010" => rgb <= "000000";
					when "01111100010110011" => rgb <= "000000";
					when "01111100010110100" => rgb <= "000000";
					when "01111100010110101" => rgb <= "000000";
					when "01111100010110110" => rgb <= "000000";
					when "01111100010110111" => rgb <= "000000";
					when "01111100010111000" => rgb <= "000000";
					when "01111100010111001" => rgb <= "000000";
					when "01111100010111010" => rgb <= "000000";
					when "01111100010111011" => rgb <= "000000";
					when "01111100010111100" => rgb <= "000000";
					when "01111100010111101" => rgb <= "000000";
					when "01111100010111110" => rgb <= "000000";
					when "01111100010111111" => rgb <= "000000";
					when "01111100011000000" => rgb <= "000000";
					when "01111100011000001" => rgb <= "000000";
					when "01111100011000010" => rgb <= "000000";
					when "01111100011000011" => rgb <= "000000";
					when "01111100011000100" => rgb <= "000000";
					when "01111100011000101" => rgb <= "000000";
					when "01111100011000110" => rgb <= "000000";
					when "01111100011000111" => rgb <= "000000";
					when "01111100011001000" => rgb <= "000000";
					when "01111100011001001" => rgb <= "000000";
					when "01111100011001010" => rgb <= "000000";
					when "01111100011001011" => rgb <= "000000";
					when "01111100011001100" => rgb <= "000000";
					when "01111100011001101" => rgb <= "000000";
					when "01111100011001110" => rgb <= "000000";
					when "01111100011001111" => rgb <= "000000";
					when "01111100011010000" => rgb <= "000000";
					when "01111100011010001" => rgb <= "000000";
					when "01111100011010010" => rgb <= "000000";
					when "01111100011010011" => rgb <= "000000";
					when "01111100011010100" => rgb <= "000000";
					when "01111100011010101" => rgb <= "000000";
					when "01111100011010110" => rgb <= "000000";
					when "01111100011010111" => rgb <= "000000";
					when "01111100011011000" => rgb <= "000000";
					when "01111100011011001" => rgb <= "000000";
					when "01111100011011010" => rgb <= "000000";
					when "01111100011011011" => rgb <= "000000";
					when "01111100011011100" => rgb <= "000000";
					when "01111100011011101" => rgb <= "000000";
					when "01111100011011110" => rgb <= "000000";
					when "01111100011011111" => rgb <= "000000";
					when "01111100011100000" => rgb <= "000000";
					when "01111100011100001" => rgb <= "000000";
					when "01111100011100010" => rgb <= "000000";
					when "01111100011100011" => rgb <= "000000";
					when "01111100011100100" => rgb <= "000000";
					when "01111100011100101" => rgb <= "000000";
					when "01111100011100110" => rgb <= "000000";
					when "01111100011100111" => rgb <= "000000";
					when "01111100011101000" => rgb <= "000000";
					when "01111100011101001" => rgb <= "000000";
					when "01111100011101010" => rgb <= "000000";
					when "01111100011101011" => rgb <= "000000";
					when "01111100011101100" => rgb <= "000000";
					when "01111100011101101" => rgb <= "000000";
					when "01111100011101110" => rgb <= "000000";
					when "01111100011101111" => rgb <= "000000";
					when "01111100011110000" => rgb <= "000000";
					when "01111100011110001" => rgb <= "000000";
					when "01111100011110010" => rgb <= "000000";
					when "01111100011110011" => rgb <= "000000";
					when "01111100011110100" => rgb <= "000000";
					when "01111100011110101" => rgb <= "000000";
					when "01111100011110110" => rgb <= "000000";
					when "01111100011110111" => rgb <= "000000";
					when "01111100011111000" => rgb <= "000000";
					when "01111100011111001" => rgb <= "000000";
					when "01111100011111010" => rgb <= "000000";
					when "01111100011111011" => rgb <= "000000";
					when "01111100011111100" => rgb <= "000000";
					when "01111100011111101" => rgb <= "000000";
					when "01111100011111110" => rgb <= "000000";
					when "01111100011111111" => rgb <= "000000";
					when "01111100100000000" => rgb <= "000000";
					when "01111100100000001" => rgb <= "000000";
					when "01111100100000010" => rgb <= "000000";
					when "01111100100000011" => rgb <= "000000";
					when "01111100100000100" => rgb <= "000000";
					when "01111100100000101" => rgb <= "000000";
					when "01111100100000110" => rgb <= "000000";
					when "01111100100000111" => rgb <= "000000";
					when "01111100100001000" => rgb <= "000000";
					when "01111100100001001" => rgb <= "000000";
					when "01111100100001010" => rgb <= "000000";
					when "01111100100001011" => rgb <= "000000";
					when "01111100100001100" => rgb <= "000000";
					when "01111100100001101" => rgb <= "000000";
					when "01111100100001110" => rgb <= "000000";
					when "01111100100001111" => rgb <= "000000";
					when "01111100100010000" => rgb <= "000000";
					when "01111100100010001" => rgb <= "000000";
					when "01111100100010010" => rgb <= "000000";
					when "01111100100010011" => rgb <= "000000";
					when "01111100100010100" => rgb <= "000000";
					when "01111100100010101" => rgb <= "000000";
					when "01111100100010110" => rgb <= "000000";
					when "01111100100010111" => rgb <= "000000";
					when "01111100100011000" => rgb <= "000000";
					when "01111100100011001" => rgb <= "000000";
					when "01111100100011010" => rgb <= "000000";
					when "01111100100011011" => rgb <= "000000";
					when "01111100100011100" => rgb <= "000000";
					when "01111100100011101" => rgb <= "000000";
					when "01111100100011110" => rgb <= "000000";
					when "01111100100011111" => rgb <= "000000";
					when "01111100100100000" => rgb <= "000000";
					when "01111100100100001" => rgb <= "000000";
					when "01111100100100010" => rgb <= "000000";
					when "01111100100100011" => rgb <= "000000";
					when "01111100100100100" => rgb <= "000000";
					when "01111100100100101" => rgb <= "000000";
					when "01111100100100110" => rgb <= "000000";
					when "01111100100100111" => rgb <= "000000";
					when "01111100100101000" => rgb <= "000000";
					when "01111100100101001" => rgb <= "000000";
					when "01111100100101010" => rgb <= "000000";
					when "01111100100101011" => rgb <= "000000";
					when "01111100100101100" => rgb <= "000000";
					when "01111100100101101" => rgb <= "000000";
					when "01111100100101110" => rgb <= "000000";
					when "01111100100101111" => rgb <= "000000";
					when "01111100100110000" => rgb <= "000000";
					when "01111100100110001" => rgb <= "000000";
					when "01111100100110010" => rgb <= "000000";
					when "01111100100110011" => rgb <= "000000";
					when "01111100100110100" => rgb <= "000000";
					when "01111100100110101" => rgb <= "000000";
					when "01111100100110110" => rgb <= "000000";
					when "01111100100110111" => rgb <= "000000";
					when "01111100100111000" => rgb <= "000000";
					when "01111100100111001" => rgb <= "000000";
					when "01111100100111010" => rgb <= "000000";
					when "01111100100111011" => rgb <= "000000";
					when "01111100100111100" => rgb <= "000000";
					when "01111100100111101" => rgb <= "000000";
					when "01111100100111110" => rgb <= "000000";
					when "01111100100111111" => rgb <= "000000";
					when "01111101000000000" => rgb <= "000000";
					when "01111101000000001" => rgb <= "000000";
					when "01111101000000010" => rgb <= "000000";
					when "01111101000000011" => rgb <= "000000";
					when "01111101000000100" => rgb <= "000000";
					when "01111101000000101" => rgb <= "000000";
					when "01111101000000110" => rgb <= "000000";
					when "01111101000000111" => rgb <= "000000";
					when "01111101000001000" => rgb <= "000000";
					when "01111101000001001" => rgb <= "000000";
					when "01111101000001010" => rgb <= "000000";
					when "01111101000001011" => rgb <= "000000";
					when "01111101000001100" => rgb <= "000000";
					when "01111101000001101" => rgb <= "000000";
					when "01111101000001110" => rgb <= "000000";
					when "01111101000001111" => rgb <= "000000";
					when "01111101000010000" => rgb <= "000000";
					when "01111101000010001" => rgb <= "000000";
					when "01111101000010010" => rgb <= "000000";
					when "01111101000010011" => rgb <= "000000";
					when "01111101000010100" => rgb <= "000000";
					when "01111101000010101" => rgb <= "000000";
					when "01111101000010110" => rgb <= "000000";
					when "01111101000010111" => rgb <= "000000";
					when "01111101000011000" => rgb <= "000000";
					when "01111101000011001" => rgb <= "000000";
					when "01111101000011010" => rgb <= "000000";
					when "01111101000011011" => rgb <= "000000";
					when "01111101000011100" => rgb <= "000000";
					when "01111101000011101" => rgb <= "000000";
					when "01111101000011110" => rgb <= "000000";
					when "01111101000011111" => rgb <= "000000";
					when "01111101000100000" => rgb <= "000000";
					when "01111101000100001" => rgb <= "000000";
					when "01111101000100010" => rgb <= "000000";
					when "01111101000100011" => rgb <= "000000";
					when "01111101000100100" => rgb <= "000000";
					when "01111101000100101" => rgb <= "000000";
					when "01111101000100110" => rgb <= "000000";
					when "01111101000100111" => rgb <= "000000";
					when "01111101000101000" => rgb <= "000000";
					when "01111101000101001" => rgb <= "000000";
					when "01111101000101010" => rgb <= "000000";
					when "01111101000101011" => rgb <= "000000";
					when "01111101000101100" => rgb <= "000000";
					when "01111101000101101" => rgb <= "000000";
					when "01111101000101110" => rgb <= "000000";
					when "01111101000101111" => rgb <= "000000";
					when "01111101000110000" => rgb <= "000000";
					when "01111101000110001" => rgb <= "000000";
					when "01111101000110010" => rgb <= "000000";
					when "01111101000110011" => rgb <= "000000";
					when "01111101000110100" => rgb <= "000000";
					when "01111101000110101" => rgb <= "000000";
					when "01111101000110110" => rgb <= "000000";
					when "01111101000110111" => rgb <= "000000";
					when "01111101000111000" => rgb <= "000000";
					when "01111101000111001" => rgb <= "000000";
					when "01111101000111010" => rgb <= "000000";
					when "01111101000111011" => rgb <= "000000";
					when "01111101000111100" => rgb <= "000000";
					when "01111101000111101" => rgb <= "000000";
					when "01111101000111110" => rgb <= "000000";
					when "01111101000111111" => rgb <= "000000";
					when "01111101001000000" => rgb <= "000000";
					when "01111101001000001" => rgb <= "000000";
					when "01111101001000010" => rgb <= "000000";
					when "01111101001000011" => rgb <= "000000";
					when "01111101001000100" => rgb <= "000000";
					when "01111101001000101" => rgb <= "000000";
					when "01111101001000110" => rgb <= "000000";
					when "01111101001000111" => rgb <= "000000";
					when "01111101001001000" => rgb <= "000000";
					when "01111101001001001" => rgb <= "000000";
					when "01111101001001010" => rgb <= "000000";
					when "01111101001001011" => rgb <= "000000";
					when "01111101001001100" => rgb <= "000000";
					when "01111101001001101" => rgb <= "000000";
					when "01111101001001110" => rgb <= "000000";
					when "01111101001001111" => rgb <= "000000";
					when "01111101001010000" => rgb <= "000000";
					when "01111101001010001" => rgb <= "000000";
					when "01111101001010010" => rgb <= "000000";
					when "01111101001010011" => rgb <= "000000";
					when "01111101001010100" => rgb <= "000000";
					when "01111101001010101" => rgb <= "000000";
					when "01111101001010110" => rgb <= "000000";
					when "01111101001010111" => rgb <= "000000";
					when "01111101001011000" => rgb <= "000000";
					when "01111101001011001" => rgb <= "000000";
					when "01111101001011010" => rgb <= "000000";
					when "01111101001011011" => rgb <= "000000";
					when "01111101001011100" => rgb <= "000000";
					when "01111101001011101" => rgb <= "000000";
					when "01111101001011110" => rgb <= "000000";
					when "01111101001011111" => rgb <= "000000";
					when "01111101001100000" => rgb <= "000000";
					when "01111101001100001" => rgb <= "000000";
					when "01111101001100010" => rgb <= "000000";
					when "01111101001100011" => rgb <= "000000";
					when "01111101001100100" => rgb <= "000000";
					when "01111101001100101" => rgb <= "000000";
					when "01111101001100110" => rgb <= "000000";
					when "01111101001100111" => rgb <= "000000";
					when "01111101001101000" => rgb <= "000000";
					when "01111101001101001" => rgb <= "000000";
					when "01111101001101010" => rgb <= "000000";
					when "01111101001101011" => rgb <= "000000";
					when "01111101001101100" => rgb <= "000000";
					when "01111101001101101" => rgb <= "000000";
					when "01111101001101110" => rgb <= "000000";
					when "01111101001101111" => rgb <= "000000";
					when "01111101001110000" => rgb <= "000000";
					when "01111101001110001" => rgb <= "000000";
					when "01111101001110010" => rgb <= "000000";
					when "01111101001110011" => rgb <= "000000";
					when "01111101001110100" => rgb <= "000000";
					when "01111101001110101" => rgb <= "000000";
					when "01111101001110110" => rgb <= "000000";
					when "01111101001110111" => rgb <= "000000";
					when "01111101001111000" => rgb <= "000000";
					when "01111101001111001" => rgb <= "000000";
					when "01111101001111010" => rgb <= "000000";
					when "01111101001111011" => rgb <= "000000";
					when "01111101001111100" => rgb <= "000000";
					when "01111101001111101" => rgb <= "000000";
					when "01111101001111110" => rgb <= "000000";
					when "01111101001111111" => rgb <= "000000";
					when "01111101010000000" => rgb <= "000000";
					when "01111101010000001" => rgb <= "000000";
					when "01111101010000010" => rgb <= "000000";
					when "01111101010000011" => rgb <= "000000";
					when "01111101010000100" => rgb <= "000000";
					when "01111101010000101" => rgb <= "000000";
					when "01111101010000110" => rgb <= "000000";
					when "01111101010000111" => rgb <= "000000";
					when "01111101010001000" => rgb <= "000000";
					when "01111101010001001" => rgb <= "000000";
					when "01111101010001010" => rgb <= "000000";
					when "01111101010001011" => rgb <= "000000";
					when "01111101010001100" => rgb <= "000000";
					when "01111101010001101" => rgb <= "000000";
					when "01111101010001110" => rgb <= "000000";
					when "01111101010001111" => rgb <= "000000";
					when "01111101010010000" => rgb <= "000000";
					when "01111101010010001" => rgb <= "000000";
					when "01111101010010010" => rgb <= "000000";
					when "01111101010010011" => rgb <= "000000";
					when "01111101010010100" => rgb <= "000000";
					when "01111101010010101" => rgb <= "000000";
					when "01111101010010110" => rgb <= "000000";
					when "01111101010010111" => rgb <= "000000";
					when "01111101010011000" => rgb <= "000000";
					when "01111101010011001" => rgb <= "000000";
					when "01111101010011010" => rgb <= "000000";
					when "01111101010011011" => rgb <= "000000";
					when "01111101010011100" => rgb <= "000000";
					when "01111101010011101" => rgb <= "000000";
					when "01111101010011110" => rgb <= "000000";
					when "01111101010011111" => rgb <= "000000";
					when "01111101010100000" => rgb <= "000000";
					when "01111101010100001" => rgb <= "000000";
					when "01111101010100010" => rgb <= "000000";
					when "01111101010100011" => rgb <= "000000";
					when "01111101010100100" => rgb <= "000000";
					when "01111101010100101" => rgb <= "000000";
					when "01111101010100110" => rgb <= "000000";
					when "01111101010100111" => rgb <= "000000";
					when "01111101010101000" => rgb <= "000000";
					when "01111101010101001" => rgb <= "000000";
					when "01111101010101010" => rgb <= "000000";
					when "01111101010101011" => rgb <= "000000";
					when "01111101010101100" => rgb <= "000000";
					when "01111101010101101" => rgb <= "000000";
					when "01111101010101110" => rgb <= "000000";
					when "01111101010101111" => rgb <= "000000";
					when "01111101010110000" => rgb <= "000000";
					when "01111101010110001" => rgb <= "000000";
					when "01111101010110010" => rgb <= "000000";
					when "01111101010110011" => rgb <= "000000";
					when "01111101010110100" => rgb <= "000000";
					when "01111101010110101" => rgb <= "000000";
					when "01111101010110110" => rgb <= "000000";
					when "01111101010110111" => rgb <= "000000";
					when "01111101010111000" => rgb <= "000000";
					when "01111101010111001" => rgb <= "000000";
					when "01111101010111010" => rgb <= "000000";
					when "01111101010111011" => rgb <= "000000";
					when "01111101010111100" => rgb <= "000000";
					when "01111101010111101" => rgb <= "000000";
					when "01111101010111110" => rgb <= "000000";
					when "01111101010111111" => rgb <= "000000";
					when "01111101011000000" => rgb <= "000000";
					when "01111101011000001" => rgb <= "000000";
					when "01111101011000010" => rgb <= "000000";
					when "01111101011000011" => rgb <= "000000";
					when "01111101011000100" => rgb <= "000000";
					when "01111101011000101" => rgb <= "000000";
					when "01111101011000110" => rgb <= "000000";
					when "01111101011000111" => rgb <= "000000";
					when "01111101011001000" => rgb <= "000000";
					when "01111101011001001" => rgb <= "000000";
					when "01111101011001010" => rgb <= "000000";
					when "01111101011001011" => rgb <= "000000";
					when "01111101011001100" => rgb <= "000000";
					when "01111101011001101" => rgb <= "000000";
					when "01111101011001110" => rgb <= "000000";
					when "01111101011001111" => rgb <= "000000";
					when "01111101011010000" => rgb <= "000000";
					when "01111101011010001" => rgb <= "000000";
					when "01111101011010010" => rgb <= "000000";
					when "01111101011010011" => rgb <= "000000";
					when "01111101011010100" => rgb <= "000000";
					when "01111101011010101" => rgb <= "000000";
					when "01111101011010110" => rgb <= "000000";
					when "01111101011010111" => rgb <= "000000";
					when "01111101011011000" => rgb <= "000000";
					when "01111101011011001" => rgb <= "000000";
					when "01111101011011010" => rgb <= "000000";
					when "01111101011011011" => rgb <= "000000";
					when "01111101011011100" => rgb <= "000000";
					when "01111101011011101" => rgb <= "000000";
					when "01111101011011110" => rgb <= "000000";
					when "01111101011011111" => rgb <= "000000";
					when "01111101011100000" => rgb <= "000000";
					when "01111101011100001" => rgb <= "000000";
					when "01111101011100010" => rgb <= "000000";
					when "01111101011100011" => rgb <= "000000";
					when "01111101011100100" => rgb <= "000000";
					when "01111101011100101" => rgb <= "000000";
					when "01111101011100110" => rgb <= "000000";
					when "01111101011100111" => rgb <= "000000";
					when "01111101011101000" => rgb <= "000000";
					when "01111101011101001" => rgb <= "000000";
					when "01111101011101010" => rgb <= "000000";
					when "01111101011101011" => rgb <= "000000";
					when "01111101011101100" => rgb <= "000000";
					when "01111101011101101" => rgb <= "000000";
					when "01111101011101110" => rgb <= "000000";
					when "01111101011101111" => rgb <= "000000";
					when "01111101011110000" => rgb <= "000000";
					when "01111101011110001" => rgb <= "000000";
					when "01111101011110010" => rgb <= "000000";
					when "01111101011110011" => rgb <= "000000";
					when "01111101011110100" => rgb <= "000000";
					when "01111101011110101" => rgb <= "000000";
					when "01111101011110110" => rgb <= "000000";
					when "01111101011110111" => rgb <= "000000";
					when "01111101011111000" => rgb <= "000000";
					when "01111101011111001" => rgb <= "000000";
					when "01111101011111010" => rgb <= "000000";
					when "01111101011111011" => rgb <= "000000";
					when "01111101011111100" => rgb <= "000000";
					when "01111101011111101" => rgb <= "000000";
					when "01111101011111110" => rgb <= "000000";
					when "01111101011111111" => rgb <= "000000";
					when "01111101100000000" => rgb <= "000000";
					when "01111101100000001" => rgb <= "000000";
					when "01111101100000010" => rgb <= "000000";
					when "01111101100000011" => rgb <= "000000";
					when "01111101100000100" => rgb <= "000000";
					when "01111101100000101" => rgb <= "000000";
					when "01111101100000110" => rgb <= "000000";
					when "01111101100000111" => rgb <= "000000";
					when "01111101100001000" => rgb <= "000000";
					when "01111101100001001" => rgb <= "000000";
					when "01111101100001010" => rgb <= "000000";
					when "01111101100001011" => rgb <= "000000";
					when "01111101100001100" => rgb <= "000000";
					when "01111101100001101" => rgb <= "000000";
					when "01111101100001110" => rgb <= "000000";
					when "01111101100001111" => rgb <= "000000";
					when "01111101100010000" => rgb <= "000000";
					when "01111101100010001" => rgb <= "000000";
					when "01111101100010010" => rgb <= "000000";
					when "01111101100010011" => rgb <= "000000";
					when "01111101100010100" => rgb <= "000000";
					when "01111101100010101" => rgb <= "000000";
					when "01111101100010110" => rgb <= "000000";
					when "01111101100010111" => rgb <= "000000";
					when "01111101100011000" => rgb <= "000000";
					when "01111101100011001" => rgb <= "000000";
					when "01111101100011010" => rgb <= "000000";
					when "01111101100011011" => rgb <= "000000";
					when "01111101100011100" => rgb <= "000000";
					when "01111101100011101" => rgb <= "000000";
					when "01111101100011110" => rgb <= "000000";
					when "01111101100011111" => rgb <= "000000";
					when "01111101100100000" => rgb <= "000000";
					when "01111101100100001" => rgb <= "000000";
					when "01111101100100010" => rgb <= "000000";
					when "01111101100100011" => rgb <= "000000";
					when "01111101100100100" => rgb <= "000000";
					when "01111101100100101" => rgb <= "000000";
					when "01111101100100110" => rgb <= "000000";
					when "01111101100100111" => rgb <= "000000";
					when "01111101100101000" => rgb <= "000000";
					when "01111101100101001" => rgb <= "000000";
					when "01111101100101010" => rgb <= "000000";
					when "01111101100101011" => rgb <= "000000";
					when "01111101100101100" => rgb <= "000000";
					when "01111101100101101" => rgb <= "000000";
					when "01111101100101110" => rgb <= "000000";
					when "01111101100101111" => rgb <= "000000";
					when "01111101100110000" => rgb <= "000000";
					when "01111101100110001" => rgb <= "000000";
					when "01111101100110010" => rgb <= "000000";
					when "01111101100110011" => rgb <= "000000";
					when "01111101100110100" => rgb <= "000000";
					when "01111101100110101" => rgb <= "000000";
					when "01111101100110110" => rgb <= "000000";
					when "01111101100110111" => rgb <= "000000";
					when "01111101100111000" => rgb <= "000000";
					when "01111101100111001" => rgb <= "000000";
					when "01111101100111010" => rgb <= "000000";
					when "01111101100111011" => rgb <= "000000";
					when "01111101100111100" => rgb <= "000000";
					when "01111101100111101" => rgb <= "000000";
					when "01111101100111110" => rgb <= "000000";
					when "01111101100111111" => rgb <= "000000";
					when "01111110000000000" => rgb <= "000000";
					when "01111110000000001" => rgb <= "000000";
					when "01111110000000010" => rgb <= "000000";
					when "01111110000000011" => rgb <= "000000";
					when "01111110000000100" => rgb <= "000000";
					when "01111110000000101" => rgb <= "000000";
					when "01111110000000110" => rgb <= "000000";
					when "01111110000000111" => rgb <= "000000";
					when "01111110000001000" => rgb <= "000000";
					when "01111110000001001" => rgb <= "000000";
					when "01111110000001010" => rgb <= "000000";
					when "01111110000001011" => rgb <= "000000";
					when "01111110000001100" => rgb <= "000000";
					when "01111110000001101" => rgb <= "000000";
					when "01111110000001110" => rgb <= "000000";
					when "01111110000001111" => rgb <= "000000";
					when "01111110000010000" => rgb <= "000000";
					when "01111110000010001" => rgb <= "000000";
					when "01111110000010010" => rgb <= "000000";
					when "01111110000010011" => rgb <= "000000";
					when "01111110000010100" => rgb <= "000000";
					when "01111110000010101" => rgb <= "000000";
					when "01111110000010110" => rgb <= "000000";
					when "01111110000010111" => rgb <= "000000";
					when "01111110000011000" => rgb <= "000000";
					when "01111110000011001" => rgb <= "000000";
					when "01111110000011010" => rgb <= "000000";
					when "01111110000011011" => rgb <= "000000";
					when "01111110000011100" => rgb <= "000000";
					when "01111110000011101" => rgb <= "000000";
					when "01111110000011110" => rgb <= "000000";
					when "01111110000011111" => rgb <= "000000";
					when "01111110000100000" => rgb <= "000000";
					when "01111110000100001" => rgb <= "000000";
					when "01111110000100010" => rgb <= "000000";
					when "01111110000100011" => rgb <= "000000";
					when "01111110000100100" => rgb <= "000000";
					when "01111110000100101" => rgb <= "000000";
					when "01111110000100110" => rgb <= "000000";
					when "01111110000100111" => rgb <= "000000";
					when "01111110000101000" => rgb <= "000000";
					when "01111110000101001" => rgb <= "000000";
					when "01111110000101010" => rgb <= "000000";
					when "01111110000101011" => rgb <= "000000";
					when "01111110000101100" => rgb <= "000000";
					when "01111110000101101" => rgb <= "000000";
					when "01111110000101110" => rgb <= "000000";
					when "01111110000101111" => rgb <= "000000";
					when "01111110000110000" => rgb <= "000000";
					when "01111110000110001" => rgb <= "000000";
					when "01111110000110010" => rgb <= "000000";
					when "01111110000110011" => rgb <= "000000";
					when "01111110000110100" => rgb <= "000000";
					when "01111110000110101" => rgb <= "000000";
					when "01111110000110110" => rgb <= "000000";
					when "01111110000110111" => rgb <= "000000";
					when "01111110000111000" => rgb <= "000000";
					when "01111110000111001" => rgb <= "000000";
					when "01111110000111010" => rgb <= "000000";
					when "01111110000111011" => rgb <= "000000";
					when "01111110000111100" => rgb <= "000000";
					when "01111110000111101" => rgb <= "000000";
					when "01111110000111110" => rgb <= "000000";
					when "01111110000111111" => rgb <= "000000";
					when "01111110001000000" => rgb <= "000000";
					when "01111110001000001" => rgb <= "000000";
					when "01111110001000010" => rgb <= "000000";
					when "01111110001000011" => rgb <= "000000";
					when "01111110001000100" => rgb <= "000000";
					when "01111110001000101" => rgb <= "000000";
					when "01111110001000110" => rgb <= "000000";
					when "01111110001000111" => rgb <= "000000";
					when "01111110001001000" => rgb <= "000000";
					when "01111110001001001" => rgb <= "000000";
					when "01111110001001010" => rgb <= "000000";
					when "01111110001001011" => rgb <= "000000";
					when "01111110001001100" => rgb <= "000000";
					when "01111110001001101" => rgb <= "000000";
					when "01111110001001110" => rgb <= "000000";
					when "01111110001001111" => rgb <= "000000";
					when "01111110001010000" => rgb <= "000000";
					when "01111110001010001" => rgb <= "000000";
					when "01111110001010010" => rgb <= "000000";
					when "01111110001010011" => rgb <= "000000";
					when "01111110001010100" => rgb <= "000000";
					when "01111110001010101" => rgb <= "000000";
					when "01111110001010110" => rgb <= "000000";
					when "01111110001010111" => rgb <= "000000";
					when "01111110001011000" => rgb <= "000000";
					when "01111110001011001" => rgb <= "000000";
					when "01111110001011010" => rgb <= "000000";
					when "01111110001011011" => rgb <= "000000";
					when "01111110001011100" => rgb <= "000000";
					when "01111110001011101" => rgb <= "000000";
					when "01111110001011110" => rgb <= "000000";
					when "01111110001011111" => rgb <= "000000";
					when "01111110001100000" => rgb <= "000000";
					when "01111110001100001" => rgb <= "000000";
					when "01111110001100010" => rgb <= "000000";
					when "01111110001100011" => rgb <= "000000";
					when "01111110001100100" => rgb <= "000000";
					when "01111110001100101" => rgb <= "000000";
					when "01111110001100110" => rgb <= "000000";
					when "01111110001100111" => rgb <= "000000";
					when "01111110001101000" => rgb <= "000000";
					when "01111110001101001" => rgb <= "000000";
					when "01111110001101010" => rgb <= "000000";
					when "01111110001101011" => rgb <= "000000";
					when "01111110001101100" => rgb <= "000000";
					when "01111110001101101" => rgb <= "000000";
					when "01111110001101110" => rgb <= "000000";
					when "01111110001101111" => rgb <= "000000";
					when "01111110001110000" => rgb <= "000000";
					when "01111110001110001" => rgb <= "000000";
					when "01111110001110010" => rgb <= "000000";
					when "01111110001110011" => rgb <= "000000";
					when "01111110001110100" => rgb <= "000000";
					when "01111110001110101" => rgb <= "000000";
					when "01111110001110110" => rgb <= "000000";
					when "01111110001110111" => rgb <= "000000";
					when "01111110001111000" => rgb <= "000000";
					when "01111110001111001" => rgb <= "000000";
					when "01111110001111010" => rgb <= "000000";
					when "01111110001111011" => rgb <= "000000";
					when "01111110001111100" => rgb <= "000000";
					when "01111110001111101" => rgb <= "000000";
					when "01111110001111110" => rgb <= "000000";
					when "01111110001111111" => rgb <= "000000";
					when "01111110010000000" => rgb <= "000000";
					when "01111110010000001" => rgb <= "000000";
					when "01111110010000010" => rgb <= "000000";
					when "01111110010000011" => rgb <= "000000";
					when "01111110010000100" => rgb <= "000000";
					when "01111110010000101" => rgb <= "000000";
					when "01111110010000110" => rgb <= "000000";
					when "01111110010000111" => rgb <= "000000";
					when "01111110010001000" => rgb <= "000000";
					when "01111110010001001" => rgb <= "000000";
					when "01111110010001010" => rgb <= "000000";
					when "01111110010001011" => rgb <= "000000";
					when "01111110010001100" => rgb <= "000000";
					when "01111110010001101" => rgb <= "000000";
					when "01111110010001110" => rgb <= "000000";
					when "01111110010001111" => rgb <= "000000";
					when "01111110010010000" => rgb <= "000000";
					when "01111110010010001" => rgb <= "000000";
					when "01111110010010010" => rgb <= "000000";
					when "01111110010010011" => rgb <= "000000";
					when "01111110010010100" => rgb <= "000000";
					when "01111110010010101" => rgb <= "000000";
					when "01111110010010110" => rgb <= "000000";
					when "01111110010010111" => rgb <= "000000";
					when "01111110010011000" => rgb <= "000000";
					when "01111110010011001" => rgb <= "000000";
					when "01111110010011010" => rgb <= "000000";
					when "01111110010011011" => rgb <= "000000";
					when "01111110010011100" => rgb <= "000000";
					when "01111110010011101" => rgb <= "000000";
					when "01111110010011110" => rgb <= "000000";
					when "01111110010011111" => rgb <= "000000";
					when "01111110010100000" => rgb <= "000000";
					when "01111110010100001" => rgb <= "000000";
					when "01111110010100010" => rgb <= "000000";
					when "01111110010100011" => rgb <= "000000";
					when "01111110010100100" => rgb <= "000000";
					when "01111110010100101" => rgb <= "000000";
					when "01111110010100110" => rgb <= "000000";
					when "01111110010100111" => rgb <= "000000";
					when "01111110010101000" => rgb <= "000000";
					when "01111110010101001" => rgb <= "000000";
					when "01111110010101010" => rgb <= "000000";
					when "01111110010101011" => rgb <= "000000";
					when "01111110010101100" => rgb <= "000000";
					when "01111110010101101" => rgb <= "000000";
					when "01111110010101110" => rgb <= "000000";
					when "01111110010101111" => rgb <= "000000";
					when "01111110010110000" => rgb <= "000000";
					when "01111110010110001" => rgb <= "000000";
					when "01111110010110010" => rgb <= "000000";
					when "01111110010110011" => rgb <= "000000";
					when "01111110010110100" => rgb <= "000000";
					when "01111110010110101" => rgb <= "000000";
					when "01111110010110110" => rgb <= "000000";
					when "01111110010110111" => rgb <= "000000";
					when "01111110010111000" => rgb <= "000000";
					when "01111110010111001" => rgb <= "000000";
					when "01111110010111010" => rgb <= "000000";
					when "01111110010111011" => rgb <= "000000";
					when "01111110010111100" => rgb <= "000000";
					when "01111110010111101" => rgb <= "000000";
					when "01111110010111110" => rgb <= "000000";
					when "01111110010111111" => rgb <= "000000";
					when "01111110011000000" => rgb <= "000000";
					when "01111110011000001" => rgb <= "000000";
					when "01111110011000010" => rgb <= "000000";
					when "01111110011000011" => rgb <= "000000";
					when "01111110011000100" => rgb <= "000000";
					when "01111110011000101" => rgb <= "000000";
					when "01111110011000110" => rgb <= "000000";
					when "01111110011000111" => rgb <= "000000";
					when "01111110011001000" => rgb <= "000000";
					when "01111110011001001" => rgb <= "000000";
					when "01111110011001010" => rgb <= "000000";
					when "01111110011001011" => rgb <= "000000";
					when "01111110011001100" => rgb <= "000000";
					when "01111110011001101" => rgb <= "000000";
					when "01111110011001110" => rgb <= "000000";
					when "01111110011001111" => rgb <= "000000";
					when "01111110011010000" => rgb <= "000000";
					when "01111110011010001" => rgb <= "000000";
					when "01111110011010010" => rgb <= "000000";
					when "01111110011010011" => rgb <= "000000";
					when "01111110011010100" => rgb <= "000000";
					when "01111110011010101" => rgb <= "000000";
					when "01111110011010110" => rgb <= "000000";
					when "01111110011010111" => rgb <= "000000";
					when "01111110011011000" => rgb <= "000000";
					when "01111110011011001" => rgb <= "000000";
					when "01111110011011010" => rgb <= "000000";
					when "01111110011011011" => rgb <= "000000";
					when "01111110011011100" => rgb <= "000000";
					when "01111110011011101" => rgb <= "000000";
					when "01111110011011110" => rgb <= "000000";
					when "01111110011011111" => rgb <= "000000";
					when "01111110011100000" => rgb <= "000000";
					when "01111110011100001" => rgb <= "000000";
					when "01111110011100010" => rgb <= "000000";
					when "01111110011100011" => rgb <= "000000";
					when "01111110011100100" => rgb <= "000000";
					when "01111110011100101" => rgb <= "000000";
					when "01111110011100110" => rgb <= "000000";
					when "01111110011100111" => rgb <= "000000";
					when "01111110011101000" => rgb <= "000000";
					when "01111110011101001" => rgb <= "000000";
					when "01111110011101010" => rgb <= "000000";
					when "01111110011101011" => rgb <= "000000";
					when "01111110011101100" => rgb <= "000000";
					when "01111110011101101" => rgb <= "000000";
					when "01111110011101110" => rgb <= "000000";
					when "01111110011101111" => rgb <= "000000";
					when "01111110011110000" => rgb <= "000000";
					when "01111110011110001" => rgb <= "000000";
					when "01111110011110010" => rgb <= "000000";
					when "01111110011110011" => rgb <= "000000";
					when "01111110011110100" => rgb <= "000000";
					when "01111110011110101" => rgb <= "000000";
					when "01111110011110110" => rgb <= "000000";
					when "01111110011110111" => rgb <= "000000";
					when "01111110011111000" => rgb <= "000000";
					when "01111110011111001" => rgb <= "000000";
					when "01111110011111010" => rgb <= "000000";
					when "01111110011111011" => rgb <= "000000";
					when "01111110011111100" => rgb <= "000000";
					when "01111110011111101" => rgb <= "000000";
					when "01111110011111110" => rgb <= "000000";
					when "01111110011111111" => rgb <= "000000";
					when "01111110100000000" => rgb <= "000000";
					when "01111110100000001" => rgb <= "000000";
					when "01111110100000010" => rgb <= "000000";
					when "01111110100000011" => rgb <= "000000";
					when "01111110100000100" => rgb <= "000000";
					when "01111110100000101" => rgb <= "000000";
					when "01111110100000110" => rgb <= "000000";
					when "01111110100000111" => rgb <= "000000";
					when "01111110100001000" => rgb <= "000000";
					when "01111110100001001" => rgb <= "000000";
					when "01111110100001010" => rgb <= "000000";
					when "01111110100001011" => rgb <= "000000";
					when "01111110100001100" => rgb <= "000000";
					when "01111110100001101" => rgb <= "000000";
					when "01111110100001110" => rgb <= "000000";
					when "01111110100001111" => rgb <= "000000";
					when "01111110100010000" => rgb <= "000000";
					when "01111110100010001" => rgb <= "000000";
					when "01111110100010010" => rgb <= "000000";
					when "01111110100010011" => rgb <= "000000";
					when "01111110100010100" => rgb <= "000000";
					when "01111110100010101" => rgb <= "000000";
					when "01111110100010110" => rgb <= "000000";
					when "01111110100010111" => rgb <= "000000";
					when "01111110100011000" => rgb <= "000000";
					when "01111110100011001" => rgb <= "000000";
					when "01111110100011010" => rgb <= "000000";
					when "01111110100011011" => rgb <= "000000";
					when "01111110100011100" => rgb <= "000000";
					when "01111110100011101" => rgb <= "000000";
					when "01111110100011110" => rgb <= "000000";
					when "01111110100011111" => rgb <= "000000";
					when "01111110100100000" => rgb <= "000000";
					when "01111110100100001" => rgb <= "000000";
					when "01111110100100010" => rgb <= "000000";
					when "01111110100100011" => rgb <= "000000";
					when "01111110100100100" => rgb <= "000000";
					when "01111110100100101" => rgb <= "000000";
					when "01111110100100110" => rgb <= "000000";
					when "01111110100100111" => rgb <= "000000";
					when "01111110100101000" => rgb <= "000000";
					when "01111110100101001" => rgb <= "000000";
					when "01111110100101010" => rgb <= "000000";
					when "01111110100101011" => rgb <= "000000";
					when "01111110100101100" => rgb <= "000000";
					when "01111110100101101" => rgb <= "000000";
					when "01111110100101110" => rgb <= "000000";
					when "01111110100101111" => rgb <= "000000";
					when "01111110100110000" => rgb <= "000000";
					when "01111110100110001" => rgb <= "000000";
					when "01111110100110010" => rgb <= "000000";
					when "01111110100110011" => rgb <= "000000";
					when "01111110100110100" => rgb <= "000000";
					when "01111110100110101" => rgb <= "000000";
					when "01111110100110110" => rgb <= "000000";
					when "01111110100110111" => rgb <= "000000";
					when "01111110100111000" => rgb <= "000000";
					when "01111110100111001" => rgb <= "000000";
					when "01111110100111010" => rgb <= "000000";
					when "01111110100111011" => rgb <= "000000";
					when "01111110100111100" => rgb <= "000000";
					when "01111110100111101" => rgb <= "000000";
					when "01111110100111110" => rgb <= "000000";
					when "01111110100111111" => rgb <= "000000";
					when "01111111000000000" => rgb <= "000000";
					when "01111111000000001" => rgb <= "000000";
					when "01111111000000010" => rgb <= "000000";
					when "01111111000000011" => rgb <= "000000";
					when "01111111000000100" => rgb <= "000000";
					when "01111111000000101" => rgb <= "000000";
					when "01111111000000110" => rgb <= "000000";
					when "01111111000000111" => rgb <= "000000";
					when "01111111000001000" => rgb <= "000000";
					when "01111111000001001" => rgb <= "000000";
					when "01111111000001010" => rgb <= "000000";
					when "01111111000001011" => rgb <= "000000";
					when "01111111000001100" => rgb <= "000000";
					when "01111111000001101" => rgb <= "000000";
					when "01111111000001110" => rgb <= "000000";
					when "01111111000001111" => rgb <= "000000";
					when "01111111000010000" => rgb <= "000000";
					when "01111111000010001" => rgb <= "000000";
					when "01111111000010010" => rgb <= "000000";
					when "01111111000010011" => rgb <= "000000";
					when "01111111000010100" => rgb <= "000000";
					when "01111111000010101" => rgb <= "000000";
					when "01111111000010110" => rgb <= "000000";
					when "01111111000010111" => rgb <= "000000";
					when "01111111000011000" => rgb <= "000000";
					when "01111111000011001" => rgb <= "000000";
					when "01111111000011010" => rgb <= "000000";
					when "01111111000011011" => rgb <= "000000";
					when "01111111000011100" => rgb <= "000000";
					when "01111111000011101" => rgb <= "000000";
					when "01111111000011110" => rgb <= "000000";
					when "01111111000011111" => rgb <= "000000";
					when "01111111000100000" => rgb <= "000000";
					when "01111111000100001" => rgb <= "000000";
					when "01111111000100010" => rgb <= "000000";
					when "01111111000100011" => rgb <= "000000";
					when "01111111000100100" => rgb <= "000000";
					when "01111111000100101" => rgb <= "000000";
					when "01111111000100110" => rgb <= "000000";
					when "01111111000100111" => rgb <= "000000";
					when "01111111000101000" => rgb <= "000000";
					when "01111111000101001" => rgb <= "000000";
					when "01111111000101010" => rgb <= "000000";
					when "01111111000101011" => rgb <= "000000";
					when "01111111000101100" => rgb <= "000000";
					when "01111111000101101" => rgb <= "000000";
					when "01111111000101110" => rgb <= "000000";
					when "01111111000101111" => rgb <= "000000";
					when "01111111000110000" => rgb <= "000000";
					when "01111111000110001" => rgb <= "000000";
					when "01111111000110010" => rgb <= "000000";
					when "01111111000110011" => rgb <= "000000";
					when "01111111000110100" => rgb <= "000000";
					when "01111111000110101" => rgb <= "000000";
					when "01111111000110110" => rgb <= "000000";
					when "01111111000110111" => rgb <= "000000";
					when "01111111000111000" => rgb <= "000000";
					when "01111111000111001" => rgb <= "000000";
					when "01111111000111010" => rgb <= "000000";
					when "01111111000111011" => rgb <= "000000";
					when "01111111000111100" => rgb <= "000000";
					when "01111111000111101" => rgb <= "000000";
					when "01111111000111110" => rgb <= "000000";
					when "01111111000111111" => rgb <= "000000";
					when "01111111001000000" => rgb <= "000000";
					when "01111111001000001" => rgb <= "000000";
					when "01111111001000010" => rgb <= "000000";
					when "01111111001000011" => rgb <= "000000";
					when "01111111001000100" => rgb <= "000000";
					when "01111111001000101" => rgb <= "000000";
					when "01111111001000110" => rgb <= "000000";
					when "01111111001000111" => rgb <= "000000";
					when "01111111001001000" => rgb <= "000000";
					when "01111111001001001" => rgb <= "000000";
					when "01111111001001010" => rgb <= "000000";
					when "01111111001001011" => rgb <= "000000";
					when "01111111001001100" => rgb <= "000000";
					when "01111111001001101" => rgb <= "000000";
					when "01111111001001110" => rgb <= "000000";
					when "01111111001001111" => rgb <= "000000";
					when "01111111001010000" => rgb <= "000000";
					when "01111111001010001" => rgb <= "000000";
					when "01111111001010010" => rgb <= "000000";
					when "01111111001010011" => rgb <= "000000";
					when "01111111001010100" => rgb <= "000000";
					when "01111111001010101" => rgb <= "000000";
					when "01111111001010110" => rgb <= "000000";
					when "01111111001010111" => rgb <= "000000";
					when "01111111001011000" => rgb <= "000000";
					when "01111111001011001" => rgb <= "000000";
					when "01111111001011010" => rgb <= "000000";
					when "01111111001011011" => rgb <= "000000";
					when "01111111001011100" => rgb <= "000000";
					when "01111111001011101" => rgb <= "000000";
					when "01111111001011110" => rgb <= "000000";
					when "01111111001011111" => rgb <= "000000";
					when "01111111001100000" => rgb <= "000000";
					when "01111111001100001" => rgb <= "000000";
					when "01111111001100010" => rgb <= "000000";
					when "01111111001100011" => rgb <= "000000";
					when "01111111001100100" => rgb <= "000000";
					when "01111111001100101" => rgb <= "000000";
					when "01111111001100110" => rgb <= "000000";
					when "01111111001100111" => rgb <= "000000";
					when "01111111001101000" => rgb <= "000000";
					when "01111111001101001" => rgb <= "000000";
					when "01111111001101010" => rgb <= "000000";
					when "01111111001101011" => rgb <= "000000";
					when "01111111001101100" => rgb <= "000000";
					when "01111111001101101" => rgb <= "000000";
					when "01111111001101110" => rgb <= "000000";
					when "01111111001101111" => rgb <= "000000";
					when "01111111001110000" => rgb <= "000000";
					when "01111111001110001" => rgb <= "000000";
					when "01111111001110010" => rgb <= "000000";
					when "01111111001110011" => rgb <= "000000";
					when "01111111001110100" => rgb <= "000000";
					when "01111111001110101" => rgb <= "000000";
					when "01111111001110110" => rgb <= "000000";
					when "01111111001110111" => rgb <= "000000";
					when "01111111001111000" => rgb <= "000000";
					when "01111111001111001" => rgb <= "000000";
					when "01111111001111010" => rgb <= "000000";
					when "01111111001111011" => rgb <= "000000";
					when "01111111001111100" => rgb <= "000000";
					when "01111111001111101" => rgb <= "000000";
					when "01111111001111110" => rgb <= "000000";
					when "01111111001111111" => rgb <= "000000";
					when "01111111010000000" => rgb <= "000000";
					when "01111111010000001" => rgb <= "000000";
					when "01111111010000010" => rgb <= "000000";
					when "01111111010000011" => rgb <= "000000";
					when "01111111010000100" => rgb <= "000000";
					when "01111111010000101" => rgb <= "000000";
					when "01111111010000110" => rgb <= "000000";
					when "01111111010000111" => rgb <= "000000";
					when "01111111010001000" => rgb <= "000000";
					when "01111111010001001" => rgb <= "000000";
					when "01111111010001010" => rgb <= "000000";
					when "01111111010001011" => rgb <= "000000";
					when "01111111010001100" => rgb <= "000000";
					when "01111111010001101" => rgb <= "000000";
					when "01111111010001110" => rgb <= "000000";
					when "01111111010001111" => rgb <= "000000";
					when "01111111010010000" => rgb <= "000000";
					when "01111111010010001" => rgb <= "000000";
					when "01111111010010010" => rgb <= "000000";
					when "01111111010010011" => rgb <= "000000";
					when "01111111010010100" => rgb <= "000000";
					when "01111111010010101" => rgb <= "000000";
					when "01111111010010110" => rgb <= "000000";
					when "01111111010010111" => rgb <= "000000";
					when "01111111010011000" => rgb <= "000000";
					when "01111111010011001" => rgb <= "000000";
					when "01111111010011010" => rgb <= "000000";
					when "01111111010011011" => rgb <= "000000";
					when "01111111010011100" => rgb <= "000000";
					when "01111111010011101" => rgb <= "000000";
					when "01111111010011110" => rgb <= "000000";
					when "01111111010011111" => rgb <= "000000";
					when "01111111010100000" => rgb <= "000000";
					when "01111111010100001" => rgb <= "000000";
					when "01111111010100010" => rgb <= "000000";
					when "01111111010100011" => rgb <= "000000";
					when "01111111010100100" => rgb <= "000000";
					when "01111111010100101" => rgb <= "000000";
					when "01111111010100110" => rgb <= "000000";
					when "01111111010100111" => rgb <= "000000";
					when "01111111010101000" => rgb <= "000000";
					when "01111111010101001" => rgb <= "000000";
					when "01111111010101010" => rgb <= "000000";
					when "01111111010101011" => rgb <= "000000";
					when "01111111010101100" => rgb <= "000000";
					when "01111111010101101" => rgb <= "000000";
					when "01111111010101110" => rgb <= "000000";
					when "01111111010101111" => rgb <= "000000";
					when "01111111010110000" => rgb <= "000000";
					when "01111111010110001" => rgb <= "000000";
					when "01111111010110010" => rgb <= "000000";
					when "01111111010110011" => rgb <= "000000";
					when "01111111010110100" => rgb <= "000000";
					when "01111111010110101" => rgb <= "000000";
					when "01111111010110110" => rgb <= "000000";
					when "01111111010110111" => rgb <= "000000";
					when "01111111010111000" => rgb <= "000000";
					when "01111111010111001" => rgb <= "000000";
					when "01111111010111010" => rgb <= "000000";
					when "01111111010111011" => rgb <= "000000";
					when "01111111010111100" => rgb <= "000000";
					when "01111111010111101" => rgb <= "000000";
					when "01111111010111110" => rgb <= "000000";
					when "01111111010111111" => rgb <= "000000";
					when "01111111011000000" => rgb <= "000000";
					when "01111111011000001" => rgb <= "000000";
					when "01111111011000010" => rgb <= "000000";
					when "01111111011000011" => rgb <= "000000";
					when "01111111011000100" => rgb <= "000000";
					when "01111111011000101" => rgb <= "000000";
					when "01111111011000110" => rgb <= "000000";
					when "01111111011000111" => rgb <= "000000";
					when "01111111011001000" => rgb <= "000000";
					when "01111111011001001" => rgb <= "000000";
					when "01111111011001010" => rgb <= "000000";
					when "01111111011001011" => rgb <= "000000";
					when "01111111011001100" => rgb <= "000000";
					when "01111111011001101" => rgb <= "000000";
					when "01111111011001110" => rgb <= "000000";
					when "01111111011001111" => rgb <= "000000";
					when "01111111011010000" => rgb <= "000000";
					when "01111111011010001" => rgb <= "000000";
					when "01111111011010010" => rgb <= "000000";
					when "01111111011010011" => rgb <= "000000";
					when "01111111011010100" => rgb <= "000000";
					when "01111111011010101" => rgb <= "000000";
					when "01111111011010110" => rgb <= "000000";
					when "01111111011010111" => rgb <= "000000";
					when "01111111011011000" => rgb <= "000000";
					when "01111111011011001" => rgb <= "000000";
					when "01111111011011010" => rgb <= "000000";
					when "01111111011011011" => rgb <= "000000";
					when "01111111011011100" => rgb <= "000000";
					when "01111111011011101" => rgb <= "000000";
					when "01111111011011110" => rgb <= "000000";
					when "01111111011011111" => rgb <= "000000";
					when "01111111011100000" => rgb <= "000000";
					when "01111111011100001" => rgb <= "000000";
					when "01111111011100010" => rgb <= "000000";
					when "01111111011100011" => rgb <= "000000";
					when "01111111011100100" => rgb <= "000000";
					when "01111111011100101" => rgb <= "000000";
					when "01111111011100110" => rgb <= "000000";
					when "01111111011100111" => rgb <= "000000";
					when "01111111011101000" => rgb <= "000000";
					when "01111111011101001" => rgb <= "000000";
					when "01111111011101010" => rgb <= "000000";
					when "01111111011101011" => rgb <= "000000";
					when "01111111011101100" => rgb <= "000000";
					when "01111111011101101" => rgb <= "000000";
					when "01111111011101110" => rgb <= "000000";
					when "01111111011101111" => rgb <= "000000";
					when "01111111011110000" => rgb <= "000000";
					when "01111111011110001" => rgb <= "000000";
					when "01111111011110010" => rgb <= "000000";
					when "01111111011110011" => rgb <= "000000";
					when "01111111011110100" => rgb <= "000000";
					when "01111111011110101" => rgb <= "000000";
					when "01111111011110110" => rgb <= "000000";
					when "01111111011110111" => rgb <= "000000";
					when "01111111011111000" => rgb <= "000000";
					when "01111111011111001" => rgb <= "000000";
					when "01111111011111010" => rgb <= "000000";
					when "01111111011111011" => rgb <= "000000";
					when "01111111011111100" => rgb <= "000000";
					when "01111111011111101" => rgb <= "000000";
					when "01111111011111110" => rgb <= "000000";
					when "01111111011111111" => rgb <= "000000";
					when "01111111100000000" => rgb <= "000000";
					when "01111111100000001" => rgb <= "000000";
					when "01111111100000010" => rgb <= "000000";
					when "01111111100000011" => rgb <= "000000";
					when "01111111100000100" => rgb <= "000000";
					when "01111111100000101" => rgb <= "000000";
					when "01111111100000110" => rgb <= "000000";
					when "01111111100000111" => rgb <= "000000";
					when "01111111100001000" => rgb <= "000000";
					when "01111111100001001" => rgb <= "000000";
					when "01111111100001010" => rgb <= "000000";
					when "01111111100001011" => rgb <= "000000";
					when "01111111100001100" => rgb <= "000000";
					when "01111111100001101" => rgb <= "000000";
					when "01111111100001110" => rgb <= "000000";
					when "01111111100001111" => rgb <= "000000";
					when "01111111100010000" => rgb <= "000000";
					when "01111111100010001" => rgb <= "000000";
					when "01111111100010010" => rgb <= "000000";
					when "01111111100010011" => rgb <= "000000";
					when "01111111100010100" => rgb <= "000000";
					when "01111111100010101" => rgb <= "000000";
					when "01111111100010110" => rgb <= "000000";
					when "01111111100010111" => rgb <= "000000";
					when "01111111100011000" => rgb <= "000000";
					when "01111111100011001" => rgb <= "000000";
					when "01111111100011010" => rgb <= "000000";
					when "01111111100011011" => rgb <= "000000";
					when "01111111100011100" => rgb <= "000000";
					when "01111111100011101" => rgb <= "000000";
					when "01111111100011110" => rgb <= "000000";
					when "01111111100011111" => rgb <= "000000";
					when "01111111100100000" => rgb <= "000000";
					when "01111111100100001" => rgb <= "000000";
					when "01111111100100010" => rgb <= "000000";
					when "01111111100100011" => rgb <= "000000";
					when "01111111100100100" => rgb <= "000000";
					when "01111111100100101" => rgb <= "000000";
					when "01111111100100110" => rgb <= "000000";
					when "01111111100100111" => rgb <= "000000";
					when "01111111100101000" => rgb <= "000000";
					when "01111111100101001" => rgb <= "000000";
					when "01111111100101010" => rgb <= "000000";
					when "01111111100101011" => rgb <= "000000";
					when "01111111100101100" => rgb <= "000000";
					when "01111111100101101" => rgb <= "000000";
					when "01111111100101110" => rgb <= "000000";
					when "01111111100101111" => rgb <= "000000";
					when "01111111100110000" => rgb <= "000000";
					when "01111111100110001" => rgb <= "000000";
					when "01111111100110010" => rgb <= "000000";
					when "01111111100110011" => rgb <= "000000";
					when "01111111100110100" => rgb <= "000000";
					when "01111111100110101" => rgb <= "000000";
					when "01111111100110110" => rgb <= "000000";
					when "01111111100110111" => rgb <= "000000";
					when "01111111100111000" => rgb <= "000000";
					when "01111111100111001" => rgb <= "000000";
					when "01111111100111010" => rgb <= "000000";
					when "01111111100111011" => rgb <= "000000";
					when "01111111100111100" => rgb <= "000000";
					when "01111111100111101" => rgb <= "000000";
					when "01111111100111110" => rgb <= "000000";
					when "01111111100111111" => rgb <= "000000";
					when "10000000000000000" => rgb <= "000000";
					when "10000000000000001" => rgb <= "000000";
					when "10000000000000010" => rgb <= "000000";
					when "10000000000000011" => rgb <= "000000";
					when "10000000000000100" => rgb <= "000000";
					when "10000000000000101" => rgb <= "000000";
					when "10000000000000110" => rgb <= "000000";
					when "10000000000000111" => rgb <= "000000";
					when "10000000000001000" => rgb <= "000000";
					when "10000000000001001" => rgb <= "000000";
					when "10000000000001010" => rgb <= "000000";
					when "10000000000001011" => rgb <= "000000";
					when "10000000000001100" => rgb <= "000000";
					when "10000000000001101" => rgb <= "000000";
					when "10000000000001110" => rgb <= "000000";
					when "10000000000001111" => rgb <= "000000";
					when "10000000000010000" => rgb <= "000000";
					when "10000000000010001" => rgb <= "000000";
					when "10000000000010010" => rgb <= "000000";
					when "10000000000010011" => rgb <= "000000";
					when "10000000000010100" => rgb <= "000000";
					when "10000000000010101" => rgb <= "000000";
					when "10000000000010110" => rgb <= "000000";
					when "10000000000010111" => rgb <= "000000";
					when "10000000000011000" => rgb <= "000000";
					when "10000000000011001" => rgb <= "000000";
					when "10000000000011010" => rgb <= "000000";
					when "10000000000011011" => rgb <= "000000";
					when "10000000000011100" => rgb <= "000000";
					when "10000000000011101" => rgb <= "000000";
					when "10000000000011110" => rgb <= "000000";
					when "10000000000011111" => rgb <= "000000";
					when "10000000000100000" => rgb <= "000000";
					when "10000000000100001" => rgb <= "000000";
					when "10000000000100010" => rgb <= "000000";
					when "10000000000100011" => rgb <= "000000";
					when "10000000000100100" => rgb <= "000000";
					when "10000000000100101" => rgb <= "000000";
					when "10000000000100110" => rgb <= "000000";
					when "10000000000100111" => rgb <= "000000";
					when "10000000000101000" => rgb <= "000000";
					when "10000000000101001" => rgb <= "000000";
					when "10000000000101010" => rgb <= "000000";
					when "10000000000101011" => rgb <= "000000";
					when "10000000000101100" => rgb <= "000000";
					when "10000000000101101" => rgb <= "000000";
					when "10000000000101110" => rgb <= "000000";
					when "10000000000101111" => rgb <= "000000";
					when "10000000000110000" => rgb <= "000000";
					when "10000000000110001" => rgb <= "000000";
					when "10000000000110010" => rgb <= "000000";
					when "10000000000110011" => rgb <= "000000";
					when "10000000000110100" => rgb <= "000000";
					when "10000000000110101" => rgb <= "000000";
					when "10000000000110110" => rgb <= "000000";
					when "10000000000110111" => rgb <= "000000";
					when "10000000000111000" => rgb <= "000000";
					when "10000000000111001" => rgb <= "000000";
					when "10000000000111010" => rgb <= "000000";
					when "10000000000111011" => rgb <= "000000";
					when "10000000000111100" => rgb <= "000000";
					when "10000000000111101" => rgb <= "000000";
					when "10000000000111110" => rgb <= "000000";
					when "10000000000111111" => rgb <= "000000";
					when "10000000001000000" => rgb <= "000000";
					when "10000000001000001" => rgb <= "000000";
					when "10000000001000010" => rgb <= "000000";
					when "10000000001000011" => rgb <= "000000";
					when "10000000001000100" => rgb <= "000000";
					when "10000000001000101" => rgb <= "000000";
					when "10000000001000110" => rgb <= "000000";
					when "10000000001000111" => rgb <= "000000";
					when "10000000001001000" => rgb <= "000000";
					when "10000000001001001" => rgb <= "000000";
					when "10000000001001010" => rgb <= "000000";
					when "10000000001001011" => rgb <= "000000";
					when "10000000001001100" => rgb <= "000000";
					when "10000000001001101" => rgb <= "000000";
					when "10000000001001110" => rgb <= "000000";
					when "10000000001001111" => rgb <= "000000";
					when "10000000001010000" => rgb <= "000000";
					when "10000000001010001" => rgb <= "000000";
					when "10000000001010010" => rgb <= "000000";
					when "10000000001010011" => rgb <= "000000";
					when "10000000001010100" => rgb <= "000000";
					when "10000000001010101" => rgb <= "000000";
					when "10000000001010110" => rgb <= "000000";
					when "10000000001010111" => rgb <= "000000";
					when "10000000001011000" => rgb <= "000000";
					when "10000000001011001" => rgb <= "000000";
					when "10000000001011010" => rgb <= "000000";
					when "10000000001011011" => rgb <= "000000";
					when "10000000001011100" => rgb <= "000000";
					when "10000000001011101" => rgb <= "000000";
					when "10000000001011110" => rgb <= "000000";
					when "10000000001011111" => rgb <= "000000";
					when "10000000001100000" => rgb <= "000000";
					when "10000000001100001" => rgb <= "000000";
					when "10000000001100010" => rgb <= "000000";
					when "10000000001100011" => rgb <= "000000";
					when "10000000001100100" => rgb <= "000000";
					when "10000000001100101" => rgb <= "000000";
					when "10000000001100110" => rgb <= "000000";
					when "10000000001100111" => rgb <= "000000";
					when "10000000001101000" => rgb <= "000000";
					when "10000000001101001" => rgb <= "000000";
					when "10000000001101010" => rgb <= "000000";
					when "10000000001101011" => rgb <= "000000";
					when "10000000001101100" => rgb <= "000000";
					when "10000000001101101" => rgb <= "000000";
					when "10000000001101110" => rgb <= "000000";
					when "10000000001101111" => rgb <= "000000";
					when "10000000001110000" => rgb <= "000000";
					when "10000000001110001" => rgb <= "000000";
					when "10000000001110010" => rgb <= "000000";
					when "10000000001110011" => rgb <= "000000";
					when "10000000001110100" => rgb <= "000000";
					when "10000000001110101" => rgb <= "000000";
					when "10000000001110110" => rgb <= "000000";
					when "10000000001110111" => rgb <= "000000";
					when "10000000001111000" => rgb <= "000000";
					when "10000000001111001" => rgb <= "000000";
					when "10000000001111010" => rgb <= "000000";
					when "10000000001111011" => rgb <= "000000";
					when "10000000001111100" => rgb <= "000000";
					when "10000000001111101" => rgb <= "000000";
					when "10000000001111110" => rgb <= "000000";
					when "10000000001111111" => rgb <= "000000";
					when "10000000010000000" => rgb <= "000000";
					when "10000000010000001" => rgb <= "000000";
					when "10000000010000010" => rgb <= "000000";
					when "10000000010000011" => rgb <= "000000";
					when "10000000010000100" => rgb <= "000000";
					when "10000000010000101" => rgb <= "000000";
					when "10000000010000110" => rgb <= "000000";
					when "10000000010000111" => rgb <= "000000";
					when "10000000010001000" => rgb <= "000000";
					when "10000000010001001" => rgb <= "000000";
					when "10000000010001010" => rgb <= "000000";
					when "10000000010001011" => rgb <= "000000";
					when "10000000010001100" => rgb <= "000000";
					when "10000000010001101" => rgb <= "000000";
					when "10000000010001110" => rgb <= "000000";
					when "10000000010001111" => rgb <= "000000";
					when "10000000010010000" => rgb <= "000000";
					when "10000000010010001" => rgb <= "000000";
					when "10000000010010010" => rgb <= "000000";
					when "10000000010010011" => rgb <= "000000";
					when "10000000010010100" => rgb <= "000000";
					when "10000000010010101" => rgb <= "000000";
					when "10000000010010110" => rgb <= "000000";
					when "10000000010010111" => rgb <= "000000";
					when "10000000010011000" => rgb <= "000000";
					when "10000000010011001" => rgb <= "000000";
					when "10000000010011010" => rgb <= "000000";
					when "10000000010011011" => rgb <= "000000";
					when "10000000010011100" => rgb <= "000000";
					when "10000000010011101" => rgb <= "000000";
					when "10000000010011110" => rgb <= "000000";
					when "10000000010011111" => rgb <= "000000";
					when "10000000010100000" => rgb <= "000000";
					when "10000000010100001" => rgb <= "000000";
					when "10000000010100010" => rgb <= "000000";
					when "10000000010100011" => rgb <= "000000";
					when "10000000010100100" => rgb <= "000000";
					when "10000000010100101" => rgb <= "000000";
					when "10000000010100110" => rgb <= "000000";
					when "10000000010100111" => rgb <= "000000";
					when "10000000010101000" => rgb <= "000000";
					when "10000000010101001" => rgb <= "000000";
					when "10000000010101010" => rgb <= "000000";
					when "10000000010101011" => rgb <= "000000";
					when "10000000010101100" => rgb <= "000000";
					when "10000000010101101" => rgb <= "000000";
					when "10000000010101110" => rgb <= "000000";
					when "10000000010101111" => rgb <= "000000";
					when "10000000010110000" => rgb <= "000000";
					when "10000000010110001" => rgb <= "000000";
					when "10000000010110010" => rgb <= "000000";
					when "10000000010110011" => rgb <= "000000";
					when "10000000010110100" => rgb <= "000000";
					when "10000000010110101" => rgb <= "000000";
					when "10000000010110110" => rgb <= "000000";
					when "10000000010110111" => rgb <= "000000";
					when "10000000010111000" => rgb <= "000000";
					when "10000000010111001" => rgb <= "000000";
					when "10000000010111010" => rgb <= "000000";
					when "10000000010111011" => rgb <= "000000";
					when "10000000010111100" => rgb <= "000000";
					when "10000000010111101" => rgb <= "000000";
					when "10000000010111110" => rgb <= "000000";
					when "10000000010111111" => rgb <= "000000";
					when "10000000011000000" => rgb <= "000000";
					when "10000000011000001" => rgb <= "000000";
					when "10000000011000010" => rgb <= "000000";
					when "10000000011000011" => rgb <= "000000";
					when "10000000011000100" => rgb <= "000000";
					when "10000000011000101" => rgb <= "000000";
					when "10000000011000110" => rgb <= "000000";
					when "10000000011000111" => rgb <= "000000";
					when "10000000011001000" => rgb <= "000000";
					when "10000000011001001" => rgb <= "000000";
					when "10000000011001010" => rgb <= "000000";
					when "10000000011001011" => rgb <= "000000";
					when "10000000011001100" => rgb <= "000000";
					when "10000000011001101" => rgb <= "000000";
					when "10000000011001110" => rgb <= "000000";
					when "10000000011001111" => rgb <= "000000";
					when "10000000011010000" => rgb <= "000000";
					when "10000000011010001" => rgb <= "000000";
					when "10000000011010010" => rgb <= "000000";
					when "10000000011010011" => rgb <= "000000";
					when "10000000011010100" => rgb <= "000000";
					when "10000000011010101" => rgb <= "000000";
					when "10000000011010110" => rgb <= "000000";
					when "10000000011010111" => rgb <= "000000";
					when "10000000011011000" => rgb <= "000000";
					when "10000000011011001" => rgb <= "000000";
					when "10000000011011010" => rgb <= "000000";
					when "10000000011011011" => rgb <= "000000";
					when "10000000011011100" => rgb <= "000000";
					when "10000000011011101" => rgb <= "000000";
					when "10000000011011110" => rgb <= "000000";
					when "10000000011011111" => rgb <= "000000";
					when "10000000011100000" => rgb <= "000000";
					when "10000000011100001" => rgb <= "000000";
					when "10000000011100010" => rgb <= "000000";
					when "10000000011100011" => rgb <= "000000";
					when "10000000011100100" => rgb <= "000000";
					when "10000000011100101" => rgb <= "000000";
					when "10000000011100110" => rgb <= "000000";
					when "10000000011100111" => rgb <= "000000";
					when "10000000011101000" => rgb <= "000000";
					when "10000000011101001" => rgb <= "000000";
					when "10000000011101010" => rgb <= "000000";
					when "10000000011101011" => rgb <= "000000";
					when "10000000011101100" => rgb <= "000000";
					when "10000000011101101" => rgb <= "000000";
					when "10000000011101110" => rgb <= "000000";
					when "10000000011101111" => rgb <= "000000";
					when "10000000011110000" => rgb <= "000000";
					when "10000000011110001" => rgb <= "000000";
					when "10000000011110010" => rgb <= "000000";
					when "10000000011110011" => rgb <= "000000";
					when "10000000011110100" => rgb <= "000000";
					when "10000000011110101" => rgb <= "000000";
					when "10000000011110110" => rgb <= "000000";
					when "10000000011110111" => rgb <= "000000";
					when "10000000011111000" => rgb <= "000000";
					when "10000000011111001" => rgb <= "000000";
					when "10000000011111010" => rgb <= "000000";
					when "10000000011111011" => rgb <= "000000";
					when "10000000011111100" => rgb <= "000000";
					when "10000000011111101" => rgb <= "000000";
					when "10000000011111110" => rgb <= "000000";
					when "10000000011111111" => rgb <= "000000";
					when "10000000100000000" => rgb <= "000000";
					when "10000000100000001" => rgb <= "000000";
					when "10000000100000010" => rgb <= "000000";
					when "10000000100000011" => rgb <= "000000";
					when "10000000100000100" => rgb <= "000000";
					when "10000000100000101" => rgb <= "000000";
					when "10000000100000110" => rgb <= "000000";
					when "10000000100000111" => rgb <= "000000";
					when "10000000100001000" => rgb <= "000000";
					when "10000000100001001" => rgb <= "000000";
					when "10000000100001010" => rgb <= "000000";
					when "10000000100001011" => rgb <= "000000";
					when "10000000100001100" => rgb <= "000000";
					when "10000000100001101" => rgb <= "000000";
					when "10000000100001110" => rgb <= "000000";
					when "10000000100001111" => rgb <= "000000";
					when "10000000100010000" => rgb <= "000000";
					when "10000000100010001" => rgb <= "000000";
					when "10000000100010010" => rgb <= "000000";
					when "10000000100010011" => rgb <= "000000";
					when "10000000100010100" => rgb <= "000000";
					when "10000000100010101" => rgb <= "000000";
					when "10000000100010110" => rgb <= "000000";
					when "10000000100010111" => rgb <= "000000";
					when "10000000100011000" => rgb <= "000000";
					when "10000000100011001" => rgb <= "000000";
					when "10000000100011010" => rgb <= "000000";
					when "10000000100011011" => rgb <= "000000";
					when "10000000100011100" => rgb <= "000000";
					when "10000000100011101" => rgb <= "000000";
					when "10000000100011110" => rgb <= "000000";
					when "10000000100011111" => rgb <= "000000";
					when "10000000100100000" => rgb <= "000000";
					when "10000000100100001" => rgb <= "000000";
					when "10000000100100010" => rgb <= "000000";
					when "10000000100100011" => rgb <= "000000";
					when "10000000100100100" => rgb <= "000000";
					when "10000000100100101" => rgb <= "000000";
					when "10000000100100110" => rgb <= "000000";
					when "10000000100100111" => rgb <= "000000";
					when "10000000100101000" => rgb <= "000000";
					when "10000000100101001" => rgb <= "000000";
					when "10000000100101010" => rgb <= "000000";
					when "10000000100101011" => rgb <= "000000";
					when "10000000100101100" => rgb <= "000000";
					when "10000000100101101" => rgb <= "000000";
					when "10000000100101110" => rgb <= "000000";
					when "10000000100101111" => rgb <= "000000";
					when "10000000100110000" => rgb <= "000000";
					when "10000000100110001" => rgb <= "000000";
					when "10000000100110010" => rgb <= "000000";
					when "10000000100110011" => rgb <= "000000";
					when "10000000100110100" => rgb <= "000000";
					when "10000000100110101" => rgb <= "000000";
					when "10000000100110110" => rgb <= "000000";
					when "10000000100110111" => rgb <= "000000";
					when "10000000100111000" => rgb <= "000000";
					when "10000000100111001" => rgb <= "000000";
					when "10000000100111010" => rgb <= "000000";
					when "10000000100111011" => rgb <= "000000";
					when "10000000100111100" => rgb <= "000000";
					when "10000000100111101" => rgb <= "000000";
					when "10000000100111110" => rgb <= "000000";
					when "10000000100111111" => rgb <= "000000";
					when "10000001000000000" => rgb <= "000000";
					when "10000001000000001" => rgb <= "000000";
					when "10000001000000010" => rgb <= "000000";
					when "10000001000000011" => rgb <= "000000";
					when "10000001000000100" => rgb <= "000000";
					when "10000001000000101" => rgb <= "000000";
					when "10000001000000110" => rgb <= "000000";
					when "10000001000000111" => rgb <= "000000";
					when "10000001000001000" => rgb <= "000000";
					when "10000001000001001" => rgb <= "000000";
					when "10000001000001010" => rgb <= "000000";
					when "10000001000001011" => rgb <= "000000";
					when "10000001000001100" => rgb <= "000000";
					when "10000001000001101" => rgb <= "000000";
					when "10000001000001110" => rgb <= "000000";
					when "10000001000001111" => rgb <= "000000";
					when "10000001000010000" => rgb <= "000000";
					when "10000001000010001" => rgb <= "000000";
					when "10000001000010010" => rgb <= "000000";
					when "10000001000010011" => rgb <= "000000";
					when "10000001000010100" => rgb <= "000000";
					when "10000001000010101" => rgb <= "000000";
					when "10000001000010110" => rgb <= "000000";
					when "10000001000010111" => rgb <= "000000";
					when "10000001000011000" => rgb <= "000000";
					when "10000001000011001" => rgb <= "000000";
					when "10000001000011010" => rgb <= "000000";
					when "10000001000011011" => rgb <= "000000";
					when "10000001000011100" => rgb <= "000000";
					when "10000001000011101" => rgb <= "000000";
					when "10000001000011110" => rgb <= "000000";
					when "10000001000011111" => rgb <= "000000";
					when "10000001000100000" => rgb <= "000000";
					when "10000001000100001" => rgb <= "000000";
					when "10000001000100010" => rgb <= "000000";
					when "10000001000100011" => rgb <= "000000";
					when "10000001000100100" => rgb <= "000000";
					when "10000001000100101" => rgb <= "000000";
					when "10000001000100110" => rgb <= "000000";
					when "10000001000100111" => rgb <= "000000";
					when "10000001000101000" => rgb <= "000000";
					when "10000001000101001" => rgb <= "000000";
					when "10000001000101010" => rgb <= "000000";
					when "10000001000101011" => rgb <= "000000";
					when "10000001000101100" => rgb <= "000000";
					when "10000001000101101" => rgb <= "000000";
					when "10000001000101110" => rgb <= "000000";
					when "10000001000101111" => rgb <= "000000";
					when "10000001000110000" => rgb <= "000000";
					when "10000001000110001" => rgb <= "000000";
					when "10000001000110010" => rgb <= "000000";
					when "10000001000110011" => rgb <= "000000";
					when "10000001000110100" => rgb <= "000000";
					when "10000001000110101" => rgb <= "000000";
					when "10000001000110110" => rgb <= "000000";
					when "10000001000110111" => rgb <= "000000";
					when "10000001000111000" => rgb <= "000000";
					when "10000001000111001" => rgb <= "000000";
					when "10000001000111010" => rgb <= "000000";
					when "10000001000111011" => rgb <= "000000";
					when "10000001000111100" => rgb <= "000000";
					when "10000001000111101" => rgb <= "000000";
					when "10000001000111110" => rgb <= "000000";
					when "10000001000111111" => rgb <= "000000";
					when "10000001001000000" => rgb <= "000000";
					when "10000001001000001" => rgb <= "000000";
					when "10000001001000010" => rgb <= "000000";
					when "10000001001000011" => rgb <= "000000";
					when "10000001001000100" => rgb <= "000000";
					when "10000001001000101" => rgb <= "000000";
					when "10000001001000110" => rgb <= "000000";
					when "10000001001000111" => rgb <= "000000";
					when "10000001001001000" => rgb <= "000000";
					when "10000001001001001" => rgb <= "000000";
					when "10000001001001010" => rgb <= "000000";
					when "10000001001001011" => rgb <= "000000";
					when "10000001001001100" => rgb <= "000000";
					when "10000001001001101" => rgb <= "000000";
					when "10000001001001110" => rgb <= "000000";
					when "10000001001001111" => rgb <= "000000";
					when "10000001001010000" => rgb <= "000000";
					when "10000001001010001" => rgb <= "000000";
					when "10000001001010010" => rgb <= "000000";
					when "10000001001010011" => rgb <= "000000";
					when "10000001001010100" => rgb <= "000000";
					when "10000001001010101" => rgb <= "000000";
					when "10000001001010110" => rgb <= "000000";
					when "10000001001010111" => rgb <= "000000";
					when "10000001001011000" => rgb <= "000000";
					when "10000001001011001" => rgb <= "000000";
					when "10000001001011010" => rgb <= "000000";
					when "10000001001011011" => rgb <= "000000";
					when "10000001001011100" => rgb <= "000000";
					when "10000001001011101" => rgb <= "000000";
					when "10000001001011110" => rgb <= "000000";
					when "10000001001011111" => rgb <= "000000";
					when "10000001001100000" => rgb <= "000000";
					when "10000001001100001" => rgb <= "000000";
					when "10000001001100010" => rgb <= "000000";
					when "10000001001100011" => rgb <= "000000";
					when "10000001001100100" => rgb <= "000000";
					when "10000001001100101" => rgb <= "000000";
					when "10000001001100110" => rgb <= "000000";
					when "10000001001100111" => rgb <= "000000";
					when "10000001001101000" => rgb <= "000000";
					when "10000001001101001" => rgb <= "000000";
					when "10000001001101010" => rgb <= "000000";
					when "10000001001101011" => rgb <= "000000";
					when "10000001001101100" => rgb <= "000000";
					when "10000001001101101" => rgb <= "000000";
					when "10000001001101110" => rgb <= "000000";
					when "10000001001101111" => rgb <= "000000";
					when "10000001001110000" => rgb <= "000000";
					when "10000001001110001" => rgb <= "000000";
					when "10000001001110010" => rgb <= "000000";
					when "10000001001110011" => rgb <= "000000";
					when "10000001001110100" => rgb <= "000000";
					when "10000001001110101" => rgb <= "000000";
					when "10000001001110110" => rgb <= "000000";
					when "10000001001110111" => rgb <= "000000";
					when "10000001001111000" => rgb <= "000000";
					when "10000001001111001" => rgb <= "000000";
					when "10000001001111010" => rgb <= "000000";
					when "10000001001111011" => rgb <= "000000";
					when "10000001001111100" => rgb <= "000000";
					when "10000001001111101" => rgb <= "000000";
					when "10000001001111110" => rgb <= "000000";
					when "10000001001111111" => rgb <= "000000";
					when "10000001010000000" => rgb <= "000000";
					when "10000001010000001" => rgb <= "000000";
					when "10000001010000010" => rgb <= "000000";
					when "10000001010000011" => rgb <= "000000";
					when "10000001010000100" => rgb <= "000000";
					when "10000001010000101" => rgb <= "000000";
					when "10000001010000110" => rgb <= "000000";
					when "10000001010000111" => rgb <= "000000";
					when "10000001010001000" => rgb <= "000000";
					when "10000001010001001" => rgb <= "000000";
					when "10000001010001010" => rgb <= "000000";
					when "10000001010001011" => rgb <= "000000";
					when "10000001010001100" => rgb <= "000000";
					when "10000001010001101" => rgb <= "000000";
					when "10000001010001110" => rgb <= "000000";
					when "10000001010001111" => rgb <= "000000";
					when "10000001010010000" => rgb <= "000000";
					when "10000001010010001" => rgb <= "000000";
					when "10000001010010010" => rgb <= "000000";
					when "10000001010010011" => rgb <= "000000";
					when "10000001010010100" => rgb <= "000000";
					when "10000001010010101" => rgb <= "000000";
					when "10000001010010110" => rgb <= "000000";
					when "10000001010010111" => rgb <= "000000";
					when "10000001010011000" => rgb <= "000000";
					when "10000001010011001" => rgb <= "000000";
					when "10000001010011010" => rgb <= "000000";
					when "10000001010011011" => rgb <= "000000";
					when "10000001010011100" => rgb <= "000000";
					when "10000001010011101" => rgb <= "000000";
					when "10000001010011110" => rgb <= "000000";
					when "10000001010011111" => rgb <= "000000";
					when "10000001010100000" => rgb <= "000000";
					when "10000001010100001" => rgb <= "000000";
					when "10000001010100010" => rgb <= "000000";
					when "10000001010100011" => rgb <= "000000";
					when "10000001010100100" => rgb <= "000000";
					when "10000001010100101" => rgb <= "000000";
					when "10000001010100110" => rgb <= "000000";
					when "10000001010100111" => rgb <= "000000";
					when "10000001010101000" => rgb <= "000000";
					when "10000001010101001" => rgb <= "000000";
					when "10000001010101010" => rgb <= "000000";
					when "10000001010101011" => rgb <= "000000";
					when "10000001010101100" => rgb <= "000000";
					when "10000001010101101" => rgb <= "000000";
					when "10000001010101110" => rgb <= "000000";
					when "10000001010101111" => rgb <= "000000";
					when "10000001010110000" => rgb <= "000000";
					when "10000001010110001" => rgb <= "000000";
					when "10000001010110010" => rgb <= "000000";
					when "10000001010110011" => rgb <= "000000";
					when "10000001010110100" => rgb <= "000000";
					when "10000001010110101" => rgb <= "000000";
					when "10000001010110110" => rgb <= "000000";
					when "10000001010110111" => rgb <= "000000";
					when "10000001010111000" => rgb <= "000000";
					when "10000001010111001" => rgb <= "000000";
					when "10000001010111010" => rgb <= "000000";
					when "10000001010111011" => rgb <= "000000";
					when "10000001010111100" => rgb <= "000000";
					when "10000001010111101" => rgb <= "000000";
					when "10000001010111110" => rgb <= "000000";
					when "10000001010111111" => rgb <= "000000";
					when "10000001011000000" => rgb <= "000000";
					when "10000001011000001" => rgb <= "000000";
					when "10000001011000010" => rgb <= "000000";
					when "10000001011000011" => rgb <= "000000";
					when "10000001011000100" => rgb <= "000000";
					when "10000001011000101" => rgb <= "000000";
					when "10000001011000110" => rgb <= "000000";
					when "10000001011000111" => rgb <= "000000";
					when "10000001011001000" => rgb <= "000000";
					when "10000001011001001" => rgb <= "000000";
					when "10000001011001010" => rgb <= "000000";
					when "10000001011001011" => rgb <= "000000";
					when "10000001011001100" => rgb <= "000000";
					when "10000001011001101" => rgb <= "000000";
					when "10000001011001110" => rgb <= "000000";
					when "10000001011001111" => rgb <= "000000";
					when "10000001011010000" => rgb <= "000000";
					when "10000001011010001" => rgb <= "000000";
					when "10000001011010010" => rgb <= "000000";
					when "10000001011010011" => rgb <= "000000";
					when "10000001011010100" => rgb <= "000000";
					when "10000001011010101" => rgb <= "000000";
					when "10000001011010110" => rgb <= "000000";
					when "10000001011010111" => rgb <= "000000";
					when "10000001011011000" => rgb <= "000000";
					when "10000001011011001" => rgb <= "000000";
					when "10000001011011010" => rgb <= "000000";
					when "10000001011011011" => rgb <= "000000";
					when "10000001011011100" => rgb <= "000000";
					when "10000001011011101" => rgb <= "000000";
					when "10000001011011110" => rgb <= "000000";
					when "10000001011011111" => rgb <= "000000";
					when "10000001011100000" => rgb <= "000000";
					when "10000001011100001" => rgb <= "000000";
					when "10000001011100010" => rgb <= "000000";
					when "10000001011100011" => rgb <= "000000";
					when "10000001011100100" => rgb <= "000000";
					when "10000001011100101" => rgb <= "000000";
					when "10000001011100110" => rgb <= "000000";
					when "10000001011100111" => rgb <= "000000";
					when "10000001011101000" => rgb <= "000000";
					when "10000001011101001" => rgb <= "000000";
					when "10000001011101010" => rgb <= "000000";
					when "10000001011101011" => rgb <= "000000";
					when "10000001011101100" => rgb <= "000000";
					when "10000001011101101" => rgb <= "000000";
					when "10000001011101110" => rgb <= "000000";
					when "10000001011101111" => rgb <= "000000";
					when "10000001011110000" => rgb <= "000000";
					when "10000001011110001" => rgb <= "000000";
					when "10000001011110010" => rgb <= "000000";
					when "10000001011110011" => rgb <= "000000";
					when "10000001011110100" => rgb <= "000000";
					when "10000001011110101" => rgb <= "000000";
					when "10000001011110110" => rgb <= "000000";
					when "10000001011110111" => rgb <= "000000";
					when "10000001011111000" => rgb <= "000000";
					when "10000001011111001" => rgb <= "000000";
					when "10000001011111010" => rgb <= "000000";
					when "10000001011111011" => rgb <= "000000";
					when "10000001011111100" => rgb <= "000000";
					when "10000001011111101" => rgb <= "000000";
					when "10000001011111110" => rgb <= "000000";
					when "10000001011111111" => rgb <= "000000";
					when "10000001100000000" => rgb <= "000000";
					when "10000001100000001" => rgb <= "000000";
					when "10000001100000010" => rgb <= "000000";
					when "10000001100000011" => rgb <= "000000";
					when "10000001100000100" => rgb <= "000000";
					when "10000001100000101" => rgb <= "000000";
					when "10000001100000110" => rgb <= "000000";
					when "10000001100000111" => rgb <= "000000";
					when "10000001100001000" => rgb <= "000000";
					when "10000001100001001" => rgb <= "000000";
					when "10000001100001010" => rgb <= "000000";
					when "10000001100001011" => rgb <= "000000";
					when "10000001100001100" => rgb <= "000000";
					when "10000001100001101" => rgb <= "000000";
					when "10000001100001110" => rgb <= "000000";
					when "10000001100001111" => rgb <= "000000";
					when "10000001100010000" => rgb <= "000000";
					when "10000001100010001" => rgb <= "000000";
					when "10000001100010010" => rgb <= "000000";
					when "10000001100010011" => rgb <= "000000";
					when "10000001100010100" => rgb <= "000000";
					when "10000001100010101" => rgb <= "000000";
					when "10000001100010110" => rgb <= "000000";
					when "10000001100010111" => rgb <= "000000";
					when "10000001100011000" => rgb <= "000000";
					when "10000001100011001" => rgb <= "000000";
					when "10000001100011010" => rgb <= "000000";
					when "10000001100011011" => rgb <= "000000";
					when "10000001100011100" => rgb <= "000000";
					when "10000001100011101" => rgb <= "000000";
					when "10000001100011110" => rgb <= "000000";
					when "10000001100011111" => rgb <= "000000";
					when "10000001100100000" => rgb <= "000000";
					when "10000001100100001" => rgb <= "000000";
					when "10000001100100010" => rgb <= "000000";
					when "10000001100100011" => rgb <= "000000";
					when "10000001100100100" => rgb <= "000000";
					when "10000001100100101" => rgb <= "000000";
					when "10000001100100110" => rgb <= "000000";
					when "10000001100100111" => rgb <= "000000";
					when "10000001100101000" => rgb <= "000000";
					when "10000001100101001" => rgb <= "000000";
					when "10000001100101010" => rgb <= "000000";
					when "10000001100101011" => rgb <= "000000";
					when "10000001100101100" => rgb <= "000000";
					when "10000001100101101" => rgb <= "000000";
					when "10000001100101110" => rgb <= "000000";
					when "10000001100101111" => rgb <= "000000";
					when "10000001100110000" => rgb <= "000000";
					when "10000001100110001" => rgb <= "000000";
					when "10000001100110010" => rgb <= "000000";
					when "10000001100110011" => rgb <= "000000";
					when "10000001100110100" => rgb <= "000000";
					when "10000001100110101" => rgb <= "000000";
					when "10000001100110110" => rgb <= "000000";
					when "10000001100110111" => rgb <= "000000";
					when "10000001100111000" => rgb <= "000000";
					when "10000001100111001" => rgb <= "000000";
					when "10000001100111010" => rgb <= "000000";
					when "10000001100111011" => rgb <= "000000";
					when "10000001100111100" => rgb <= "000000";
					when "10000001100111101" => rgb <= "000000";
					when "10000001100111110" => rgb <= "000000";
					when "10000001100111111" => rgb <= "000000";
					when "10000010000000000" => rgb <= "000000";
					when "10000010000000001" => rgb <= "000000";
					when "10000010000000010" => rgb <= "000000";
					when "10000010000000011" => rgb <= "000000";
					when "10000010000000100" => rgb <= "000000";
					when "10000010000000101" => rgb <= "000000";
					when "10000010000000110" => rgb <= "000000";
					when "10000010000000111" => rgb <= "000000";
					when "10000010000001000" => rgb <= "000000";
					when "10000010000001001" => rgb <= "000000";
					when "10000010000001010" => rgb <= "000000";
					when "10000010000001011" => rgb <= "000000";
					when "10000010000001100" => rgb <= "000000";
					when "10000010000001101" => rgb <= "000000";
					when "10000010000001110" => rgb <= "000000";
					when "10000010000001111" => rgb <= "000000";
					when "10000010000010000" => rgb <= "000000";
					when "10000010000010001" => rgb <= "000000";
					when "10000010000010010" => rgb <= "000000";
					when "10000010000010011" => rgb <= "000000";
					when "10000010000010100" => rgb <= "000000";
					when "10000010000010101" => rgb <= "000000";
					when "10000010000010110" => rgb <= "000000";
					when "10000010000010111" => rgb <= "000000";
					when "10000010000011000" => rgb <= "000000";
					when "10000010000011001" => rgb <= "000000";
					when "10000010000011010" => rgb <= "000000";
					when "10000010000011011" => rgb <= "000000";
					when "10000010000011100" => rgb <= "000000";
					when "10000010000011101" => rgb <= "000000";
					when "10000010000011110" => rgb <= "000000";
					when "10000010000011111" => rgb <= "000000";
					when "10000010000100000" => rgb <= "000000";
					when "10000010000100001" => rgb <= "000000";
					when "10000010000100010" => rgb <= "000000";
					when "10000010000100011" => rgb <= "000000";
					when "10000010000100100" => rgb <= "000000";
					when "10000010000100101" => rgb <= "000000";
					when "10000010000100110" => rgb <= "000000";
					when "10000010000100111" => rgb <= "000000";
					when "10000010000101000" => rgb <= "000000";
					when "10000010000101001" => rgb <= "000000";
					when "10000010000101010" => rgb <= "000000";
					when "10000010000101011" => rgb <= "000000";
					when "10000010000101100" => rgb <= "000000";
					when "10000010000101101" => rgb <= "000000";
					when "10000010000101110" => rgb <= "000000";
					when "10000010000101111" => rgb <= "000000";
					when "10000010000110000" => rgb <= "000000";
					when "10000010000110001" => rgb <= "000000";
					when "10000010000110010" => rgb <= "000000";
					when "10000010000110011" => rgb <= "000000";
					when "10000010000110100" => rgb <= "000000";
					when "10000010000110101" => rgb <= "000000";
					when "10000010000110110" => rgb <= "000000";
					when "10000010000110111" => rgb <= "000000";
					when "10000010000111000" => rgb <= "000000";
					when "10000010000111001" => rgb <= "000000";
					when "10000010000111010" => rgb <= "000000";
					when "10000010000111011" => rgb <= "000000";
					when "10000010000111100" => rgb <= "000000";
					when "10000010000111101" => rgb <= "000000";
					when "10000010000111110" => rgb <= "000000";
					when "10000010000111111" => rgb <= "000000";
					when "10000010001000000" => rgb <= "000000";
					when "10000010001000001" => rgb <= "000000";
					when "10000010001000010" => rgb <= "000000";
					when "10000010001000011" => rgb <= "000000";
					when "10000010001000100" => rgb <= "000000";
					when "10000010001000101" => rgb <= "000000";
					when "10000010001000110" => rgb <= "000000";
					when "10000010001000111" => rgb <= "000000";
					when "10000010001001000" => rgb <= "000000";
					when "10000010001001001" => rgb <= "000000";
					when "10000010001001010" => rgb <= "000000";
					when "10000010001001011" => rgb <= "000000";
					when "10000010001001100" => rgb <= "000000";
					when "10000010001001101" => rgb <= "000000";
					when "10000010001001110" => rgb <= "000000";
					when "10000010001001111" => rgb <= "000000";
					when "10000010001010000" => rgb <= "000000";
					when "10000010001010001" => rgb <= "000000";
					when "10000010001010010" => rgb <= "000000";
					when "10000010001010011" => rgb <= "000000";
					when "10000010001010100" => rgb <= "000000";
					when "10000010001010101" => rgb <= "000000";
					when "10000010001010110" => rgb <= "000000";
					when "10000010001010111" => rgb <= "000000";
					when "10000010001011000" => rgb <= "000000";
					when "10000010001011001" => rgb <= "000000";
					when "10000010001011010" => rgb <= "000000";
					when "10000010001011011" => rgb <= "000000";
					when "10000010001011100" => rgb <= "000000";
					when "10000010001011101" => rgb <= "000000";
					when "10000010001011110" => rgb <= "000000";
					when "10000010001011111" => rgb <= "000000";
					when "10000010001100000" => rgb <= "000000";
					when "10000010001100001" => rgb <= "000000";
					when "10000010001100010" => rgb <= "000000";
					when "10000010001100011" => rgb <= "000000";
					when "10000010001100100" => rgb <= "000000";
					when "10000010001100101" => rgb <= "000000";
					when "10000010001100110" => rgb <= "000000";
					when "10000010001100111" => rgb <= "000000";
					when "10000010001101000" => rgb <= "000000";
					when "10000010001101001" => rgb <= "000000";
					when "10000010001101010" => rgb <= "000000";
					when "10000010001101011" => rgb <= "000000";
					when "10000010001101100" => rgb <= "000000";
					when "10000010001101101" => rgb <= "000000";
					when "10000010001101110" => rgb <= "000000";
					when "10000010001101111" => rgb <= "000000";
					when "10000010001110000" => rgb <= "000000";
					when "10000010001110001" => rgb <= "000000";
					when "10000010001110010" => rgb <= "000000";
					when "10000010001110011" => rgb <= "000000";
					when "10000010001110100" => rgb <= "000000";
					when "10000010001110101" => rgb <= "000000";
					when "10000010001110110" => rgb <= "000000";
					when "10000010001110111" => rgb <= "000000";
					when "10000010001111000" => rgb <= "000000";
					when "10000010001111001" => rgb <= "000000";
					when "10000010001111010" => rgb <= "000000";
					when "10000010001111011" => rgb <= "000000";
					when "10000010001111100" => rgb <= "000000";
					when "10000010001111101" => rgb <= "000000";
					when "10000010001111110" => rgb <= "000000";
					when "10000010001111111" => rgb <= "000000";
					when "10000010010000000" => rgb <= "000000";
					when "10000010010000001" => rgb <= "000000";
					when "10000010010000010" => rgb <= "000000";
					when "10000010010000011" => rgb <= "000000";
					when "10000010010000100" => rgb <= "000000";
					when "10000010010000101" => rgb <= "000000";
					when "10000010010000110" => rgb <= "000000";
					when "10000010010000111" => rgb <= "000000";
					when "10000010010001000" => rgb <= "000000";
					when "10000010010001001" => rgb <= "000000";
					when "10000010010001010" => rgb <= "000000";
					when "10000010010001011" => rgb <= "000000";
					when "10000010010001100" => rgb <= "000000";
					when "10000010010001101" => rgb <= "000000";
					when "10000010010001110" => rgb <= "000000";
					when "10000010010001111" => rgb <= "000000";
					when "10000010010010000" => rgb <= "000000";
					when "10000010010010001" => rgb <= "000000";
					when "10000010010010010" => rgb <= "000000";
					when "10000010010010011" => rgb <= "000000";
					when "10000010010010100" => rgb <= "000000";
					when "10000010010010101" => rgb <= "000000";
					when "10000010010010110" => rgb <= "000000";
					when "10000010010010111" => rgb <= "000000";
					when "10000010010011000" => rgb <= "000000";
					when "10000010010011001" => rgb <= "000000";
					when "10000010010011010" => rgb <= "000000";
					when "10000010010011011" => rgb <= "000000";
					when "10000010010011100" => rgb <= "000000";
					when "10000010010011101" => rgb <= "000000";
					when "10000010010011110" => rgb <= "000000";
					when "10000010010011111" => rgb <= "000000";
					when "10000010010100000" => rgb <= "000000";
					when "10000010010100001" => rgb <= "000000";
					when "10000010010100010" => rgb <= "000000";
					when "10000010010100011" => rgb <= "000000";
					when "10000010010100100" => rgb <= "000000";
					when "10000010010100101" => rgb <= "000000";
					when "10000010010100110" => rgb <= "000000";
					when "10000010010100111" => rgb <= "000000";
					when "10000010010101000" => rgb <= "000000";
					when "10000010010101001" => rgb <= "000000";
					when "10000010010101010" => rgb <= "000000";
					when "10000010010101011" => rgb <= "000000";
					when "10000010010101100" => rgb <= "000000";
					when "10000010010101101" => rgb <= "000000";
					when "10000010010101110" => rgb <= "000000";
					when "10000010010101111" => rgb <= "000000";
					when "10000010010110000" => rgb <= "000000";
					when "10000010010110001" => rgb <= "000000";
					when "10000010010110010" => rgb <= "000000";
					when "10000010010110011" => rgb <= "000000";
					when "10000010010110100" => rgb <= "000000";
					when "10000010010110101" => rgb <= "000000";
					when "10000010010110110" => rgb <= "000000";
					when "10000010010110111" => rgb <= "000000";
					when "10000010010111000" => rgb <= "000000";
					when "10000010010111001" => rgb <= "000000";
					when "10000010010111010" => rgb <= "000000";
					when "10000010010111011" => rgb <= "000000";
					when "10000010010111100" => rgb <= "000000";
					when "10000010010111101" => rgb <= "000000";
					when "10000010010111110" => rgb <= "000000";
					when "10000010010111111" => rgb <= "000000";
					when "10000010011000000" => rgb <= "000000";
					when "10000010011000001" => rgb <= "000000";
					when "10000010011000010" => rgb <= "000000";
					when "10000010011000011" => rgb <= "000000";
					when "10000010011000100" => rgb <= "000000";
					when "10000010011000101" => rgb <= "000000";
					when "10000010011000110" => rgb <= "000000";
					when "10000010011000111" => rgb <= "000000";
					when "10000010011001000" => rgb <= "000000";
					when "10000010011001001" => rgb <= "000000";
					when "10000010011001010" => rgb <= "000000";
					when "10000010011001011" => rgb <= "000000";
					when "10000010011001100" => rgb <= "000000";
					when "10000010011001101" => rgb <= "000000";
					when "10000010011001110" => rgb <= "000000";
					when "10000010011001111" => rgb <= "000000";
					when "10000010011010000" => rgb <= "000000";
					when "10000010011010001" => rgb <= "000000";
					when "10000010011010010" => rgb <= "000000";
					when "10000010011010011" => rgb <= "000000";
					when "10000010011010100" => rgb <= "000000";
					when "10000010011010101" => rgb <= "000000";
					when "10000010011010110" => rgb <= "000000";
					when "10000010011010111" => rgb <= "000000";
					when "10000010011011000" => rgb <= "000000";
					when "10000010011011001" => rgb <= "000000";
					when "10000010011011010" => rgb <= "000000";
					when "10000010011011011" => rgb <= "000000";
					when "10000010011011100" => rgb <= "000000";
					when "10000010011011101" => rgb <= "000000";
					when "10000010011011110" => rgb <= "000000";
					when "10000010011011111" => rgb <= "000000";
					when "10000010011100000" => rgb <= "000000";
					when "10000010011100001" => rgb <= "000000";
					when "10000010011100010" => rgb <= "000000";
					when "10000010011100011" => rgb <= "000000";
					when "10000010011100100" => rgb <= "000000";
					when "10000010011100101" => rgb <= "000000";
					when "10000010011100110" => rgb <= "000000";
					when "10000010011100111" => rgb <= "000000";
					when "10000010011101000" => rgb <= "000000";
					when "10000010011101001" => rgb <= "000000";
					when "10000010011101010" => rgb <= "000000";
					when "10000010011101011" => rgb <= "000000";
					when "10000010011101100" => rgb <= "000000";
					when "10000010011101101" => rgb <= "000000";
					when "10000010011101110" => rgb <= "000000";
					when "10000010011101111" => rgb <= "000000";
					when "10000010011110000" => rgb <= "000000";
					when "10000010011110001" => rgb <= "000000";
					when "10000010011110010" => rgb <= "000000";
					when "10000010011110011" => rgb <= "000000";
					when "10000010011110100" => rgb <= "000000";
					when "10000010011110101" => rgb <= "000000";
					when "10000010011110110" => rgb <= "000000";
					when "10000010011110111" => rgb <= "000000";
					when "10000010011111000" => rgb <= "000000";
					when "10000010011111001" => rgb <= "000000";
					when "10000010011111010" => rgb <= "000000";
					when "10000010011111011" => rgb <= "000000";
					when "10000010011111100" => rgb <= "000000";
					when "10000010011111101" => rgb <= "000000";
					when "10000010011111110" => rgb <= "000000";
					when "10000010011111111" => rgb <= "000000";
					when "10000010100000000" => rgb <= "000000";
					when "10000010100000001" => rgb <= "000000";
					when "10000010100000010" => rgb <= "000000";
					when "10000010100000011" => rgb <= "000000";
					when "10000010100000100" => rgb <= "000000";
					when "10000010100000101" => rgb <= "000000";
					when "10000010100000110" => rgb <= "000000";
					when "10000010100000111" => rgb <= "000000";
					when "10000010100001000" => rgb <= "000000";
					when "10000010100001001" => rgb <= "000000";
					when "10000010100001010" => rgb <= "000000";
					when "10000010100001011" => rgb <= "000000";
					when "10000010100001100" => rgb <= "000000";
					when "10000010100001101" => rgb <= "000000";
					when "10000010100001110" => rgb <= "000000";
					when "10000010100001111" => rgb <= "000000";
					when "10000010100010000" => rgb <= "000000";
					when "10000010100010001" => rgb <= "000000";
					when "10000010100010010" => rgb <= "000000";
					when "10000010100010011" => rgb <= "000000";
					when "10000010100010100" => rgb <= "000000";
					when "10000010100010101" => rgb <= "000000";
					when "10000010100010110" => rgb <= "000000";
					when "10000010100010111" => rgb <= "000000";
					when "10000010100011000" => rgb <= "000000";
					when "10000010100011001" => rgb <= "000000";
					when "10000010100011010" => rgb <= "000000";
					when "10000010100011011" => rgb <= "000000";
					when "10000010100011100" => rgb <= "000000";
					when "10000010100011101" => rgb <= "000000";
					when "10000010100011110" => rgb <= "000000";
					when "10000010100011111" => rgb <= "000000";
					when "10000010100100000" => rgb <= "000000";
					when "10000010100100001" => rgb <= "000000";
					when "10000010100100010" => rgb <= "000000";
					when "10000010100100011" => rgb <= "000000";
					when "10000010100100100" => rgb <= "000000";
					when "10000010100100101" => rgb <= "000000";
					when "10000010100100110" => rgb <= "000000";
					when "10000010100100111" => rgb <= "000000";
					when "10000010100101000" => rgb <= "000000";
					when "10000010100101001" => rgb <= "000000";
					when "10000010100101010" => rgb <= "000000";
					when "10000010100101011" => rgb <= "000000";
					when "10000010100101100" => rgb <= "000000";
					when "10000010100101101" => rgb <= "000000";
					when "10000010100101110" => rgb <= "000000";
					when "10000010100101111" => rgb <= "000000";
					when "10000010100110000" => rgb <= "000000";
					when "10000010100110001" => rgb <= "000000";
					when "10000010100110010" => rgb <= "000000";
					when "10000010100110011" => rgb <= "000000";
					when "10000010100110100" => rgb <= "000000";
					when "10000010100110101" => rgb <= "000000";
					when "10000010100110110" => rgb <= "000000";
					when "10000010100110111" => rgb <= "000000";
					when "10000010100111000" => rgb <= "000000";
					when "10000010100111001" => rgb <= "000000";
					when "10000010100111010" => rgb <= "000000";
					when "10000010100111011" => rgb <= "000000";
					when "10000010100111100" => rgb <= "000000";
					when "10000010100111101" => rgb <= "000000";
					when "10000010100111110" => rgb <= "000000";
					when "10000010100111111" => rgb <= "000000";
					when "10000011000000000" => rgb <= "000000";
					when "10000011000000001" => rgb <= "000000";
					when "10000011000000010" => rgb <= "000000";
					when "10000011000000011" => rgb <= "000000";
					when "10000011000000100" => rgb <= "000000";
					when "10000011000000101" => rgb <= "000000";
					when "10000011000000110" => rgb <= "000000";
					when "10000011000000111" => rgb <= "000000";
					when "10000011000001000" => rgb <= "000000";
					when "10000011000001001" => rgb <= "000000";
					when "10000011000001010" => rgb <= "000000";
					when "10000011000001011" => rgb <= "000000";
					when "10000011000001100" => rgb <= "000000";
					when "10000011000001101" => rgb <= "000000";
					when "10000011000001110" => rgb <= "000000";
					when "10000011000001111" => rgb <= "000000";
					when "10000011000010000" => rgb <= "000000";
					when "10000011000010001" => rgb <= "000000";
					when "10000011000010010" => rgb <= "000000";
					when "10000011000010011" => rgb <= "000000";
					when "10000011000010100" => rgb <= "000000";
					when "10000011000010101" => rgb <= "000000";
					when "10000011000010110" => rgb <= "000000";
					when "10000011000010111" => rgb <= "000000";
					when "10000011000011000" => rgb <= "000000";
					when "10000011000011001" => rgb <= "000000";
					when "10000011000011010" => rgb <= "000000";
					when "10000011000011011" => rgb <= "000000";
					when "10000011000011100" => rgb <= "000000";
					when "10000011000011101" => rgb <= "000000";
					when "10000011000011110" => rgb <= "000000";
					when "10000011000011111" => rgb <= "000000";
					when "10000011000100000" => rgb <= "000000";
					when "10000011000100001" => rgb <= "000000";
					when "10000011000100010" => rgb <= "000000";
					when "10000011000100011" => rgb <= "000000";
					when "10000011000100100" => rgb <= "000000";
					when "10000011000100101" => rgb <= "000000";
					when "10000011000100110" => rgb <= "000000";
					when "10000011000100111" => rgb <= "000000";
					when "10000011000101000" => rgb <= "000000";
					when "10000011000101001" => rgb <= "000000";
					when "10000011000101010" => rgb <= "000000";
					when "10000011000101011" => rgb <= "000000";
					when "10000011000101100" => rgb <= "000000";
					when "10000011000101101" => rgb <= "000000";
					when "10000011000101110" => rgb <= "000000";
					when "10000011000101111" => rgb <= "000000";
					when "10000011000110000" => rgb <= "000000";
					when "10000011000110001" => rgb <= "000000";
					when "10000011000110010" => rgb <= "000000";
					when "10000011000110011" => rgb <= "000000";
					when "10000011000110100" => rgb <= "000000";
					when "10000011000110101" => rgb <= "000000";
					when "10000011000110110" => rgb <= "000000";
					when "10000011000110111" => rgb <= "000000";
					when "10000011000111000" => rgb <= "000000";
					when "10000011000111001" => rgb <= "000000";
					when "10000011000111010" => rgb <= "000000";
					when "10000011000111011" => rgb <= "000000";
					when "10000011000111100" => rgb <= "000000";
					when "10000011000111101" => rgb <= "000000";
					when "10000011000111110" => rgb <= "000000";
					when "10000011000111111" => rgb <= "000000";
					when "10000011001000000" => rgb <= "000000";
					when "10000011001000001" => rgb <= "000000";
					when "10000011001000010" => rgb <= "000000";
					when "10000011001000011" => rgb <= "000000";
					when "10000011001000100" => rgb <= "000000";
					when "10000011001000101" => rgb <= "000000";
					when "10000011001000110" => rgb <= "000000";
					when "10000011001000111" => rgb <= "000000";
					when "10000011001001000" => rgb <= "000000";
					when "10000011001001001" => rgb <= "000000";
					when "10000011001001010" => rgb <= "000000";
					when "10000011001001011" => rgb <= "000000";
					when "10000011001001100" => rgb <= "000000";
					when "10000011001001101" => rgb <= "000000";
					when "10000011001001110" => rgb <= "000000";
					when "10000011001001111" => rgb <= "000000";
					when "10000011001010000" => rgb <= "000000";
					when "10000011001010001" => rgb <= "000000";
					when "10000011001010010" => rgb <= "000000";
					when "10000011001010011" => rgb <= "000000";
					when "10000011001010100" => rgb <= "000000";
					when "10000011001010101" => rgb <= "000000";
					when "10000011001010110" => rgb <= "000000";
					when "10000011001010111" => rgb <= "000000";
					when "10000011001011000" => rgb <= "000000";
					when "10000011001011001" => rgb <= "000000";
					when "10000011001011010" => rgb <= "000000";
					when "10000011001011011" => rgb <= "000000";
					when "10000011001011100" => rgb <= "000000";
					when "10000011001011101" => rgb <= "000000";
					when "10000011001011110" => rgb <= "000000";
					when "10000011001011111" => rgb <= "000000";
					when "10000011001100000" => rgb <= "000000";
					when "10000011001100001" => rgb <= "000000";
					when "10000011001100010" => rgb <= "000000";
					when "10000011001100011" => rgb <= "000000";
					when "10000011001100100" => rgb <= "000000";
					when "10000011001100101" => rgb <= "000000";
					when "10000011001100110" => rgb <= "000000";
					when "10000011001100111" => rgb <= "000000";
					when "10000011001101000" => rgb <= "000000";
					when "10000011001101001" => rgb <= "000000";
					when "10000011001101010" => rgb <= "000000";
					when "10000011001101011" => rgb <= "000000";
					when "10000011001101100" => rgb <= "000000";
					when "10000011001101101" => rgb <= "000000";
					when "10000011001101110" => rgb <= "000000";
					when "10000011001101111" => rgb <= "000000";
					when "10000011001110000" => rgb <= "000000";
					when "10000011001110001" => rgb <= "000000";
					when "10000011001110010" => rgb <= "000000";
					when "10000011001110011" => rgb <= "000000";
					when "10000011001110100" => rgb <= "000000";
					when "10000011001110101" => rgb <= "000000";
					when "10000011001110110" => rgb <= "000000";
					when "10000011001110111" => rgb <= "000000";
					when "10000011001111000" => rgb <= "000000";
					when "10000011001111001" => rgb <= "000000";
					when "10000011001111010" => rgb <= "000000";
					when "10000011001111011" => rgb <= "000000";
					when "10000011001111100" => rgb <= "000000";
					when "10000011001111101" => rgb <= "000000";
					when "10000011001111110" => rgb <= "000000";
					when "10000011001111111" => rgb <= "000000";
					when "10000011010000000" => rgb <= "000000";
					when "10000011010000001" => rgb <= "000000";
					when "10000011010000010" => rgb <= "000000";
					when "10000011010000011" => rgb <= "000000";
					when "10000011010000100" => rgb <= "000000";
					when "10000011010000101" => rgb <= "000000";
					when "10000011010000110" => rgb <= "000000";
					when "10000011010000111" => rgb <= "000000";
					when "10000011010001000" => rgb <= "000000";
					when "10000011010001001" => rgb <= "000000";
					when "10000011010001010" => rgb <= "000000";
					when "10000011010001011" => rgb <= "000000";
					when "10000011010001100" => rgb <= "000000";
					when "10000011010001101" => rgb <= "000000";
					when "10000011010001110" => rgb <= "000000";
					when "10000011010001111" => rgb <= "000000";
					when "10000011010010000" => rgb <= "000000";
					when "10000011010010001" => rgb <= "000000";
					when "10000011010010010" => rgb <= "000000";
					when "10000011010010011" => rgb <= "000000";
					when "10000011010010100" => rgb <= "000000";
					when "10000011010010101" => rgb <= "000000";
					when "10000011010010110" => rgb <= "000000";
					when "10000011010010111" => rgb <= "000000";
					when "10000011010011000" => rgb <= "000000";
					when "10000011010011001" => rgb <= "000000";
					when "10000011010011010" => rgb <= "000000";
					when "10000011010011011" => rgb <= "000000";
					when "10000011010011100" => rgb <= "000000";
					when "10000011010011101" => rgb <= "000000";
					when "10000011010011110" => rgb <= "000000";
					when "10000011010011111" => rgb <= "000000";
					when "10000011010100000" => rgb <= "000000";
					when "10000011010100001" => rgb <= "000000";
					when "10000011010100010" => rgb <= "000000";
					when "10000011010100011" => rgb <= "000000";
					when "10000011010100100" => rgb <= "000000";
					when "10000011010100101" => rgb <= "000000";
					when "10000011010100110" => rgb <= "000000";
					when "10000011010100111" => rgb <= "000000";
					when "10000011010101000" => rgb <= "000000";
					when "10000011010101001" => rgb <= "000000";
					when "10000011010101010" => rgb <= "000000";
					when "10000011010101011" => rgb <= "000000";
					when "10000011010101100" => rgb <= "000000";
					when "10000011010101101" => rgb <= "000000";
					when "10000011010101110" => rgb <= "000000";
					when "10000011010101111" => rgb <= "000000";
					when "10000011010110000" => rgb <= "000000";
					when "10000011010110001" => rgb <= "000000";
					when "10000011010110010" => rgb <= "000000";
					when "10000011010110011" => rgb <= "000000";
					when "10000011010110100" => rgb <= "000000";
					when "10000011010110101" => rgb <= "000000";
					when "10000011010110110" => rgb <= "000000";
					when "10000011010110111" => rgb <= "000000";
					when "10000011010111000" => rgb <= "000000";
					when "10000011010111001" => rgb <= "000000";
					when "10000011010111010" => rgb <= "000000";
					when "10000011010111011" => rgb <= "000000";
					when "10000011010111100" => rgb <= "000000";
					when "10000011010111101" => rgb <= "000000";
					when "10000011010111110" => rgb <= "000000";
					when "10000011010111111" => rgb <= "000000";
					when "10000011011000000" => rgb <= "000000";
					when "10000011011000001" => rgb <= "000000";
					when "10000011011000010" => rgb <= "000000";
					when "10000011011000011" => rgb <= "000000";
					when "10000011011000100" => rgb <= "000000";
					when "10000011011000101" => rgb <= "000000";
					when "10000011011000110" => rgb <= "000000";
					when "10000011011000111" => rgb <= "000000";
					when "10000011011001000" => rgb <= "000000";
					when "10000011011001001" => rgb <= "000000";
					when "10000011011001010" => rgb <= "000000";
					when "10000011011001011" => rgb <= "000000";
					when "10000011011001100" => rgb <= "000000";
					when "10000011011001101" => rgb <= "000000";
					when "10000011011001110" => rgb <= "000000";
					when "10000011011001111" => rgb <= "000000";
					when "10000011011010000" => rgb <= "000000";
					when "10000011011010001" => rgb <= "000000";
					when "10000011011010010" => rgb <= "000000";
					when "10000011011010011" => rgb <= "000000";
					when "10000011011010100" => rgb <= "000000";
					when "10000011011010101" => rgb <= "000000";
					when "10000011011010110" => rgb <= "000000";
					when "10000011011010111" => rgb <= "000000";
					when "10000011011011000" => rgb <= "000000";
					when "10000011011011001" => rgb <= "000000";
					when "10000011011011010" => rgb <= "000000";
					when "10000011011011011" => rgb <= "000000";
					when "10000011011011100" => rgb <= "000000";
					when "10000011011011101" => rgb <= "000000";
					when "10000011011011110" => rgb <= "000000";
					when "10000011011011111" => rgb <= "000000";
					when "10000011011100000" => rgb <= "000000";
					when "10000011011100001" => rgb <= "000000";
					when "10000011011100010" => rgb <= "000000";
					when "10000011011100011" => rgb <= "000000";
					when "10000011011100100" => rgb <= "000000";
					when "10000011011100101" => rgb <= "000000";
					when "10000011011100110" => rgb <= "000000";
					when "10000011011100111" => rgb <= "000000";
					when "10000011011101000" => rgb <= "000000";
					when "10000011011101001" => rgb <= "000000";
					when "10000011011101010" => rgb <= "000000";
					when "10000011011101011" => rgb <= "000000";
					when "10000011011101100" => rgb <= "000000";
					when "10000011011101101" => rgb <= "000000";
					when "10000011011101110" => rgb <= "000000";
					when "10000011011101111" => rgb <= "000000";
					when "10000011011110000" => rgb <= "000000";
					when "10000011011110001" => rgb <= "000000";
					when "10000011011110010" => rgb <= "000000";
					when "10000011011110011" => rgb <= "000000";
					when "10000011011110100" => rgb <= "000000";
					when "10000011011110101" => rgb <= "000000";
					when "10000011011110110" => rgb <= "000000";
					when "10000011011110111" => rgb <= "000000";
					when "10000011011111000" => rgb <= "000000";
					when "10000011011111001" => rgb <= "000000";
					when "10000011011111010" => rgb <= "000000";
					when "10000011011111011" => rgb <= "000000";
					when "10000011011111100" => rgb <= "000000";
					when "10000011011111101" => rgb <= "000000";
					when "10000011011111110" => rgb <= "000000";
					when "10000011011111111" => rgb <= "000000";
					when "10000011100000000" => rgb <= "000000";
					when "10000011100000001" => rgb <= "000000";
					when "10000011100000010" => rgb <= "000000";
					when "10000011100000011" => rgb <= "000000";
					when "10000011100000100" => rgb <= "000000";
					when "10000011100000101" => rgb <= "000000";
					when "10000011100000110" => rgb <= "000000";
					when "10000011100000111" => rgb <= "000000";
					when "10000011100001000" => rgb <= "000000";
					when "10000011100001001" => rgb <= "000000";
					when "10000011100001010" => rgb <= "000000";
					when "10000011100001011" => rgb <= "000000";
					when "10000011100001100" => rgb <= "000000";
					when "10000011100001101" => rgb <= "000000";
					when "10000011100001110" => rgb <= "000000";
					when "10000011100001111" => rgb <= "000000";
					when "10000011100010000" => rgb <= "000000";
					when "10000011100010001" => rgb <= "000000";
					when "10000011100010010" => rgb <= "000000";
					when "10000011100010011" => rgb <= "000000";
					when "10000011100010100" => rgb <= "000000";
					when "10000011100010101" => rgb <= "000000";
					when "10000011100010110" => rgb <= "000000";
					when "10000011100010111" => rgb <= "000000";
					when "10000011100011000" => rgb <= "000000";
					when "10000011100011001" => rgb <= "000000";
					when "10000011100011010" => rgb <= "000000";
					when "10000011100011011" => rgb <= "000000";
					when "10000011100011100" => rgb <= "000000";
					when "10000011100011101" => rgb <= "000000";
					when "10000011100011110" => rgb <= "000000";
					when "10000011100011111" => rgb <= "000000";
					when "10000011100100000" => rgb <= "000000";
					when "10000011100100001" => rgb <= "000000";
					when "10000011100100010" => rgb <= "000000";
					when "10000011100100011" => rgb <= "000000";
					when "10000011100100100" => rgb <= "000000";
					when "10000011100100101" => rgb <= "000000";
					when "10000011100100110" => rgb <= "000000";
					when "10000011100100111" => rgb <= "000000";
					when "10000011100101000" => rgb <= "000000";
					when "10000011100101001" => rgb <= "000000";
					when "10000011100101010" => rgb <= "000000";
					when "10000011100101011" => rgb <= "000000";
					when "10000011100101100" => rgb <= "000000";
					when "10000011100101101" => rgb <= "000000";
					when "10000011100101110" => rgb <= "000000";
					when "10000011100101111" => rgb <= "000000";
					when "10000011100110000" => rgb <= "000000";
					when "10000011100110001" => rgb <= "000000";
					when "10000011100110010" => rgb <= "000000";
					when "10000011100110011" => rgb <= "000000";
					when "10000011100110100" => rgb <= "000000";
					when "10000011100110101" => rgb <= "000000";
					when "10000011100110110" => rgb <= "000000";
					when "10000011100110111" => rgb <= "000000";
					when "10000011100111000" => rgb <= "000000";
					when "10000011100111001" => rgb <= "000000";
					when "10000011100111010" => rgb <= "000000";
					when "10000011100111011" => rgb <= "000000";
					when "10000011100111100" => rgb <= "000000";
					when "10000011100111101" => rgb <= "000000";
					when "10000011100111110" => rgb <= "000000";
					when "10000011100111111" => rgb <= "000000";
					when "10000100000000000" => rgb <= "000000";
					when "10000100000000001" => rgb <= "000000";
					when "10000100000000010" => rgb <= "000000";
					when "10000100000000011" => rgb <= "000000";
					when "10000100000000100" => rgb <= "000000";
					when "10000100000000101" => rgb <= "000000";
					when "10000100000000110" => rgb <= "000000";
					when "10000100000000111" => rgb <= "000000";
					when "10000100000001000" => rgb <= "000000";
					when "10000100000001001" => rgb <= "000000";
					when "10000100000001010" => rgb <= "000000";
					when "10000100000001011" => rgb <= "000000";
					when "10000100000001100" => rgb <= "000000";
					when "10000100000001101" => rgb <= "000000";
					when "10000100000001110" => rgb <= "000000";
					when "10000100000001111" => rgb <= "000000";
					when "10000100000010000" => rgb <= "000000";
					when "10000100000010001" => rgb <= "000000";
					when "10000100000010010" => rgb <= "000000";
					when "10000100000010011" => rgb <= "000000";
					when "10000100000010100" => rgb <= "000000";
					when "10000100000010101" => rgb <= "000000";
					when "10000100000010110" => rgb <= "000000";
					when "10000100000010111" => rgb <= "000000";
					when "10000100000011000" => rgb <= "000000";
					when "10000100000011001" => rgb <= "000000";
					when "10000100000011010" => rgb <= "000000";
					when "10000100000011011" => rgb <= "000000";
					when "10000100000011100" => rgb <= "000000";
					when "10000100000011101" => rgb <= "000000";
					when "10000100000011110" => rgb <= "000000";
					when "10000100000011111" => rgb <= "000000";
					when "10000100000100000" => rgb <= "000000";
					when "10000100000100001" => rgb <= "000000";
					when "10000100000100010" => rgb <= "000000";
					when "10000100000100011" => rgb <= "000000";
					when "10000100000100100" => rgb <= "000000";
					when "10000100000100101" => rgb <= "000000";
					when "10000100000100110" => rgb <= "000000";
					when "10000100000100111" => rgb <= "000000";
					when "10000100000101000" => rgb <= "000000";
					when "10000100000101001" => rgb <= "000000";
					when "10000100000101010" => rgb <= "000000";
					when "10000100000101011" => rgb <= "000000";
					when "10000100000101100" => rgb <= "000000";
					when "10000100000101101" => rgb <= "000000";
					when "10000100000101110" => rgb <= "000000";
					when "10000100000101111" => rgb <= "000000";
					when "10000100000110000" => rgb <= "000000";
					when "10000100000110001" => rgb <= "000000";
					when "10000100000110010" => rgb <= "000000";
					when "10000100000110011" => rgb <= "000000";
					when "10000100000110100" => rgb <= "000000";
					when "10000100000110101" => rgb <= "000000";
					when "10000100000110110" => rgb <= "000000";
					when "10000100000110111" => rgb <= "000000";
					when "10000100000111000" => rgb <= "000000";
					when "10000100000111001" => rgb <= "000000";
					when "10000100000111010" => rgb <= "000000";
					when "10000100000111011" => rgb <= "000000";
					when "10000100000111100" => rgb <= "000000";
					when "10000100000111101" => rgb <= "000000";
					when "10000100000111110" => rgb <= "000000";
					when "10000100000111111" => rgb <= "000000";
					when "10000100001000000" => rgb <= "000000";
					when "10000100001000001" => rgb <= "000000";
					when "10000100001000010" => rgb <= "000000";
					when "10000100001000011" => rgb <= "000000";
					when "10000100001000100" => rgb <= "000000";
					when "10000100001000101" => rgb <= "000000";
					when "10000100001000110" => rgb <= "000000";
					when "10000100001000111" => rgb <= "000000";
					when "10000100001001000" => rgb <= "000000";
					when "10000100001001001" => rgb <= "000000";
					when "10000100001001010" => rgb <= "000000";
					when "10000100001001011" => rgb <= "000000";
					when "10000100001001100" => rgb <= "000000";
					when "10000100001001101" => rgb <= "000000";
					when "10000100001001110" => rgb <= "000000";
					when "10000100001001111" => rgb <= "000000";
					when "10000100001010000" => rgb <= "000000";
					when "10000100001010001" => rgb <= "000000";
					when "10000100001010010" => rgb <= "000000";
					when "10000100001010011" => rgb <= "000000";
					when "10000100001010100" => rgb <= "000000";
					when "10000100001010101" => rgb <= "000000";
					when "10000100001010110" => rgb <= "000000";
					when "10000100001010111" => rgb <= "000000";
					when "10000100001011000" => rgb <= "000000";
					when "10000100001011001" => rgb <= "000000";
					when "10000100001011010" => rgb <= "000000";
					when "10000100001011011" => rgb <= "000000";
					when "10000100001011100" => rgb <= "000000";
					when "10000100001011101" => rgb <= "000000";
					when "10000100001011110" => rgb <= "000000";
					when "10000100001011111" => rgb <= "000000";
					when "10000100001100000" => rgb <= "000000";
					when "10000100001100001" => rgb <= "000000";
					when "10000100001100010" => rgb <= "000000";
					when "10000100001100011" => rgb <= "000000";
					when "10000100001100100" => rgb <= "000000";
					when "10000100001100101" => rgb <= "000000";
					when "10000100001100110" => rgb <= "000000";
					when "10000100001100111" => rgb <= "000000";
					when "10000100001101000" => rgb <= "000000";
					when "10000100001101001" => rgb <= "000000";
					when "10000100001101010" => rgb <= "000000";
					when "10000100001101011" => rgb <= "000000";
					when "10000100001101100" => rgb <= "000000";
					when "10000100001101101" => rgb <= "000000";
					when "10000100001101110" => rgb <= "000000";
					when "10000100001101111" => rgb <= "000000";
					when "10000100001110000" => rgb <= "000000";
					when "10000100001110001" => rgb <= "000000";
					when "10000100001110010" => rgb <= "000000";
					when "10000100001110011" => rgb <= "000000";
					when "10000100001110100" => rgb <= "000000";
					when "10000100001110101" => rgb <= "000000";
					when "10000100001110110" => rgb <= "000000";
					when "10000100001110111" => rgb <= "000000";
					when "10000100001111000" => rgb <= "000000";
					when "10000100001111001" => rgb <= "000000";
					when "10000100001111010" => rgb <= "000000";
					when "10000100001111011" => rgb <= "000000";
					when "10000100001111100" => rgb <= "000000";
					when "10000100001111101" => rgb <= "000000";
					when "10000100001111110" => rgb <= "000000";
					when "10000100001111111" => rgb <= "000000";
					when "10000100010000000" => rgb <= "000000";
					when "10000100010000001" => rgb <= "000000";
					when "10000100010000010" => rgb <= "000000";
					when "10000100010000011" => rgb <= "000000";
					when "10000100010000100" => rgb <= "000000";
					when "10000100010000101" => rgb <= "000000";
					when "10000100010000110" => rgb <= "000000";
					when "10000100010000111" => rgb <= "000000";
					when "10000100010001000" => rgb <= "000000";
					when "10000100010001001" => rgb <= "000000";
					when "10000100010001010" => rgb <= "000000";
					when "10000100010001011" => rgb <= "000000";
					when "10000100010001100" => rgb <= "000000";
					when "10000100010001101" => rgb <= "000000";
					when "10000100010001110" => rgb <= "000000";
					when "10000100010001111" => rgb <= "000000";
					when "10000100010010000" => rgb <= "000000";
					when "10000100010010001" => rgb <= "000000";
					when "10000100010010010" => rgb <= "000000";
					when "10000100010010011" => rgb <= "000000";
					when "10000100010010100" => rgb <= "000000";
					when "10000100010010101" => rgb <= "000000";
					when "10000100010010110" => rgb <= "000000";
					when "10000100010010111" => rgb <= "000000";
					when "10000100010011000" => rgb <= "000000";
					when "10000100010011001" => rgb <= "000000";
					when "10000100010011010" => rgb <= "000000";
					when "10000100010011011" => rgb <= "000000";
					when "10000100010011100" => rgb <= "000000";
					when "10000100010011101" => rgb <= "000000";
					when "10000100010011110" => rgb <= "000000";
					when "10000100010011111" => rgb <= "000000";
					when "10000100010100000" => rgb <= "000000";
					when "10000100010100001" => rgb <= "000000";
					when "10000100010100010" => rgb <= "000000";
					when "10000100010100011" => rgb <= "000000";
					when "10000100010100100" => rgb <= "000000";
					when "10000100010100101" => rgb <= "000000";
					when "10000100010100110" => rgb <= "000000";
					when "10000100010100111" => rgb <= "000000";
					when "10000100010101000" => rgb <= "000000";
					when "10000100010101001" => rgb <= "000000";
					when "10000100010101010" => rgb <= "000000";
					when "10000100010101011" => rgb <= "000000";
					when "10000100010101100" => rgb <= "000000";
					when "10000100010101101" => rgb <= "000000";
					when "10000100010101110" => rgb <= "000000";
					when "10000100010101111" => rgb <= "000000";
					when "10000100010110000" => rgb <= "000000";
					when "10000100010110001" => rgb <= "000000";
					when "10000100010110010" => rgb <= "000000";
					when "10000100010110011" => rgb <= "000000";
					when "10000100010110100" => rgb <= "000000";
					when "10000100010110101" => rgb <= "000000";
					when "10000100010110110" => rgb <= "000000";
					when "10000100010110111" => rgb <= "000000";
					when "10000100010111000" => rgb <= "000000";
					when "10000100010111001" => rgb <= "000000";
					when "10000100010111010" => rgb <= "000000";
					when "10000100010111011" => rgb <= "000000";
					when "10000100010111100" => rgb <= "000000";
					when "10000100010111101" => rgb <= "000000";
					when "10000100010111110" => rgb <= "000000";
					when "10000100010111111" => rgb <= "000000";
					when "10000100011000000" => rgb <= "000000";
					when "10000100011000001" => rgb <= "000000";
					when "10000100011000010" => rgb <= "000000";
					when "10000100011000011" => rgb <= "000000";
					when "10000100011000100" => rgb <= "000000";
					when "10000100011000101" => rgb <= "000000";
					when "10000100011000110" => rgb <= "000000";
					when "10000100011000111" => rgb <= "000000";
					when "10000100011001000" => rgb <= "000000";
					when "10000100011001001" => rgb <= "000000";
					when "10000100011001010" => rgb <= "000000";
					when "10000100011001011" => rgb <= "000000";
					when "10000100011001100" => rgb <= "000000";
					when "10000100011001101" => rgb <= "000000";
					when "10000100011001110" => rgb <= "000000";
					when "10000100011001111" => rgb <= "000000";
					when "10000100011010000" => rgb <= "000000";
					when "10000100011010001" => rgb <= "000000";
					when "10000100011010010" => rgb <= "000000";
					when "10000100011010011" => rgb <= "000000";
					when "10000100011010100" => rgb <= "000000";
					when "10000100011010101" => rgb <= "000000";
					when "10000100011010110" => rgb <= "000000";
					when "10000100011010111" => rgb <= "000000";
					when "10000100011011000" => rgb <= "000000";
					when "10000100011011001" => rgb <= "000000";
					when "10000100011011010" => rgb <= "000000";
					when "10000100011011011" => rgb <= "000000";
					when "10000100011011100" => rgb <= "000000";
					when "10000100011011101" => rgb <= "000000";
					when "10000100011011110" => rgb <= "000000";
					when "10000100011011111" => rgb <= "000000";
					when "10000100011100000" => rgb <= "000000";
					when "10000100011100001" => rgb <= "000000";
					when "10000100011100010" => rgb <= "000000";
					when "10000100011100011" => rgb <= "000000";
					when "10000100011100100" => rgb <= "000000";
					when "10000100011100101" => rgb <= "000000";
					when "10000100011100110" => rgb <= "000000";
					when "10000100011100111" => rgb <= "000000";
					when "10000100011101000" => rgb <= "000000";
					when "10000100011101001" => rgb <= "000000";
					when "10000100011101010" => rgb <= "000000";
					when "10000100011101011" => rgb <= "000000";
					when "10000100011101100" => rgb <= "000000";
					when "10000100011101101" => rgb <= "000000";
					when "10000100011101110" => rgb <= "000000";
					when "10000100011101111" => rgb <= "000000";
					when "10000100011110000" => rgb <= "000000";
					when "10000100011110001" => rgb <= "000000";
					when "10000100011110010" => rgb <= "000000";
					when "10000100011110011" => rgb <= "000000";
					when "10000100011110100" => rgb <= "000000";
					when "10000100011110101" => rgb <= "000000";
					when "10000100011110110" => rgb <= "000000";
					when "10000100011110111" => rgb <= "000000";
					when "10000100011111000" => rgb <= "000000";
					when "10000100011111001" => rgb <= "000000";
					when "10000100011111010" => rgb <= "000000";
					when "10000100011111011" => rgb <= "000000";
					when "10000100011111100" => rgb <= "000000";
					when "10000100011111101" => rgb <= "000000";
					when "10000100011111110" => rgb <= "000000";
					when "10000100011111111" => rgb <= "000000";
					when "10000100100000000" => rgb <= "000000";
					when "10000100100000001" => rgb <= "000000";
					when "10000100100000010" => rgb <= "000000";
					when "10000100100000011" => rgb <= "000000";
					when "10000100100000100" => rgb <= "000000";
					when "10000100100000101" => rgb <= "000000";
					when "10000100100000110" => rgb <= "000000";
					when "10000100100000111" => rgb <= "000000";
					when "10000100100001000" => rgb <= "000000";
					when "10000100100001001" => rgb <= "000000";
					when "10000100100001010" => rgb <= "000000";
					when "10000100100001011" => rgb <= "000000";
					when "10000100100001100" => rgb <= "000000";
					when "10000100100001101" => rgb <= "000000";
					when "10000100100001110" => rgb <= "000000";
					when "10000100100001111" => rgb <= "000000";
					when "10000100100010000" => rgb <= "000000";
					when "10000100100010001" => rgb <= "000000";
					when "10000100100010010" => rgb <= "000000";
					when "10000100100010011" => rgb <= "000000";
					when "10000100100010100" => rgb <= "000000";
					when "10000100100010101" => rgb <= "000000";
					when "10000100100010110" => rgb <= "000000";
					when "10000100100010111" => rgb <= "000000";
					when "10000100100011000" => rgb <= "000000";
					when "10000100100011001" => rgb <= "000000";
					when "10000100100011010" => rgb <= "000000";
					when "10000100100011011" => rgb <= "000000";
					when "10000100100011100" => rgb <= "000000";
					when "10000100100011101" => rgb <= "000000";
					when "10000100100011110" => rgb <= "000000";
					when "10000100100011111" => rgb <= "000000";
					when "10000100100100000" => rgb <= "000000";
					when "10000100100100001" => rgb <= "000000";
					when "10000100100100010" => rgb <= "000000";
					when "10000100100100011" => rgb <= "000000";
					when "10000100100100100" => rgb <= "000000";
					when "10000100100100101" => rgb <= "000000";
					when "10000100100100110" => rgb <= "000000";
					when "10000100100100111" => rgb <= "000000";
					when "10000100100101000" => rgb <= "000000";
					when "10000100100101001" => rgb <= "000000";
					when "10000100100101010" => rgb <= "000000";
					when "10000100100101011" => rgb <= "000000";
					when "10000100100101100" => rgb <= "000000";
					when "10000100100101101" => rgb <= "000000";
					when "10000100100101110" => rgb <= "000000";
					when "10000100100101111" => rgb <= "000000";
					when "10000100100110000" => rgb <= "000000";
					when "10000100100110001" => rgb <= "000000";
					when "10000100100110010" => rgb <= "000000";
					when "10000100100110011" => rgb <= "000000";
					when "10000100100110100" => rgb <= "000000";
					when "10000100100110101" => rgb <= "000000";
					when "10000100100110110" => rgb <= "000000";
					when "10000100100110111" => rgb <= "000000";
					when "10000100100111000" => rgb <= "000000";
					when "10000100100111001" => rgb <= "000000";
					when "10000100100111010" => rgb <= "000000";
					when "10000100100111011" => rgb <= "000000";
					when "10000100100111100" => rgb <= "000000";
					when "10000100100111101" => rgb <= "000000";
					when "10000100100111110" => rgb <= "000000";
					when "10000100100111111" => rgb <= "000000";
					when "10000101000000000" => rgb <= "000000";
					when "10000101000000001" => rgb <= "000000";
					when "10000101000000010" => rgb <= "000000";
					when "10000101000000011" => rgb <= "000000";
					when "10000101000000100" => rgb <= "000000";
					when "10000101000000101" => rgb <= "000000";
					when "10000101000000110" => rgb <= "000000";
					when "10000101000000111" => rgb <= "000000";
					when "10000101000001000" => rgb <= "000000";
					when "10000101000001001" => rgb <= "000000";
					when "10000101000001010" => rgb <= "000000";
					when "10000101000001011" => rgb <= "000000";
					when "10000101000001100" => rgb <= "000000";
					when "10000101000001101" => rgb <= "000000";
					when "10000101000001110" => rgb <= "000000";
					when "10000101000001111" => rgb <= "000000";
					when "10000101000010000" => rgb <= "000000";
					when "10000101000010001" => rgb <= "000000";
					when "10000101000010010" => rgb <= "000000";
					when "10000101000010011" => rgb <= "000000";
					when "10000101000010100" => rgb <= "000000";
					when "10000101000010101" => rgb <= "000000";
					when "10000101000010110" => rgb <= "000000";
					when "10000101000010111" => rgb <= "000000";
					when "10000101000011000" => rgb <= "000000";
					when "10000101000011001" => rgb <= "000000";
					when "10000101000011010" => rgb <= "000000";
					when "10000101000011011" => rgb <= "000000";
					when "10000101000011100" => rgb <= "000000";
					when "10000101000011101" => rgb <= "000000";
					when "10000101000011110" => rgb <= "000000";
					when "10000101000011111" => rgb <= "000000";
					when "10000101000100000" => rgb <= "000000";
					when "10000101000100001" => rgb <= "000000";
					when "10000101000100010" => rgb <= "000000";
					when "10000101000100011" => rgb <= "000000";
					when "10000101000100100" => rgb <= "000000";
					when "10000101000100101" => rgb <= "000000";
					when "10000101000100110" => rgb <= "000000";
					when "10000101000100111" => rgb <= "000000";
					when "10000101000101000" => rgb <= "000000";
					when "10000101000101001" => rgb <= "000000";
					when "10000101000101010" => rgb <= "000000";
					when "10000101000101011" => rgb <= "000000";
					when "10000101000101100" => rgb <= "000000";
					when "10000101000101101" => rgb <= "000000";
					when "10000101000101110" => rgb <= "000000";
					when "10000101000101111" => rgb <= "000000";
					when "10000101000110000" => rgb <= "000000";
					when "10000101000110001" => rgb <= "000000";
					when "10000101000110010" => rgb <= "000000";
					when "10000101000110011" => rgb <= "000000";
					when "10000101000110100" => rgb <= "000000";
					when "10000101000110101" => rgb <= "000000";
					when "10000101000110110" => rgb <= "000000";
					when "10000101000110111" => rgb <= "000000";
					when "10000101000111000" => rgb <= "000000";
					when "10000101000111001" => rgb <= "000000";
					when "10000101000111010" => rgb <= "000000";
					when "10000101000111011" => rgb <= "000000";
					when "10000101000111100" => rgb <= "000000";
					when "10000101000111101" => rgb <= "000000";
					when "10000101000111110" => rgb <= "000000";
					when "10000101000111111" => rgb <= "000000";
					when "10000101001000000" => rgb <= "000000";
					when "10000101001000001" => rgb <= "000000";
					when "10000101001000010" => rgb <= "000000";
					when "10000101001000011" => rgb <= "000000";
					when "10000101001000100" => rgb <= "000000";
					when "10000101001000101" => rgb <= "000000";
					when "10000101001000110" => rgb <= "000000";
					when "10000101001000111" => rgb <= "000000";
					when "10000101001001000" => rgb <= "000000";
					when "10000101001001001" => rgb <= "000000";
					when "10000101001001010" => rgb <= "000000";
					when "10000101001001011" => rgb <= "000000";
					when "10000101001001100" => rgb <= "000000";
					when "10000101001001101" => rgb <= "000000";
					when "10000101001001110" => rgb <= "000000";
					when "10000101001001111" => rgb <= "000000";
					when "10000101001010000" => rgb <= "000000";
					when "10000101001010001" => rgb <= "000000";
					when "10000101001010010" => rgb <= "000000";
					when "10000101001010011" => rgb <= "000000";
					when "10000101001010100" => rgb <= "000000";
					when "10000101001010101" => rgb <= "000000";
					when "10000101001010110" => rgb <= "000000";
					when "10000101001010111" => rgb <= "000000";
					when "10000101001011000" => rgb <= "000000";
					when "10000101001011001" => rgb <= "000000";
					when "10000101001011010" => rgb <= "000000";
					when "10000101001011011" => rgb <= "000000";
					when "10000101001011100" => rgb <= "000000";
					when "10000101001011101" => rgb <= "000000";
					when "10000101001011110" => rgb <= "000000";
					when "10000101001011111" => rgb <= "000000";
					when "10000101001100000" => rgb <= "000000";
					when "10000101001100001" => rgb <= "000000";
					when "10000101001100010" => rgb <= "000000";
					when "10000101001100011" => rgb <= "000000";
					when "10000101001100100" => rgb <= "000000";
					when "10000101001100101" => rgb <= "000000";
					when "10000101001100110" => rgb <= "000000";
					when "10000101001100111" => rgb <= "000000";
					when "10000101001101000" => rgb <= "000000";
					when "10000101001101001" => rgb <= "000000";
					when "10000101001101010" => rgb <= "000000";
					when "10000101001101011" => rgb <= "000000";
					when "10000101001101100" => rgb <= "000000";
					when "10000101001101101" => rgb <= "000000";
					when "10000101001101110" => rgb <= "000000";
					when "10000101001101111" => rgb <= "000000";
					when "10000101001110000" => rgb <= "000000";
					when "10000101001110001" => rgb <= "000000";
					when "10000101001110010" => rgb <= "000000";
					when "10000101001110011" => rgb <= "000000";
					when "10000101001110100" => rgb <= "000000";
					when "10000101001110101" => rgb <= "000000";
					when "10000101001110110" => rgb <= "000000";
					when "10000101001110111" => rgb <= "000000";
					when "10000101001111000" => rgb <= "000000";
					when "10000101001111001" => rgb <= "000000";
					when "10000101001111010" => rgb <= "000000";
					when "10000101001111011" => rgb <= "000000";
					when "10000101001111100" => rgb <= "000000";
					when "10000101001111101" => rgb <= "000000";
					when "10000101001111110" => rgb <= "000000";
					when "10000101001111111" => rgb <= "000000";
					when "10000101010000000" => rgb <= "000000";
					when "10000101010000001" => rgb <= "000000";
					when "10000101010000010" => rgb <= "000000";
					when "10000101010000011" => rgb <= "000000";
					when "10000101010000100" => rgb <= "000000";
					when "10000101010000101" => rgb <= "000000";
					when "10000101010000110" => rgb <= "000000";
					when "10000101010000111" => rgb <= "000000";
					when "10000101010001000" => rgb <= "000000";
					when "10000101010001001" => rgb <= "000000";
					when "10000101010001010" => rgb <= "000000";
					when "10000101010001011" => rgb <= "000000";
					when "10000101010001100" => rgb <= "000000";
					when "10000101010001101" => rgb <= "000000";
					when "10000101010001110" => rgb <= "000000";
					when "10000101010001111" => rgb <= "000000";
					when "10000101010010000" => rgb <= "000000";
					when "10000101010010001" => rgb <= "000000";
					when "10000101010010010" => rgb <= "000000";
					when "10000101010010011" => rgb <= "000000";
					when "10000101010010100" => rgb <= "000000";
					when "10000101010010101" => rgb <= "000000";
					when "10000101010010110" => rgb <= "000000";
					when "10000101010010111" => rgb <= "000000";
					when "10000101010011000" => rgb <= "000000";
					when "10000101010011001" => rgb <= "000000";
					when "10000101010011010" => rgb <= "000000";
					when "10000101010011011" => rgb <= "000000";
					when "10000101010011100" => rgb <= "000000";
					when "10000101010011101" => rgb <= "000000";
					when "10000101010011110" => rgb <= "000000";
					when "10000101010011111" => rgb <= "000000";
					when "10000101010100000" => rgb <= "000000";
					when "10000101010100001" => rgb <= "000000";
					when "10000101010100010" => rgb <= "000000";
					when "10000101010100011" => rgb <= "000000";
					when "10000101010100100" => rgb <= "000000";
					when "10000101010100101" => rgb <= "000000";
					when "10000101010100110" => rgb <= "000000";
					when "10000101010100111" => rgb <= "000000";
					when "10000101010101000" => rgb <= "000000";
					when "10000101010101001" => rgb <= "000000";
					when "10000101010101010" => rgb <= "000000";
					when "10000101010101011" => rgb <= "000000";
					when "10000101010101100" => rgb <= "000000";
					when "10000101010101101" => rgb <= "000000";
					when "10000101010101110" => rgb <= "000000";
					when "10000101010101111" => rgb <= "000000";
					when "10000101010110000" => rgb <= "000000";
					when "10000101010110001" => rgb <= "000000";
					when "10000101010110010" => rgb <= "000000";
					when "10000101010110011" => rgb <= "000000";
					when "10000101010110100" => rgb <= "000000";
					when "10000101010110101" => rgb <= "000000";
					when "10000101010110110" => rgb <= "000000";
					when "10000101010110111" => rgb <= "000000";
					when "10000101010111000" => rgb <= "000000";
					when "10000101010111001" => rgb <= "000000";
					when "10000101010111010" => rgb <= "000000";
					when "10000101010111011" => rgb <= "000000";
					when "10000101010111100" => rgb <= "000000";
					when "10000101010111101" => rgb <= "000000";
					when "10000101010111110" => rgb <= "000000";
					when "10000101010111111" => rgb <= "000000";
					when "10000101011000000" => rgb <= "000000";
					when "10000101011000001" => rgb <= "000000";
					when "10000101011000010" => rgb <= "000000";
					when "10000101011000011" => rgb <= "000000";
					when "10000101011000100" => rgb <= "000000";
					when "10000101011000101" => rgb <= "000000";
					when "10000101011000110" => rgb <= "000000";
					when "10000101011000111" => rgb <= "000000";
					when "10000101011001000" => rgb <= "000000";
					when "10000101011001001" => rgb <= "000000";
					when "10000101011001010" => rgb <= "000000";
					when "10000101011001011" => rgb <= "000000";
					when "10000101011001100" => rgb <= "000000";
					when "10000101011001101" => rgb <= "000000";
					when "10000101011001110" => rgb <= "000000";
					when "10000101011001111" => rgb <= "000000";
					when "10000101011010000" => rgb <= "000000";
					when "10000101011010001" => rgb <= "000000";
					when "10000101011010010" => rgb <= "000000";
					when "10000101011010011" => rgb <= "000000";
					when "10000101011010100" => rgb <= "000000";
					when "10000101011010101" => rgb <= "000000";
					when "10000101011010110" => rgb <= "000000";
					when "10000101011010111" => rgb <= "000000";
					when "10000101011011000" => rgb <= "000000";
					when "10000101011011001" => rgb <= "000000";
					when "10000101011011010" => rgb <= "000000";
					when "10000101011011011" => rgb <= "000000";
					when "10000101011011100" => rgb <= "000000";
					when "10000101011011101" => rgb <= "000000";
					when "10000101011011110" => rgb <= "000000";
					when "10000101011011111" => rgb <= "000000";
					when "10000101011100000" => rgb <= "000000";
					when "10000101011100001" => rgb <= "000000";
					when "10000101011100010" => rgb <= "000000";
					when "10000101011100011" => rgb <= "000000";
					when "10000101011100100" => rgb <= "000000";
					when "10000101011100101" => rgb <= "000000";
					when "10000101011100110" => rgb <= "000000";
					when "10000101011100111" => rgb <= "000000";
					when "10000101011101000" => rgb <= "000000";
					when "10000101011101001" => rgb <= "000000";
					when "10000101011101010" => rgb <= "000000";
					when "10000101011101011" => rgb <= "000000";
					when "10000101011101100" => rgb <= "000000";
					when "10000101011101101" => rgb <= "000000";
					when "10000101011101110" => rgb <= "000000";
					when "10000101011101111" => rgb <= "000000";
					when "10000101011110000" => rgb <= "000000";
					when "10000101011110001" => rgb <= "000000";
					when "10000101011110010" => rgb <= "000000";
					when "10000101011110011" => rgb <= "000000";
					when "10000101011110100" => rgb <= "000000";
					when "10000101011110101" => rgb <= "000000";
					when "10000101011110110" => rgb <= "000000";
					when "10000101011110111" => rgb <= "000000";
					when "10000101011111000" => rgb <= "000000";
					when "10000101011111001" => rgb <= "000000";
					when "10000101011111010" => rgb <= "000000";
					when "10000101011111011" => rgb <= "000000";
					when "10000101011111100" => rgb <= "000000";
					when "10000101011111101" => rgb <= "000000";
					when "10000101011111110" => rgb <= "000000";
					when "10000101011111111" => rgb <= "000000";
					when "10000101100000000" => rgb <= "000000";
					when "10000101100000001" => rgb <= "000000";
					when "10000101100000010" => rgb <= "000000";
					when "10000101100000011" => rgb <= "000000";
					when "10000101100000100" => rgb <= "000000";
					when "10000101100000101" => rgb <= "000000";
					when "10000101100000110" => rgb <= "000000";
					when "10000101100000111" => rgb <= "000000";
					when "10000101100001000" => rgb <= "000000";
					when "10000101100001001" => rgb <= "000000";
					when "10000101100001010" => rgb <= "000000";
					when "10000101100001011" => rgb <= "000000";
					when "10000101100001100" => rgb <= "000000";
					when "10000101100001101" => rgb <= "000000";
					when "10000101100001110" => rgb <= "000000";
					when "10000101100001111" => rgb <= "000000";
					when "10000101100010000" => rgb <= "000000";
					when "10000101100010001" => rgb <= "000000";
					when "10000101100010010" => rgb <= "000000";
					when "10000101100010011" => rgb <= "000000";
					when "10000101100010100" => rgb <= "000000";
					when "10000101100010101" => rgb <= "000000";
					when "10000101100010110" => rgb <= "000000";
					when "10000101100010111" => rgb <= "000000";
					when "10000101100011000" => rgb <= "000000";
					when "10000101100011001" => rgb <= "000000";
					when "10000101100011010" => rgb <= "000000";
					when "10000101100011011" => rgb <= "000000";
					when "10000101100011100" => rgb <= "000000";
					when "10000101100011101" => rgb <= "000000";
					when "10000101100011110" => rgb <= "000000";
					when "10000101100011111" => rgb <= "000000";
					when "10000101100100000" => rgb <= "000000";
					when "10000101100100001" => rgb <= "000000";
					when "10000101100100010" => rgb <= "000000";
					when "10000101100100011" => rgb <= "000000";
					when "10000101100100100" => rgb <= "000000";
					when "10000101100100101" => rgb <= "000000";
					when "10000101100100110" => rgb <= "000000";
					when "10000101100100111" => rgb <= "000000";
					when "10000101100101000" => rgb <= "000000";
					when "10000101100101001" => rgb <= "000000";
					when "10000101100101010" => rgb <= "000000";
					when "10000101100101011" => rgb <= "000000";
					when "10000101100101100" => rgb <= "000000";
					when "10000101100101101" => rgb <= "000000";
					when "10000101100101110" => rgb <= "000000";
					when "10000101100101111" => rgb <= "000000";
					when "10000101100110000" => rgb <= "000000";
					when "10000101100110001" => rgb <= "000000";
					when "10000101100110010" => rgb <= "000000";
					when "10000101100110011" => rgb <= "000000";
					when "10000101100110100" => rgb <= "000000";
					when "10000101100110101" => rgb <= "000000";
					when "10000101100110110" => rgb <= "000000";
					when "10000101100110111" => rgb <= "000000";
					when "10000101100111000" => rgb <= "000000";
					when "10000101100111001" => rgb <= "000000";
					when "10000101100111010" => rgb <= "000000";
					when "10000101100111011" => rgb <= "000000";
					when "10000101100111100" => rgb <= "000000";
					when "10000101100111101" => rgb <= "000000";
					when "10000101100111110" => rgb <= "000000";
					when "10000101100111111" => rgb <= "000000";
					when "10000110000000000" => rgb <= "000000";
					when "10000110000000001" => rgb <= "000000";
					when "10000110000000010" => rgb <= "000000";
					when "10000110000000011" => rgb <= "000000";
					when "10000110000000100" => rgb <= "000000";
					when "10000110000000101" => rgb <= "000000";
					when "10000110000000110" => rgb <= "000000";
					when "10000110000000111" => rgb <= "000000";
					when "10000110000001000" => rgb <= "000000";
					when "10000110000001001" => rgb <= "000000";
					when "10000110000001010" => rgb <= "000000";
					when "10000110000001011" => rgb <= "000000";
					when "10000110000001100" => rgb <= "000000";
					when "10000110000001101" => rgb <= "000000";
					when "10000110000001110" => rgb <= "000000";
					when "10000110000001111" => rgb <= "000000";
					when "10000110000010000" => rgb <= "000000";
					when "10000110000010001" => rgb <= "000000";
					when "10000110000010010" => rgb <= "000000";
					when "10000110000010011" => rgb <= "000000";
					when "10000110000010100" => rgb <= "000000";
					when "10000110000010101" => rgb <= "000000";
					when "10000110000010110" => rgb <= "000000";
					when "10000110000010111" => rgb <= "000000";
					when "10000110000011000" => rgb <= "000000";
					when "10000110000011001" => rgb <= "000000";
					when "10000110000011010" => rgb <= "000000";
					when "10000110000011011" => rgb <= "000000";
					when "10000110000011100" => rgb <= "000000";
					when "10000110000011101" => rgb <= "000000";
					when "10000110000011110" => rgb <= "000000";
					when "10000110000011111" => rgb <= "000000";
					when "10000110000100000" => rgb <= "000000";
					when "10000110000100001" => rgb <= "000000";
					when "10000110000100010" => rgb <= "000000";
					when "10000110000100011" => rgb <= "000000";
					when "10000110000100100" => rgb <= "000000";
					when "10000110000100101" => rgb <= "000000";
					when "10000110000100110" => rgb <= "000000";
					when "10000110000100111" => rgb <= "000000";
					when "10000110000101000" => rgb <= "000000";
					when "10000110000101001" => rgb <= "000000";
					when "10000110000101010" => rgb <= "000000";
					when "10000110000101011" => rgb <= "000000";
					when "10000110000101100" => rgb <= "000000";
					when "10000110000101101" => rgb <= "000000";
					when "10000110000101110" => rgb <= "000000";
					when "10000110000101111" => rgb <= "000000";
					when "10000110000110000" => rgb <= "000000";
					when "10000110000110001" => rgb <= "000000";
					when "10000110000110010" => rgb <= "000000";
					when "10000110000110011" => rgb <= "000000";
					when "10000110000110100" => rgb <= "000000";
					when "10000110000110101" => rgb <= "000000";
					when "10000110000110110" => rgb <= "000000";
					when "10000110000110111" => rgb <= "000000";
					when "10000110000111000" => rgb <= "000000";
					when "10000110000111001" => rgb <= "000000";
					when "10000110000111010" => rgb <= "000000";
					when "10000110000111011" => rgb <= "000000";
					when "10000110000111100" => rgb <= "000000";
					when "10000110000111101" => rgb <= "000000";
					when "10000110000111110" => rgb <= "000000";
					when "10000110000111111" => rgb <= "000000";
					when "10000110001000000" => rgb <= "000000";
					when "10000110001000001" => rgb <= "000000";
					when "10000110001000010" => rgb <= "000000";
					when "10000110001000011" => rgb <= "000000";
					when "10000110001000100" => rgb <= "000000";
					when "10000110001000101" => rgb <= "000000";
					when "10000110001000110" => rgb <= "000000";
					when "10000110001000111" => rgb <= "000000";
					when "10000110001001000" => rgb <= "000000";
					when "10000110001001001" => rgb <= "000000";
					when "10000110001001010" => rgb <= "000000";
					when "10000110001001011" => rgb <= "000000";
					when "10000110001001100" => rgb <= "000000";
					when "10000110001001101" => rgb <= "000000";
					when "10000110001001110" => rgb <= "000000";
					when "10000110001001111" => rgb <= "000000";
					when "10000110001010000" => rgb <= "000000";
					when "10000110001010001" => rgb <= "000000";
					when "10000110001010010" => rgb <= "000000";
					when "10000110001010011" => rgb <= "000000";
					when "10000110001010100" => rgb <= "000000";
					when "10000110001010101" => rgb <= "000000";
					when "10000110001010110" => rgb <= "000000";
					when "10000110001010111" => rgb <= "000000";
					when "10000110001011000" => rgb <= "000000";
					when "10000110001011001" => rgb <= "000000";
					when "10000110001011010" => rgb <= "000000";
					when "10000110001011011" => rgb <= "000000";
					when "10000110001011100" => rgb <= "000000";
					when "10000110001011101" => rgb <= "000000";
					when "10000110001011110" => rgb <= "000000";
					when "10000110001011111" => rgb <= "000000";
					when "10000110001100000" => rgb <= "000000";
					when "10000110001100001" => rgb <= "000000";
					when "10000110001100010" => rgb <= "000000";
					when "10000110001100011" => rgb <= "000000";
					when "10000110001100100" => rgb <= "000000";
					when "10000110001100101" => rgb <= "000000";
					when "10000110001100110" => rgb <= "000000";
					when "10000110001100111" => rgb <= "000000";
					when "10000110001101000" => rgb <= "000000";
					when "10000110001101001" => rgb <= "000000";
					when "10000110001101010" => rgb <= "000000";
					when "10000110001101011" => rgb <= "000000";
					when "10000110001101100" => rgb <= "000000";
					when "10000110001101101" => rgb <= "000000";
					when "10000110001101110" => rgb <= "000000";
					when "10000110001101111" => rgb <= "000000";
					when "10000110001110000" => rgb <= "000000";
					when "10000110001110001" => rgb <= "000000";
					when "10000110001110010" => rgb <= "000000";
					when "10000110001110011" => rgb <= "000000";
					when "10000110001110100" => rgb <= "000000";
					when "10000110001110101" => rgb <= "000000";
					when "10000110001110110" => rgb <= "000000";
					when "10000110001110111" => rgb <= "000000";
					when "10000110001111000" => rgb <= "000000";
					when "10000110001111001" => rgb <= "000000";
					when "10000110001111010" => rgb <= "000000";
					when "10000110001111011" => rgb <= "000000";
					when "10000110001111100" => rgb <= "000000";
					when "10000110001111101" => rgb <= "000000";
					when "10000110001111110" => rgb <= "000000";
					when "10000110001111111" => rgb <= "000000";
					when "10000110010000000" => rgb <= "000000";
					when "10000110010000001" => rgb <= "000000";
					when "10000110010000010" => rgb <= "000000";
					when "10000110010000011" => rgb <= "000000";
					when "10000110010000100" => rgb <= "000000";
					when "10000110010000101" => rgb <= "000000";
					when "10000110010000110" => rgb <= "000000";
					when "10000110010000111" => rgb <= "000000";
					when "10000110010001000" => rgb <= "000000";
					when "10000110010001001" => rgb <= "000000";
					when "10000110010001010" => rgb <= "000000";
					when "10000110010001011" => rgb <= "000000";
					when "10000110010001100" => rgb <= "000000";
					when "10000110010001101" => rgb <= "000000";
					when "10000110010001110" => rgb <= "000000";
					when "10000110010001111" => rgb <= "000000";
					when "10000110010010000" => rgb <= "000000";
					when "10000110010010001" => rgb <= "000000";
					when "10000110010010010" => rgb <= "000000";
					when "10000110010010011" => rgb <= "000000";
					when "10000110010010100" => rgb <= "000000";
					when "10000110010010101" => rgb <= "000000";
					when "10000110010010110" => rgb <= "000000";
					when "10000110010010111" => rgb <= "000000";
					when "10000110010011000" => rgb <= "000000";
					when "10000110010011001" => rgb <= "000000";
					when "10000110010011010" => rgb <= "000000";
					when "10000110010011011" => rgb <= "000000";
					when "10000110010011100" => rgb <= "000000";
					when "10000110010011101" => rgb <= "000000";
					when "10000110010011110" => rgb <= "000000";
					when "10000110010011111" => rgb <= "000000";
					when "10000110010100000" => rgb <= "000000";
					when "10000110010100001" => rgb <= "000000";
					when "10000110010100010" => rgb <= "000000";
					when "10000110010100011" => rgb <= "000000";
					when "10000110010100100" => rgb <= "000000";
					when "10000110010100101" => rgb <= "000000";
					when "10000110010100110" => rgb <= "000000";
					when "10000110010100111" => rgb <= "000000";
					when "10000110010101000" => rgb <= "000000";
					when "10000110010101001" => rgb <= "000000";
					when "10000110010101010" => rgb <= "000000";
					when "10000110010101011" => rgb <= "000000";
					when "10000110010101100" => rgb <= "000000";
					when "10000110010101101" => rgb <= "000000";
					when "10000110010101110" => rgb <= "000000";
					when "10000110010101111" => rgb <= "000000";
					when "10000110010110000" => rgb <= "000000";
					when "10000110010110001" => rgb <= "000000";
					when "10000110010110010" => rgb <= "000000";
					when "10000110010110011" => rgb <= "000000";
					when "10000110010110100" => rgb <= "000000";
					when "10000110010110101" => rgb <= "000000";
					when "10000110010110110" => rgb <= "000000";
					when "10000110010110111" => rgb <= "000000";
					when "10000110010111000" => rgb <= "000000";
					when "10000110010111001" => rgb <= "000000";
					when "10000110010111010" => rgb <= "000000";
					when "10000110010111011" => rgb <= "000000";
					when "10000110010111100" => rgb <= "000000";
					when "10000110010111101" => rgb <= "000000";
					when "10000110010111110" => rgb <= "000000";
					when "10000110010111111" => rgb <= "000000";
					when "10000110011000000" => rgb <= "000000";
					when "10000110011000001" => rgb <= "000000";
					when "10000110011000010" => rgb <= "000000";
					when "10000110011000011" => rgb <= "000000";
					when "10000110011000100" => rgb <= "000000";
					when "10000110011000101" => rgb <= "000000";
					when "10000110011000110" => rgb <= "000000";
					when "10000110011000111" => rgb <= "000000";
					when "10000110011001000" => rgb <= "000000";
					when "10000110011001001" => rgb <= "000000";
					when "10000110011001010" => rgb <= "000000";
					when "10000110011001011" => rgb <= "000000";
					when "10000110011001100" => rgb <= "000000";
					when "10000110011001101" => rgb <= "000000";
					when "10000110011001110" => rgb <= "000000";
					when "10000110011001111" => rgb <= "000000";
					when "10000110011010000" => rgb <= "000000";
					when "10000110011010001" => rgb <= "000000";
					when "10000110011010010" => rgb <= "000000";
					when "10000110011010011" => rgb <= "000000";
					when "10000110011010100" => rgb <= "000000";
					when "10000110011010101" => rgb <= "000000";
					when "10000110011010110" => rgb <= "000000";
					when "10000110011010111" => rgb <= "000000";
					when "10000110011011000" => rgb <= "000000";
					when "10000110011011001" => rgb <= "000000";
					when "10000110011011010" => rgb <= "000000";
					when "10000110011011011" => rgb <= "000000";
					when "10000110011011100" => rgb <= "000000";
					when "10000110011011101" => rgb <= "000000";
					when "10000110011011110" => rgb <= "000000";
					when "10000110011011111" => rgb <= "000000";
					when "10000110011100000" => rgb <= "000000";
					when "10000110011100001" => rgb <= "000000";
					when "10000110011100010" => rgb <= "000000";
					when "10000110011100011" => rgb <= "000000";
					when "10000110011100100" => rgb <= "000000";
					when "10000110011100101" => rgb <= "000000";
					when "10000110011100110" => rgb <= "000000";
					when "10000110011100111" => rgb <= "000000";
					when "10000110011101000" => rgb <= "000000";
					when "10000110011101001" => rgb <= "000000";
					when "10000110011101010" => rgb <= "000000";
					when "10000110011101011" => rgb <= "000000";
					when "10000110011101100" => rgb <= "000000";
					when "10000110011101101" => rgb <= "000000";
					when "10000110011101110" => rgb <= "000000";
					when "10000110011101111" => rgb <= "000000";
					when "10000110011110000" => rgb <= "000000";
					when "10000110011110001" => rgb <= "000000";
					when "10000110011110010" => rgb <= "000000";
					when "10000110011110011" => rgb <= "000000";
					when "10000110011110100" => rgb <= "000000";
					when "10000110011110101" => rgb <= "000000";
					when "10000110011110110" => rgb <= "000000";
					when "10000110011110111" => rgb <= "000000";
					when "10000110011111000" => rgb <= "000000";
					when "10000110011111001" => rgb <= "000000";
					when "10000110011111010" => rgb <= "000000";
					when "10000110011111011" => rgb <= "000000";
					when "10000110011111100" => rgb <= "000000";
					when "10000110011111101" => rgb <= "000000";
					when "10000110011111110" => rgb <= "000000";
					when "10000110011111111" => rgb <= "000000";
					when "10000110100000000" => rgb <= "000000";
					when "10000110100000001" => rgb <= "000000";
					when "10000110100000010" => rgb <= "000000";
					when "10000110100000011" => rgb <= "000000";
					when "10000110100000100" => rgb <= "000000";
					when "10000110100000101" => rgb <= "000000";
					when "10000110100000110" => rgb <= "000000";
					when "10000110100000111" => rgb <= "000000";
					when "10000110100001000" => rgb <= "000000";
					when "10000110100001001" => rgb <= "000000";
					when "10000110100001010" => rgb <= "000000";
					when "10000110100001011" => rgb <= "000000";
					when "10000110100001100" => rgb <= "000000";
					when "10000110100001101" => rgb <= "000000";
					when "10000110100001110" => rgb <= "000000";
					when "10000110100001111" => rgb <= "000000";
					when "10000110100010000" => rgb <= "000000";
					when "10000110100010001" => rgb <= "000000";
					when "10000110100010010" => rgb <= "000000";
					when "10000110100010011" => rgb <= "000000";
					when "10000110100010100" => rgb <= "000000";
					when "10000110100010101" => rgb <= "000000";
					when "10000110100010110" => rgb <= "000000";
					when "10000110100010111" => rgb <= "000000";
					when "10000110100011000" => rgb <= "000000";
					when "10000110100011001" => rgb <= "000000";
					when "10000110100011010" => rgb <= "000000";
					when "10000110100011011" => rgb <= "000000";
					when "10000110100011100" => rgb <= "000000";
					when "10000110100011101" => rgb <= "000000";
					when "10000110100011110" => rgb <= "000000";
					when "10000110100011111" => rgb <= "000000";
					when "10000110100100000" => rgb <= "000000";
					when "10000110100100001" => rgb <= "000000";
					when "10000110100100010" => rgb <= "000000";
					when "10000110100100011" => rgb <= "000000";
					when "10000110100100100" => rgb <= "000000";
					when "10000110100100101" => rgb <= "000000";
					when "10000110100100110" => rgb <= "000000";
					when "10000110100100111" => rgb <= "000000";
					when "10000110100101000" => rgb <= "000000";
					when "10000110100101001" => rgb <= "000000";
					when "10000110100101010" => rgb <= "000000";
					when "10000110100101011" => rgb <= "000000";
					when "10000110100101100" => rgb <= "000000";
					when "10000110100101101" => rgb <= "000000";
					when "10000110100101110" => rgb <= "000000";
					when "10000110100101111" => rgb <= "000000";
					when "10000110100110000" => rgb <= "000000";
					when "10000110100110001" => rgb <= "000000";
					when "10000110100110010" => rgb <= "000000";
					when "10000110100110011" => rgb <= "000000";
					when "10000110100110100" => rgb <= "000000";
					when "10000110100110101" => rgb <= "000000";
					when "10000110100110110" => rgb <= "000000";
					when "10000110100110111" => rgb <= "000000";
					when "10000110100111000" => rgb <= "000000";
					when "10000110100111001" => rgb <= "000000";
					when "10000110100111010" => rgb <= "000000";
					when "10000110100111011" => rgb <= "000000";
					when "10000110100111100" => rgb <= "000000";
					when "10000110100111101" => rgb <= "000000";
					when "10000110100111110" => rgb <= "000000";
					when "10000110100111111" => rgb <= "000000";
					when "10000111000000000" => rgb <= "000000";
					when "10000111000000001" => rgb <= "000000";
					when "10000111000000010" => rgb <= "000000";
					when "10000111000000011" => rgb <= "000000";
					when "10000111000000100" => rgb <= "000000";
					when "10000111000000101" => rgb <= "000000";
					when "10000111000000110" => rgb <= "000000";
					when "10000111000000111" => rgb <= "000000";
					when "10000111000001000" => rgb <= "000000";
					when "10000111000001001" => rgb <= "000000";
					when "10000111000001010" => rgb <= "000000";
					when "10000111000001011" => rgb <= "000000";
					when "10000111000001100" => rgb <= "000000";
					when "10000111000001101" => rgb <= "000000";
					when "10000111000001110" => rgb <= "000000";
					when "10000111000001111" => rgb <= "000000";
					when "10000111000010000" => rgb <= "000000";
					when "10000111000010001" => rgb <= "000000";
					when "10000111000010010" => rgb <= "000000";
					when "10000111000010011" => rgb <= "000000";
					when "10000111000010100" => rgb <= "000000";
					when "10000111000010101" => rgb <= "000000";
					when "10000111000010110" => rgb <= "000000";
					when "10000111000010111" => rgb <= "000000";
					when "10000111000011000" => rgb <= "000000";
					when "10000111000011001" => rgb <= "000000";
					when "10000111000011010" => rgb <= "000000";
					when "10000111000011011" => rgb <= "000000";
					when "10000111000011100" => rgb <= "000000";
					when "10000111000011101" => rgb <= "000000";
					when "10000111000011110" => rgb <= "000000";
					when "10000111000011111" => rgb <= "000000";
					when "10000111000100000" => rgb <= "000000";
					when "10000111000100001" => rgb <= "000000";
					when "10000111000100010" => rgb <= "000000";
					when "10000111000100011" => rgb <= "000000";
					when "10000111000100100" => rgb <= "000000";
					when "10000111000100101" => rgb <= "000000";
					when "10000111000100110" => rgb <= "000000";
					when "10000111000100111" => rgb <= "000000";
					when "10000111000101000" => rgb <= "000000";
					when "10000111000101001" => rgb <= "000000";
					when "10000111000101010" => rgb <= "000000";
					when "10000111000101011" => rgb <= "000000";
					when "10000111000101100" => rgb <= "000000";
					when "10000111000101101" => rgb <= "000000";
					when "10000111000101110" => rgb <= "000000";
					when "10000111000101111" => rgb <= "000000";
					when "10000111000110000" => rgb <= "000000";
					when "10000111000110001" => rgb <= "000000";
					when "10000111000110010" => rgb <= "000000";
					when "10000111000110011" => rgb <= "000000";
					when "10000111000110100" => rgb <= "000000";
					when "10000111000110101" => rgb <= "000000";
					when "10000111000110110" => rgb <= "000000";
					when "10000111000110111" => rgb <= "000000";
					when "10000111000111000" => rgb <= "000000";
					when "10000111000111001" => rgb <= "000000";
					when "10000111000111010" => rgb <= "000000";
					when "10000111000111011" => rgb <= "000000";
					when "10000111000111100" => rgb <= "000000";
					when "10000111000111101" => rgb <= "000000";
					when "10000111000111110" => rgb <= "000000";
					when "10000111000111111" => rgb <= "000000";
					when "10000111001000000" => rgb <= "000000";
					when "10000111001000001" => rgb <= "000000";
					when "10000111001000010" => rgb <= "000000";
					when "10000111001000011" => rgb <= "000000";
					when "10000111001000100" => rgb <= "000000";
					when "10000111001000101" => rgb <= "000000";
					when "10000111001000110" => rgb <= "000000";
					when "10000111001000111" => rgb <= "000000";
					when "10000111001001000" => rgb <= "000000";
					when "10000111001001001" => rgb <= "000000";
					when "10000111001001010" => rgb <= "000000";
					when "10000111001001011" => rgb <= "000000";
					when "10000111001001100" => rgb <= "000000";
					when "10000111001001101" => rgb <= "000000";
					when "10000111001001110" => rgb <= "000000";
					when "10000111001001111" => rgb <= "000000";
					when "10000111001010000" => rgb <= "000000";
					when "10000111001010001" => rgb <= "000000";
					when "10000111001010010" => rgb <= "000000";
					when "10000111001010011" => rgb <= "000000";
					when "10000111001010100" => rgb <= "000000";
					when "10000111001010101" => rgb <= "000000";
					when "10000111001010110" => rgb <= "000000";
					when "10000111001010111" => rgb <= "000000";
					when "10000111001011000" => rgb <= "000000";
					when "10000111001011001" => rgb <= "000000";
					when "10000111001011010" => rgb <= "000000";
					when "10000111001011011" => rgb <= "000000";
					when "10000111001011100" => rgb <= "000000";
					when "10000111001011101" => rgb <= "000000";
					when "10000111001011110" => rgb <= "000000";
					when "10000111001011111" => rgb <= "000000";
					when "10000111001100000" => rgb <= "000000";
					when "10000111001100001" => rgb <= "000000";
					when "10000111001100010" => rgb <= "000000";
					when "10000111001100011" => rgb <= "000000";
					when "10000111001100100" => rgb <= "000000";
					when "10000111001100101" => rgb <= "000000";
					when "10000111001100110" => rgb <= "000000";
					when "10000111001100111" => rgb <= "000000";
					when "10000111001101000" => rgb <= "000000";
					when "10000111001101001" => rgb <= "000000";
					when "10000111001101010" => rgb <= "000000";
					when "10000111001101011" => rgb <= "000000";
					when "10000111001101100" => rgb <= "000000";
					when "10000111001101101" => rgb <= "000000";
					when "10000111001101110" => rgb <= "000000";
					when "10000111001101111" => rgb <= "000000";
					when "10000111001110000" => rgb <= "000000";
					when "10000111001110001" => rgb <= "000000";
					when "10000111001110010" => rgb <= "000000";
					when "10000111001110011" => rgb <= "000000";
					when "10000111001110100" => rgb <= "000000";
					when "10000111001110101" => rgb <= "000000";
					when "10000111001110110" => rgb <= "000000";
					when "10000111001110111" => rgb <= "000000";
					when "10000111001111000" => rgb <= "000000";
					when "10000111001111001" => rgb <= "000000";
					when "10000111001111010" => rgb <= "000000";
					when "10000111001111011" => rgb <= "000000";
					when "10000111001111100" => rgb <= "000000";
					when "10000111001111101" => rgb <= "000000";
					when "10000111001111110" => rgb <= "000000";
					when "10000111001111111" => rgb <= "000000";
					when "10000111010000000" => rgb <= "000000";
					when "10000111010000001" => rgb <= "000000";
					when "10000111010000010" => rgb <= "000000";
					when "10000111010000011" => rgb <= "000000";
					when "10000111010000100" => rgb <= "000000";
					when "10000111010000101" => rgb <= "000000";
					when "10000111010000110" => rgb <= "000000";
					when "10000111010000111" => rgb <= "000000";
					when "10000111010001000" => rgb <= "000000";
					when "10000111010001001" => rgb <= "000000";
					when "10000111010001010" => rgb <= "000000";
					when "10000111010001011" => rgb <= "000000";
					when "10000111010001100" => rgb <= "000000";
					when "10000111010001101" => rgb <= "000000";
					when "10000111010001110" => rgb <= "000000";
					when "10000111010001111" => rgb <= "000000";
					when "10000111010010000" => rgb <= "000000";
					when "10000111010010001" => rgb <= "000000";
					when "10000111010010010" => rgb <= "000000";
					when "10000111010010011" => rgb <= "000000";
					when "10000111010010100" => rgb <= "000000";
					when "10000111010010101" => rgb <= "000000";
					when "10000111010010110" => rgb <= "000000";
					when "10000111010010111" => rgb <= "000000";
					when "10000111010011000" => rgb <= "000000";
					when "10000111010011001" => rgb <= "000000";
					when "10000111010011010" => rgb <= "000000";
					when "10000111010011011" => rgb <= "000000";
					when "10000111010011100" => rgb <= "000000";
					when "10000111010011101" => rgb <= "000000";
					when "10000111010011110" => rgb <= "000000";
					when "10000111010011111" => rgb <= "000000";
					when "10000111010100000" => rgb <= "000000";
					when "10000111010100001" => rgb <= "000000";
					when "10000111010100010" => rgb <= "000000";
					when "10000111010100011" => rgb <= "000000";
					when "10000111010100100" => rgb <= "000000";
					when "10000111010100101" => rgb <= "000000";
					when "10000111010100110" => rgb <= "000000";
					when "10000111010100111" => rgb <= "000000";
					when "10000111010101000" => rgb <= "000000";
					when "10000111010101001" => rgb <= "000000";
					when "10000111010101010" => rgb <= "000000";
					when "10000111010101011" => rgb <= "000000";
					when "10000111010101100" => rgb <= "000000";
					when "10000111010101101" => rgb <= "000000";
					when "10000111010101110" => rgb <= "000000";
					when "10000111010101111" => rgb <= "000000";
					when "10000111010110000" => rgb <= "000000";
					when "10000111010110001" => rgb <= "000000";
					when "10000111010110010" => rgb <= "000000";
					when "10000111010110011" => rgb <= "000000";
					when "10000111010110100" => rgb <= "000000";
					when "10000111010110101" => rgb <= "000000";
					when "10000111010110110" => rgb <= "000000";
					when "10000111010110111" => rgb <= "000000";
					when "10000111010111000" => rgb <= "000000";
					when "10000111010111001" => rgb <= "000000";
					when "10000111010111010" => rgb <= "000000";
					when "10000111010111011" => rgb <= "000000";
					when "10000111010111100" => rgb <= "000000";
					when "10000111010111101" => rgb <= "000000";
					when "10000111010111110" => rgb <= "000000";
					when "10000111010111111" => rgb <= "000000";
					when "10000111011000000" => rgb <= "000000";
					when "10000111011000001" => rgb <= "000000";
					when "10000111011000010" => rgb <= "000000";
					when "10000111011000011" => rgb <= "000000";
					when "10000111011000100" => rgb <= "000000";
					when "10000111011000101" => rgb <= "000000";
					when "10000111011000110" => rgb <= "000000";
					when "10000111011000111" => rgb <= "000000";
					when "10000111011001000" => rgb <= "000000";
					when "10000111011001001" => rgb <= "000000";
					when "10000111011001010" => rgb <= "000000";
					when "10000111011001011" => rgb <= "000000";
					when "10000111011001100" => rgb <= "000000";
					when "10000111011001101" => rgb <= "000000";
					when "10000111011001110" => rgb <= "000000";
					when "10000111011001111" => rgb <= "000000";
					when "10000111011010000" => rgb <= "000000";
					when "10000111011010001" => rgb <= "000000";
					when "10000111011010010" => rgb <= "000000";
					when "10000111011010011" => rgb <= "000000";
					when "10000111011010100" => rgb <= "000000";
					when "10000111011010101" => rgb <= "000000";
					when "10000111011010110" => rgb <= "000000";
					when "10000111011010111" => rgb <= "000000";
					when "10000111011011000" => rgb <= "000000";
					when "10000111011011001" => rgb <= "000000";
					when "10000111011011010" => rgb <= "000000";
					when "10000111011011011" => rgb <= "000000";
					when "10000111011011100" => rgb <= "000000";
					when "10000111011011101" => rgb <= "000000";
					when "10000111011011110" => rgb <= "000000";
					when "10000111011011111" => rgb <= "000000";
					when "10000111011100000" => rgb <= "000000";
					when "10000111011100001" => rgb <= "000000";
					when "10000111011100010" => rgb <= "000000";
					when "10000111011100011" => rgb <= "000000";
					when "10000111011100100" => rgb <= "000000";
					when "10000111011100101" => rgb <= "000000";
					when "10000111011100110" => rgb <= "000000";
					when "10000111011100111" => rgb <= "000000";
					when "10000111011101000" => rgb <= "000000";
					when "10000111011101001" => rgb <= "000000";
					when "10000111011101010" => rgb <= "000000";
					when "10000111011101011" => rgb <= "000000";
					when "10000111011101100" => rgb <= "000000";
					when "10000111011101101" => rgb <= "000000";
					when "10000111011101110" => rgb <= "000000";
					when "10000111011101111" => rgb <= "000000";
					when "10000111011110000" => rgb <= "000000";
					when "10000111011110001" => rgb <= "000000";
					when "10000111011110010" => rgb <= "000000";
					when "10000111011110011" => rgb <= "000000";
					when "10000111011110100" => rgb <= "000000";
					when "10000111011110101" => rgb <= "000000";
					when "10000111011110110" => rgb <= "000000";
					when "10000111011110111" => rgb <= "000000";
					when "10000111011111000" => rgb <= "000000";
					when "10000111011111001" => rgb <= "000000";
					when "10000111011111010" => rgb <= "000000";
					when "10000111011111011" => rgb <= "000000";
					when "10000111011111100" => rgb <= "000000";
					when "10000111011111101" => rgb <= "000000";
					when "10000111011111110" => rgb <= "000000";
					when "10000111011111111" => rgb <= "000000";
					when "10000111100000000" => rgb <= "000000";
					when "10000111100000001" => rgb <= "000000";
					when "10000111100000010" => rgb <= "000000";
					when "10000111100000011" => rgb <= "000000";
					when "10000111100000100" => rgb <= "000000";
					when "10000111100000101" => rgb <= "000000";
					when "10000111100000110" => rgb <= "000000";
					when "10000111100000111" => rgb <= "000000";
					when "10000111100001000" => rgb <= "000000";
					when "10000111100001001" => rgb <= "000000";
					when "10000111100001010" => rgb <= "000000";
					when "10000111100001011" => rgb <= "000000";
					when "10000111100001100" => rgb <= "000000";
					when "10000111100001101" => rgb <= "000000";
					when "10000111100001110" => rgb <= "000000";
					when "10000111100001111" => rgb <= "000000";
					when "10000111100010000" => rgb <= "000000";
					when "10000111100010001" => rgb <= "000000";
					when "10000111100010010" => rgb <= "000000";
					when "10000111100010011" => rgb <= "000000";
					when "10000111100010100" => rgb <= "000000";
					when "10000111100010101" => rgb <= "000000";
					when "10000111100010110" => rgb <= "000000";
					when "10000111100010111" => rgb <= "000000";
					when "10000111100011000" => rgb <= "000000";
					when "10000111100011001" => rgb <= "000000";
					when "10000111100011010" => rgb <= "000000";
					when "10000111100011011" => rgb <= "000000";
					when "10000111100011100" => rgb <= "000000";
					when "10000111100011101" => rgb <= "000000";
					when "10000111100011110" => rgb <= "000000";
					when "10000111100011111" => rgb <= "000000";
					when "10000111100100000" => rgb <= "000000";
					when "10000111100100001" => rgb <= "000000";
					when "10000111100100010" => rgb <= "000000";
					when "10000111100100011" => rgb <= "000000";
					when "10000111100100100" => rgb <= "000000";
					when "10000111100100101" => rgb <= "000000";
					when "10000111100100110" => rgb <= "000000";
					when "10000111100100111" => rgb <= "000000";
					when "10000111100101000" => rgb <= "000000";
					when "10000111100101001" => rgb <= "000000";
					when "10000111100101010" => rgb <= "000000";
					when "10000111100101011" => rgb <= "000000";
					when "10000111100101100" => rgb <= "000000";
					when "10000111100101101" => rgb <= "000000";
					when "10000111100101110" => rgb <= "000000";
					when "10000111100101111" => rgb <= "000000";
					when "10000111100110000" => rgb <= "000000";
					when "10000111100110001" => rgb <= "000000";
					when "10000111100110010" => rgb <= "000000";
					when "10000111100110011" => rgb <= "000000";
					when "10000111100110100" => rgb <= "000000";
					when "10000111100110101" => rgb <= "000000";
					when "10000111100110110" => rgb <= "000000";
					when "10000111100110111" => rgb <= "000000";
					when "10000111100111000" => rgb <= "000000";
					when "10000111100111001" => rgb <= "000000";
					when "10000111100111010" => rgb <= "000000";
					when "10000111100111011" => rgb <= "000000";
					when "10000111100111100" => rgb <= "000000";
					when "10000111100111101" => rgb <= "000000";
					when "10000111100111110" => rgb <= "000000";
					when "10000111100111111" => rgb <= "000000";
					when "10001000000000000" => rgb <= "000000";
					when "10001000000000001" => rgb <= "000000";
					when "10001000000000010" => rgb <= "000000";
					when "10001000000000011" => rgb <= "000000";
					when "10001000000000100" => rgb <= "000000";
					when "10001000000000101" => rgb <= "000000";
					when "10001000000000110" => rgb <= "000000";
					when "10001000000000111" => rgb <= "000000";
					when "10001000000001000" => rgb <= "000000";
					when "10001000000001001" => rgb <= "000000";
					when "10001000000001010" => rgb <= "000000";
					when "10001000000001011" => rgb <= "000000";
					when "10001000000001100" => rgb <= "000000";
					when "10001000000001101" => rgb <= "000000";
					when "10001000000001110" => rgb <= "000000";
					when "10001000000001111" => rgb <= "000000";
					when "10001000000010000" => rgb <= "000000";
					when "10001000000010001" => rgb <= "000000";
					when "10001000000010010" => rgb <= "000000";
					when "10001000000010011" => rgb <= "000000";
					when "10001000000010100" => rgb <= "000000";
					when "10001000000010101" => rgb <= "000000";
					when "10001000000010110" => rgb <= "000000";
					when "10001000000010111" => rgb <= "000000";
					when "10001000000011000" => rgb <= "000000";
					when "10001000000011001" => rgb <= "000000";
					when "10001000000011010" => rgb <= "000000";
					when "10001000000011011" => rgb <= "000000";
					when "10001000000011100" => rgb <= "000000";
					when "10001000000011101" => rgb <= "000000";
					when "10001000000011110" => rgb <= "000000";
					when "10001000000011111" => rgb <= "000000";
					when "10001000000100000" => rgb <= "000000";
					when "10001000000100001" => rgb <= "000000";
					when "10001000000100010" => rgb <= "000000";
					when "10001000000100011" => rgb <= "000000";
					when "10001000000100100" => rgb <= "000000";
					when "10001000000100101" => rgb <= "000000";
					when "10001000000100110" => rgb <= "000000";
					when "10001000000100111" => rgb <= "000000";
					when "10001000000101000" => rgb <= "000000";
					when "10001000000101001" => rgb <= "000000";
					when "10001000000101010" => rgb <= "000000";
					when "10001000000101011" => rgb <= "000000";
					when "10001000000101100" => rgb <= "000000";
					when "10001000000101101" => rgb <= "000000";
					when "10001000000101110" => rgb <= "000000";
					when "10001000000101111" => rgb <= "000000";
					when "10001000000110000" => rgb <= "000000";
					when "10001000000110001" => rgb <= "000000";
					when "10001000000110010" => rgb <= "000000";
					when "10001000000110011" => rgb <= "000000";
					when "10001000000110100" => rgb <= "000000";
					when "10001000000110101" => rgb <= "000000";
					when "10001000000110110" => rgb <= "000000";
					when "10001000000110111" => rgb <= "000000";
					when "10001000000111000" => rgb <= "000000";
					when "10001000000111001" => rgb <= "000000";
					when "10001000000111010" => rgb <= "000000";
					when "10001000000111011" => rgb <= "000000";
					when "10001000000111100" => rgb <= "000000";
					when "10001000000111101" => rgb <= "000000";
					when "10001000000111110" => rgb <= "000000";
					when "10001000000111111" => rgb <= "000000";
					when "10001000001000000" => rgb <= "000000";
					when "10001000001000001" => rgb <= "000000";
					when "10001000001000010" => rgb <= "000000";
					when "10001000001000011" => rgb <= "000000";
					when "10001000001000100" => rgb <= "000000";
					when "10001000001000101" => rgb <= "000000";
					when "10001000001000110" => rgb <= "000000";
					when "10001000001000111" => rgb <= "000000";
					when "10001000001001000" => rgb <= "000000";
					when "10001000001001001" => rgb <= "000000";
					when "10001000001001010" => rgb <= "000000";
					when "10001000001001011" => rgb <= "000000";
					when "10001000001001100" => rgb <= "000000";
					when "10001000001001101" => rgb <= "000000";
					when "10001000001001110" => rgb <= "000000";
					when "10001000001001111" => rgb <= "000000";
					when "10001000001010000" => rgb <= "000000";
					when "10001000001010001" => rgb <= "000000";
					when "10001000001010010" => rgb <= "000000";
					when "10001000001010011" => rgb <= "000000";
					when "10001000001010100" => rgb <= "000000";
					when "10001000001010101" => rgb <= "000000";
					when "10001000001010110" => rgb <= "000000";
					when "10001000001010111" => rgb <= "000000";
					when "10001000001011000" => rgb <= "000000";
					when "10001000001011001" => rgb <= "000000";
					when "10001000001011010" => rgb <= "000000";
					when "10001000001011011" => rgb <= "000000";
					when "10001000001011100" => rgb <= "000000";
					when "10001000001011101" => rgb <= "000000";
					when "10001000001011110" => rgb <= "000000";
					when "10001000001011111" => rgb <= "000000";
					when "10001000001100000" => rgb <= "000000";
					when "10001000001100001" => rgb <= "000000";
					when "10001000001100010" => rgb <= "000000";
					when "10001000001100011" => rgb <= "000000";
					when "10001000001100100" => rgb <= "000000";
					when "10001000001100101" => rgb <= "000000";
					when "10001000001100110" => rgb <= "000000";
					when "10001000001100111" => rgb <= "000000";
					when "10001000001101000" => rgb <= "000000";
					when "10001000001101001" => rgb <= "000000";
					when "10001000001101010" => rgb <= "000000";
					when "10001000001101011" => rgb <= "000000";
					when "10001000001101100" => rgb <= "000000";
					when "10001000001101101" => rgb <= "000000";
					when "10001000001101110" => rgb <= "000000";
					when "10001000001101111" => rgb <= "000000";
					when "10001000001110000" => rgb <= "000000";
					when "10001000001110001" => rgb <= "000000";
					when "10001000001110010" => rgb <= "000000";
					when "10001000001110011" => rgb <= "000000";
					when "10001000001110100" => rgb <= "000000";
					when "10001000001110101" => rgb <= "000000";
					when "10001000001110110" => rgb <= "000000";
					when "10001000001110111" => rgb <= "000000";
					when "10001000001111000" => rgb <= "000000";
					when "10001000001111001" => rgb <= "000000";
					when "10001000001111010" => rgb <= "000000";
					when "10001000001111011" => rgb <= "000000";
					when "10001000001111100" => rgb <= "000000";
					when "10001000001111101" => rgb <= "000000";
					when "10001000001111110" => rgb <= "000000";
					when "10001000001111111" => rgb <= "000000";
					when "10001000010000000" => rgb <= "000000";
					when "10001000010000001" => rgb <= "000000";
					when "10001000010000010" => rgb <= "000000";
					when "10001000010000011" => rgb <= "000000";
					when "10001000010000100" => rgb <= "000000";
					when "10001000010000101" => rgb <= "000000";
					when "10001000010000110" => rgb <= "000000";
					when "10001000010000111" => rgb <= "000000";
					when "10001000010001000" => rgb <= "000000";
					when "10001000010001001" => rgb <= "000000";
					when "10001000010001010" => rgb <= "000000";
					when "10001000010001011" => rgb <= "000000";
					when "10001000010001100" => rgb <= "000000";
					when "10001000010001101" => rgb <= "000000";
					when "10001000010001110" => rgb <= "000000";
					when "10001000010001111" => rgb <= "000000";
					when "10001000010010000" => rgb <= "000000";
					when "10001000010010001" => rgb <= "000000";
					when "10001000010010010" => rgb <= "000000";
					when "10001000010010011" => rgb <= "000000";
					when "10001000010010100" => rgb <= "000000";
					when "10001000010010101" => rgb <= "000000";
					when "10001000010010110" => rgb <= "000000";
					when "10001000010010111" => rgb <= "000000";
					when "10001000010011000" => rgb <= "000000";
					when "10001000010011001" => rgb <= "000000";
					when "10001000010011010" => rgb <= "000000";
					when "10001000010011011" => rgb <= "000000";
					when "10001000010011100" => rgb <= "000000";
					when "10001000010011101" => rgb <= "000000";
					when "10001000010011110" => rgb <= "000000";
					when "10001000010011111" => rgb <= "000000";
					when "10001000010100000" => rgb <= "000000";
					when "10001000010100001" => rgb <= "000000";
					when "10001000010100010" => rgb <= "000000";
					when "10001000010100011" => rgb <= "000000";
					when "10001000010100100" => rgb <= "000000";
					when "10001000010100101" => rgb <= "000000";
					when "10001000010100110" => rgb <= "000000";
					when "10001000010100111" => rgb <= "000000";
					when "10001000010101000" => rgb <= "000000";
					when "10001000010101001" => rgb <= "000000";
					when "10001000010101010" => rgb <= "000000";
					when "10001000010101011" => rgb <= "000000";
					when "10001000010101100" => rgb <= "000000";
					when "10001000010101101" => rgb <= "000000";
					when "10001000010101110" => rgb <= "000000";
					when "10001000010101111" => rgb <= "000000";
					when "10001000010110000" => rgb <= "000000";
					when "10001000010110001" => rgb <= "000000";
					when "10001000010110010" => rgb <= "000000";
					when "10001000010110011" => rgb <= "000000";
					when "10001000010110100" => rgb <= "000000";
					when "10001000010110101" => rgb <= "000000";
					when "10001000010110110" => rgb <= "000000";
					when "10001000010110111" => rgb <= "000000";
					when "10001000010111000" => rgb <= "000000";
					when "10001000010111001" => rgb <= "000000";
					when "10001000010111010" => rgb <= "000000";
					when "10001000010111011" => rgb <= "000000";
					when "10001000010111100" => rgb <= "000000";
					when "10001000010111101" => rgb <= "000000";
					when "10001000010111110" => rgb <= "000000";
					when "10001000010111111" => rgb <= "000000";
					when "10001000011000000" => rgb <= "000000";
					when "10001000011000001" => rgb <= "000000";
					when "10001000011000010" => rgb <= "000000";
					when "10001000011000011" => rgb <= "000000";
					when "10001000011000100" => rgb <= "000000";
					when "10001000011000101" => rgb <= "000000";
					when "10001000011000110" => rgb <= "000000";
					when "10001000011000111" => rgb <= "000000";
					when "10001000011001000" => rgb <= "000000";
					when "10001000011001001" => rgb <= "000000";
					when "10001000011001010" => rgb <= "000000";
					when "10001000011001011" => rgb <= "000000";
					when "10001000011001100" => rgb <= "000000";
					when "10001000011001101" => rgb <= "000000";
					when "10001000011001110" => rgb <= "000000";
					when "10001000011001111" => rgb <= "000000";
					when "10001000011010000" => rgb <= "000000";
					when "10001000011010001" => rgb <= "000000";
					when "10001000011010010" => rgb <= "000000";
					when "10001000011010011" => rgb <= "000000";
					when "10001000011010100" => rgb <= "000000";
					when "10001000011010101" => rgb <= "000000";
					when "10001000011010110" => rgb <= "000000";
					when "10001000011010111" => rgb <= "000000";
					when "10001000011011000" => rgb <= "000000";
					when "10001000011011001" => rgb <= "000000";
					when "10001000011011010" => rgb <= "000000";
					when "10001000011011011" => rgb <= "000000";
					when "10001000011011100" => rgb <= "000000";
					when "10001000011011101" => rgb <= "000000";
					when "10001000011011110" => rgb <= "000000";
					when "10001000011011111" => rgb <= "000000";
					when "10001000011100000" => rgb <= "000000";
					when "10001000011100001" => rgb <= "000000";
					when "10001000011100010" => rgb <= "000000";
					when "10001000011100011" => rgb <= "000000";
					when "10001000011100100" => rgb <= "000000";
					when "10001000011100101" => rgb <= "000000";
					when "10001000011100110" => rgb <= "000000";
					when "10001000011100111" => rgb <= "000000";
					when "10001000011101000" => rgb <= "000000";
					when "10001000011101001" => rgb <= "000000";
					when "10001000011101010" => rgb <= "000000";
					when "10001000011101011" => rgb <= "000000";
					when "10001000011101100" => rgb <= "000000";
					when "10001000011101101" => rgb <= "000000";
					when "10001000011101110" => rgb <= "000000";
					when "10001000011101111" => rgb <= "000000";
					when "10001000011110000" => rgb <= "000000";
					when "10001000011110001" => rgb <= "000000";
					when "10001000011110010" => rgb <= "000000";
					when "10001000011110011" => rgb <= "000000";
					when "10001000011110100" => rgb <= "000000";
					when "10001000011110101" => rgb <= "000000";
					when "10001000011110110" => rgb <= "000000";
					when "10001000011110111" => rgb <= "000000";
					when "10001000011111000" => rgb <= "000000";
					when "10001000011111001" => rgb <= "000000";
					when "10001000011111010" => rgb <= "000000";
					when "10001000011111011" => rgb <= "000000";
					when "10001000011111100" => rgb <= "000000";
					when "10001000011111101" => rgb <= "000000";
					when "10001000011111110" => rgb <= "000000";
					when "10001000011111111" => rgb <= "000000";
					when "10001000100000000" => rgb <= "000000";
					when "10001000100000001" => rgb <= "000000";
					when "10001000100000010" => rgb <= "000000";
					when "10001000100000011" => rgb <= "000000";
					when "10001000100000100" => rgb <= "000000";
					when "10001000100000101" => rgb <= "000000";
					when "10001000100000110" => rgb <= "000000";
					when "10001000100000111" => rgb <= "000000";
					when "10001000100001000" => rgb <= "000000";
					when "10001000100001001" => rgb <= "000000";
					when "10001000100001010" => rgb <= "000000";
					when "10001000100001011" => rgb <= "000000";
					when "10001000100001100" => rgb <= "000000";
					when "10001000100001101" => rgb <= "000000";
					when "10001000100001110" => rgb <= "000000";
					when "10001000100001111" => rgb <= "000000";
					when "10001000100010000" => rgb <= "000000";
					when "10001000100010001" => rgb <= "000000";
					when "10001000100010010" => rgb <= "000000";
					when "10001000100010011" => rgb <= "000000";
					when "10001000100010100" => rgb <= "000000";
					when "10001000100010101" => rgb <= "000000";
					when "10001000100010110" => rgb <= "000000";
					when "10001000100010111" => rgb <= "000000";
					when "10001000100011000" => rgb <= "000000";
					when "10001000100011001" => rgb <= "000000";
					when "10001000100011010" => rgb <= "000000";
					when "10001000100011011" => rgb <= "000000";
					when "10001000100011100" => rgb <= "000000";
					when "10001000100011101" => rgb <= "000000";
					when "10001000100011110" => rgb <= "000000";
					when "10001000100011111" => rgb <= "000000";
					when "10001000100100000" => rgb <= "000000";
					when "10001000100100001" => rgb <= "000000";
					when "10001000100100010" => rgb <= "000000";
					when "10001000100100011" => rgb <= "000000";
					when "10001000100100100" => rgb <= "000000";
					when "10001000100100101" => rgb <= "000000";
					when "10001000100100110" => rgb <= "000000";
					when "10001000100100111" => rgb <= "000000";
					when "10001000100101000" => rgb <= "000000";
					when "10001000100101001" => rgb <= "000000";
					when "10001000100101010" => rgb <= "000000";
					when "10001000100101011" => rgb <= "000000";
					when "10001000100101100" => rgb <= "000000";
					when "10001000100101101" => rgb <= "000000";
					when "10001000100101110" => rgb <= "000000";
					when "10001000100101111" => rgb <= "000000";
					when "10001000100110000" => rgb <= "000000";
					when "10001000100110001" => rgb <= "000000";
					when "10001000100110010" => rgb <= "000000";
					when "10001000100110011" => rgb <= "000000";
					when "10001000100110100" => rgb <= "000000";
					when "10001000100110101" => rgb <= "000000";
					when "10001000100110110" => rgb <= "000000";
					when "10001000100110111" => rgb <= "000000";
					when "10001000100111000" => rgb <= "000000";
					when "10001000100111001" => rgb <= "000000";
					when "10001000100111010" => rgb <= "000000";
					when "10001000100111011" => rgb <= "000000";
					when "10001000100111100" => rgb <= "000000";
					when "10001000100111101" => rgb <= "000000";
					when "10001000100111110" => rgb <= "000000";
					when "10001000100111111" => rgb <= "000000";
					when "10001001000000000" => rgb <= "000000";
					when "10001001000000001" => rgb <= "000000";
					when "10001001000000010" => rgb <= "000000";
					when "10001001000000011" => rgb <= "000000";
					when "10001001000000100" => rgb <= "000000";
					when "10001001000000101" => rgb <= "000000";
					when "10001001000000110" => rgb <= "000000";
					when "10001001000000111" => rgb <= "000000";
					when "10001001000001000" => rgb <= "000000";
					when "10001001000001001" => rgb <= "000000";
					when "10001001000001010" => rgb <= "000000";
					when "10001001000001011" => rgb <= "000000";
					when "10001001000001100" => rgb <= "000000";
					when "10001001000001101" => rgb <= "000000";
					when "10001001000001110" => rgb <= "000000";
					when "10001001000001111" => rgb <= "000000";
					when "10001001000010000" => rgb <= "000000";
					when "10001001000010001" => rgb <= "000000";
					when "10001001000010010" => rgb <= "000000";
					when "10001001000010011" => rgb <= "000000";
					when "10001001000010100" => rgb <= "000000";
					when "10001001000010101" => rgb <= "000000";
					when "10001001000010110" => rgb <= "000000";
					when "10001001000010111" => rgb <= "000000";
					when "10001001000011000" => rgb <= "000000";
					when "10001001000011001" => rgb <= "000000";
					when "10001001000011010" => rgb <= "000000";
					when "10001001000011011" => rgb <= "000000";
					when "10001001000011100" => rgb <= "000000";
					when "10001001000011101" => rgb <= "000000";
					when "10001001000011110" => rgb <= "000000";
					when "10001001000011111" => rgb <= "000000";
					when "10001001000100000" => rgb <= "000000";
					when "10001001000100001" => rgb <= "000000";
					when "10001001000100010" => rgb <= "000000";
					when "10001001000100011" => rgb <= "000000";
					when "10001001000100100" => rgb <= "000000";
					when "10001001000100101" => rgb <= "000000";
					when "10001001000100110" => rgb <= "000000";
					when "10001001000100111" => rgb <= "000000";
					when "10001001000101000" => rgb <= "000000";
					when "10001001000101001" => rgb <= "000000";
					when "10001001000101010" => rgb <= "000000";
					when "10001001000101011" => rgb <= "000000";
					when "10001001000101100" => rgb <= "000000";
					when "10001001000101101" => rgb <= "000000";
					when "10001001000101110" => rgb <= "000000";
					when "10001001000101111" => rgb <= "000000";
					when "10001001000110000" => rgb <= "000000";
					when "10001001000110001" => rgb <= "000000";
					when "10001001000110010" => rgb <= "000000";
					when "10001001000110011" => rgb <= "000000";
					when "10001001000110100" => rgb <= "000000";
					when "10001001000110101" => rgb <= "000000";
					when "10001001000110110" => rgb <= "000000";
					when "10001001000110111" => rgb <= "000000";
					when "10001001000111000" => rgb <= "000000";
					when "10001001000111001" => rgb <= "000000";
					when "10001001000111010" => rgb <= "000000";
					when "10001001000111011" => rgb <= "000000";
					when "10001001000111100" => rgb <= "000000";
					when "10001001000111101" => rgb <= "000000";
					when "10001001000111110" => rgb <= "000000";
					when "10001001000111111" => rgb <= "000000";
					when "10001001001000000" => rgb <= "000000";
					when "10001001001000001" => rgb <= "000000";
					when "10001001001000010" => rgb <= "000000";
					when "10001001001000011" => rgb <= "000000";
					when "10001001001000100" => rgb <= "000000";
					when "10001001001000101" => rgb <= "000000";
					when "10001001001000110" => rgb <= "000000";
					when "10001001001000111" => rgb <= "000000";
					when "10001001001001000" => rgb <= "000000";
					when "10001001001001001" => rgb <= "000000";
					when "10001001001001010" => rgb <= "000000";
					when "10001001001001011" => rgb <= "000000";
					when "10001001001001100" => rgb <= "000000";
					when "10001001001001101" => rgb <= "000000";
					when "10001001001001110" => rgb <= "000000";
					when "10001001001001111" => rgb <= "000000";
					when "10001001001010000" => rgb <= "000000";
					when "10001001001010001" => rgb <= "000000";
					when "10001001001010010" => rgb <= "000000";
					when "10001001001010011" => rgb <= "000000";
					when "10001001001010100" => rgb <= "000000";
					when "10001001001010101" => rgb <= "000000";
					when "10001001001010110" => rgb <= "000000";
					when "10001001001010111" => rgb <= "000000";
					when "10001001001011000" => rgb <= "000000";
					when "10001001001011001" => rgb <= "000000";
					when "10001001001011010" => rgb <= "000000";
					when "10001001001011011" => rgb <= "000000";
					when "10001001001011100" => rgb <= "000000";
					when "10001001001011101" => rgb <= "000000";
					when "10001001001011110" => rgb <= "000000";
					when "10001001001011111" => rgb <= "000000";
					when "10001001001100000" => rgb <= "000000";
					when "10001001001100001" => rgb <= "000000";
					when "10001001001100010" => rgb <= "000000";
					when "10001001001100011" => rgb <= "000000";
					when "10001001001100100" => rgb <= "000000";
					when "10001001001100101" => rgb <= "000000";
					when "10001001001100110" => rgb <= "000000";
					when "10001001001100111" => rgb <= "000000";
					when "10001001001101000" => rgb <= "000000";
					when "10001001001101001" => rgb <= "000000";
					when "10001001001101010" => rgb <= "000000";
					when "10001001001101011" => rgb <= "000000";
					when "10001001001101100" => rgb <= "000000";
					when "10001001001101101" => rgb <= "000000";
					when "10001001001101110" => rgb <= "000000";
					when "10001001001101111" => rgb <= "000000";
					when "10001001001110000" => rgb <= "000000";
					when "10001001001110001" => rgb <= "000000";
					when "10001001001110010" => rgb <= "000000";
					when "10001001001110011" => rgb <= "000000";
					when "10001001001110100" => rgb <= "000000";
					when "10001001001110101" => rgb <= "000000";
					when "10001001001110110" => rgb <= "000000";
					when "10001001001110111" => rgb <= "000000";
					when "10001001001111000" => rgb <= "000000";
					when "10001001001111001" => rgb <= "000000";
					when "10001001001111010" => rgb <= "000000";
					when "10001001001111011" => rgb <= "000000";
					when "10001001001111100" => rgb <= "000000";
					when "10001001001111101" => rgb <= "000000";
					when "10001001001111110" => rgb <= "000000";
					when "10001001001111111" => rgb <= "000000";
					when "10001001010000000" => rgb <= "000000";
					when "10001001010000001" => rgb <= "000000";
					when "10001001010000010" => rgb <= "000000";
					when "10001001010000011" => rgb <= "000000";
					when "10001001010000100" => rgb <= "000000";
					when "10001001010000101" => rgb <= "000000";
					when "10001001010000110" => rgb <= "000000";
					when "10001001010000111" => rgb <= "000000";
					when "10001001010001000" => rgb <= "000000";
					when "10001001010001001" => rgb <= "000000";
					when "10001001010001010" => rgb <= "000000";
					when "10001001010001011" => rgb <= "000000";
					when "10001001010001100" => rgb <= "000000";
					when "10001001010001101" => rgb <= "000000";
					when "10001001010001110" => rgb <= "000000";
					when "10001001010001111" => rgb <= "000000";
					when "10001001010010000" => rgb <= "000000";
					when "10001001010010001" => rgb <= "000000";
					when "10001001010010010" => rgb <= "000000";
					when "10001001010010011" => rgb <= "000000";
					when "10001001010010100" => rgb <= "000000";
					when "10001001010010101" => rgb <= "000000";
					when "10001001010010110" => rgb <= "000000";
					when "10001001010010111" => rgb <= "000000";
					when "10001001010011000" => rgb <= "000000";
					when "10001001010011001" => rgb <= "000000";
					when "10001001010011010" => rgb <= "000000";
					when "10001001010011011" => rgb <= "000000";
					when "10001001010011100" => rgb <= "000000";
					when "10001001010011101" => rgb <= "000000";
					when "10001001010011110" => rgb <= "000000";
					when "10001001010011111" => rgb <= "000000";
					when "10001001010100000" => rgb <= "000000";
					when "10001001010100001" => rgb <= "000000";
					when "10001001010100010" => rgb <= "000000";
					when "10001001010100011" => rgb <= "000000";
					when "10001001010100100" => rgb <= "000000";
					when "10001001010100101" => rgb <= "000000";
					when "10001001010100110" => rgb <= "000000";
					when "10001001010100111" => rgb <= "000000";
					when "10001001010101000" => rgb <= "000000";
					when "10001001010101001" => rgb <= "000000";
					when "10001001010101010" => rgb <= "000000";
					when "10001001010101011" => rgb <= "000000";
					when "10001001010101100" => rgb <= "000000";
					when "10001001010101101" => rgb <= "000000";
					when "10001001010101110" => rgb <= "000000";
					when "10001001010101111" => rgb <= "000000";
					when "10001001010110000" => rgb <= "000000";
					when "10001001010110001" => rgb <= "000000";
					when "10001001010110010" => rgb <= "000000";
					when "10001001010110011" => rgb <= "000000";
					when "10001001010110100" => rgb <= "000000";
					when "10001001010110101" => rgb <= "000000";
					when "10001001010110110" => rgb <= "000000";
					when "10001001010110111" => rgb <= "000000";
					when "10001001010111000" => rgb <= "000000";
					when "10001001010111001" => rgb <= "000000";
					when "10001001010111010" => rgb <= "000000";
					when "10001001010111011" => rgb <= "000000";
					when "10001001010111100" => rgb <= "000000";
					when "10001001010111101" => rgb <= "000000";
					when "10001001010111110" => rgb <= "000000";
					when "10001001010111111" => rgb <= "000000";
					when "10001001011000000" => rgb <= "000000";
					when "10001001011000001" => rgb <= "000000";
					when "10001001011000010" => rgb <= "000000";
					when "10001001011000011" => rgb <= "000000";
					when "10001001011000100" => rgb <= "000000";
					when "10001001011000101" => rgb <= "000000";
					when "10001001011000110" => rgb <= "000000";
					when "10001001011000111" => rgb <= "000000";
					when "10001001011001000" => rgb <= "000000";
					when "10001001011001001" => rgb <= "000000";
					when "10001001011001010" => rgb <= "000000";
					when "10001001011001011" => rgb <= "000000";
					when "10001001011001100" => rgb <= "000000";
					when "10001001011001101" => rgb <= "000000";
					when "10001001011001110" => rgb <= "000000";
					when "10001001011001111" => rgb <= "000000";
					when "10001001011010000" => rgb <= "000000";
					when "10001001011010001" => rgb <= "000000";
					when "10001001011010010" => rgb <= "000000";
					when "10001001011010011" => rgb <= "000000";
					when "10001001011010100" => rgb <= "000000";
					when "10001001011010101" => rgb <= "000000";
					when "10001001011010110" => rgb <= "000000";
					when "10001001011010111" => rgb <= "000000";
					when "10001001011011000" => rgb <= "000000";
					when "10001001011011001" => rgb <= "000000";
					when "10001001011011010" => rgb <= "000000";
					when "10001001011011011" => rgb <= "000000";
					when "10001001011011100" => rgb <= "000000";
					when "10001001011011101" => rgb <= "000000";
					when "10001001011011110" => rgb <= "000000";
					when "10001001011011111" => rgb <= "000000";
					when "10001001011100000" => rgb <= "000000";
					when "10001001011100001" => rgb <= "000000";
					when "10001001011100010" => rgb <= "000000";
					when "10001001011100011" => rgb <= "000000";
					when "10001001011100100" => rgb <= "000000";
					when "10001001011100101" => rgb <= "000000";
					when "10001001011100110" => rgb <= "000000";
					when "10001001011100111" => rgb <= "000000";
					when "10001001011101000" => rgb <= "000000";
					when "10001001011101001" => rgb <= "000000";
					when "10001001011101010" => rgb <= "000000";
					when "10001001011101011" => rgb <= "000000";
					when "10001001011101100" => rgb <= "000000";
					when "10001001011101101" => rgb <= "000000";
					when "10001001011101110" => rgb <= "000000";
					when "10001001011101111" => rgb <= "000000";
					when "10001001011110000" => rgb <= "000000";
					when "10001001011110001" => rgb <= "000000";
					when "10001001011110010" => rgb <= "000000";
					when "10001001011110011" => rgb <= "000000";
					when "10001001011110100" => rgb <= "000000";
					when "10001001011110101" => rgb <= "000000";
					when "10001001011110110" => rgb <= "000000";
					when "10001001011110111" => rgb <= "000000";
					when "10001001011111000" => rgb <= "000000";
					when "10001001011111001" => rgb <= "000000";
					when "10001001011111010" => rgb <= "000000";
					when "10001001011111011" => rgb <= "000000";
					when "10001001011111100" => rgb <= "000000";
					when "10001001011111101" => rgb <= "000000";
					when "10001001011111110" => rgb <= "000000";
					when "10001001011111111" => rgb <= "000000";
					when "10001001100000000" => rgb <= "000000";
					when "10001001100000001" => rgb <= "000000";
					when "10001001100000010" => rgb <= "000000";
					when "10001001100000011" => rgb <= "000000";
					when "10001001100000100" => rgb <= "000000";
					when "10001001100000101" => rgb <= "000000";
					when "10001001100000110" => rgb <= "000000";
					when "10001001100000111" => rgb <= "000000";
					when "10001001100001000" => rgb <= "000000";
					when "10001001100001001" => rgb <= "000000";
					when "10001001100001010" => rgb <= "000000";
					when "10001001100001011" => rgb <= "000000";
					when "10001001100001100" => rgb <= "000000";
					when "10001001100001101" => rgb <= "000000";
					when "10001001100001110" => rgb <= "000000";
					when "10001001100001111" => rgb <= "000000";
					when "10001001100010000" => rgb <= "000000";
					when "10001001100010001" => rgb <= "000000";
					when "10001001100010010" => rgb <= "000000";
					when "10001001100010011" => rgb <= "000000";
					when "10001001100010100" => rgb <= "000000";
					when "10001001100010101" => rgb <= "000000";
					when "10001001100010110" => rgb <= "000000";
					when "10001001100010111" => rgb <= "000000";
					when "10001001100011000" => rgb <= "000000";
					when "10001001100011001" => rgb <= "000000";
					when "10001001100011010" => rgb <= "000000";
					when "10001001100011011" => rgb <= "000000";
					when "10001001100011100" => rgb <= "000000";
					when "10001001100011101" => rgb <= "000000";
					when "10001001100011110" => rgb <= "000000";
					when "10001001100011111" => rgb <= "000000";
					when "10001001100100000" => rgb <= "000000";
					when "10001001100100001" => rgb <= "000000";
					when "10001001100100010" => rgb <= "000000";
					when "10001001100100011" => rgb <= "000000";
					when "10001001100100100" => rgb <= "000000";
					when "10001001100100101" => rgb <= "000000";
					when "10001001100100110" => rgb <= "000000";
					when "10001001100100111" => rgb <= "000000";
					when "10001001100101000" => rgb <= "000000";
					when "10001001100101001" => rgb <= "000000";
					when "10001001100101010" => rgb <= "000000";
					when "10001001100101011" => rgb <= "000000";
					when "10001001100101100" => rgb <= "000000";
					when "10001001100101101" => rgb <= "000000";
					when "10001001100101110" => rgb <= "000000";
					when "10001001100101111" => rgb <= "000000";
					when "10001001100110000" => rgb <= "000000";
					when "10001001100110001" => rgb <= "000000";
					when "10001001100110010" => rgb <= "000000";
					when "10001001100110011" => rgb <= "000000";
					when "10001001100110100" => rgb <= "000000";
					when "10001001100110101" => rgb <= "000000";
					when "10001001100110110" => rgb <= "000000";
					when "10001001100110111" => rgb <= "000000";
					when "10001001100111000" => rgb <= "000000";
					when "10001001100111001" => rgb <= "000000";
					when "10001001100111010" => rgb <= "000000";
					when "10001001100111011" => rgb <= "000000";
					when "10001001100111100" => rgb <= "000000";
					when "10001001100111101" => rgb <= "000000";
					when "10001001100111110" => rgb <= "000000";
					when "10001001100111111" => rgb <= "000000";
					when "10001010000000000" => rgb <= "000000";
					when "10001010000000001" => rgb <= "000000";
					when "10001010000000010" => rgb <= "000000";
					when "10001010000000011" => rgb <= "000000";
					when "10001010000000100" => rgb <= "000000";
					when "10001010000000101" => rgb <= "000000";
					when "10001010000000110" => rgb <= "000000";
					when "10001010000000111" => rgb <= "000000";
					when "10001010000001000" => rgb <= "000000";
					when "10001010000001001" => rgb <= "000000";
					when "10001010000001010" => rgb <= "000000";
					when "10001010000001011" => rgb <= "000000";
					when "10001010000001100" => rgb <= "000000";
					when "10001010000001101" => rgb <= "000000";
					when "10001010000001110" => rgb <= "000000";
					when "10001010000001111" => rgb <= "000000";
					when "10001010000010000" => rgb <= "000000";
					when "10001010000010001" => rgb <= "000000";
					when "10001010000010010" => rgb <= "000000";
					when "10001010000010011" => rgb <= "000000";
					when "10001010000010100" => rgb <= "000000";
					when "10001010000010101" => rgb <= "000000";
					when "10001010000010110" => rgb <= "000000";
					when "10001010000010111" => rgb <= "000000";
					when "10001010000011000" => rgb <= "000000";
					when "10001010000011001" => rgb <= "000000";
					when "10001010000011010" => rgb <= "000000";
					when "10001010000011011" => rgb <= "000000";
					when "10001010000011100" => rgb <= "000000";
					when "10001010000011101" => rgb <= "000000";
					when "10001010000011110" => rgb <= "000000";
					when "10001010000011111" => rgb <= "000000";
					when "10001010000100000" => rgb <= "000000";
					when "10001010000100001" => rgb <= "000000";
					when "10001010000100010" => rgb <= "000000";
					when "10001010000100011" => rgb <= "000000";
					when "10001010000100100" => rgb <= "000000";
					when "10001010000100101" => rgb <= "000000";
					when "10001010000100110" => rgb <= "000000";
					when "10001010000100111" => rgb <= "000000";
					when "10001010000101000" => rgb <= "000000";
					when "10001010000101001" => rgb <= "000000";
					when "10001010000101010" => rgb <= "000000";
					when "10001010000101011" => rgb <= "000000";
					when "10001010000101100" => rgb <= "000000";
					when "10001010000101101" => rgb <= "000000";
					when "10001010000101110" => rgb <= "000000";
					when "10001010000101111" => rgb <= "000000";
					when "10001010000110000" => rgb <= "000000";
					when "10001010000110001" => rgb <= "000000";
					when "10001010000110010" => rgb <= "000000";
					when "10001010000110011" => rgb <= "000000";
					when "10001010000110100" => rgb <= "000000";
					when "10001010000110101" => rgb <= "000000";
					when "10001010000110110" => rgb <= "000000";
					when "10001010000110111" => rgb <= "000000";
					when "10001010000111000" => rgb <= "000000";
					when "10001010000111001" => rgb <= "000000";
					when "10001010000111010" => rgb <= "000000";
					when "10001010000111011" => rgb <= "000000";
					when "10001010000111100" => rgb <= "000000";
					when "10001010000111101" => rgb <= "000000";
					when "10001010000111110" => rgb <= "000000";
					when "10001010000111111" => rgb <= "000000";
					when "10001010001000000" => rgb <= "000000";
					when "10001010001000001" => rgb <= "000000";
					when "10001010001000010" => rgb <= "000000";
					when "10001010001000011" => rgb <= "000000";
					when "10001010001000100" => rgb <= "000000";
					when "10001010001000101" => rgb <= "000000";
					when "10001010001000110" => rgb <= "000000";
					when "10001010001000111" => rgb <= "000000";
					when "10001010001001000" => rgb <= "000000";
					when "10001010001001001" => rgb <= "000000";
					when "10001010001001010" => rgb <= "000000";
					when "10001010001001011" => rgb <= "000000";
					when "10001010001001100" => rgb <= "000000";
					when "10001010001001101" => rgb <= "000000";
					when "10001010001001110" => rgb <= "000000";
					when "10001010001001111" => rgb <= "000000";
					when "10001010001010000" => rgb <= "000000";
					when "10001010001010001" => rgb <= "000000";
					when "10001010001010010" => rgb <= "000000";
					when "10001010001010011" => rgb <= "000000";
					when "10001010001010100" => rgb <= "000000";
					when "10001010001010101" => rgb <= "000000";
					when "10001010001010110" => rgb <= "000000";
					when "10001010001010111" => rgb <= "000000";
					when "10001010001011000" => rgb <= "000000";
					when "10001010001011001" => rgb <= "000000";
					when "10001010001011010" => rgb <= "000000";
					when "10001010001011011" => rgb <= "000000";
					when "10001010001011100" => rgb <= "000000";
					when "10001010001011101" => rgb <= "000000";
					when "10001010001011110" => rgb <= "000000";
					when "10001010001011111" => rgb <= "000000";
					when "10001010001100000" => rgb <= "000000";
					when "10001010001100001" => rgb <= "000000";
					when "10001010001100010" => rgb <= "000000";
					when "10001010001100011" => rgb <= "000000";
					when "10001010001100100" => rgb <= "000000";
					when "10001010001100101" => rgb <= "000000";
					when "10001010001100110" => rgb <= "000000";
					when "10001010001100111" => rgb <= "000000";
					when "10001010001101000" => rgb <= "000000";
					when "10001010001101001" => rgb <= "000000";
					when "10001010001101010" => rgb <= "000000";
					when "10001010001101011" => rgb <= "000000";
					when "10001010001101100" => rgb <= "000000";
					when "10001010001101101" => rgb <= "000000";
					when "10001010001101110" => rgb <= "000000";
					when "10001010001101111" => rgb <= "000000";
					when "10001010001110000" => rgb <= "000000";
					when "10001010001110001" => rgb <= "000000";
					when "10001010001110010" => rgb <= "000000";
					when "10001010001110011" => rgb <= "000000";
					when "10001010001110100" => rgb <= "000000";
					when "10001010001110101" => rgb <= "000000";
					when "10001010001110110" => rgb <= "000000";
					when "10001010001110111" => rgb <= "000000";
					when "10001010001111000" => rgb <= "000000";
					when "10001010001111001" => rgb <= "000000";
					when "10001010001111010" => rgb <= "000000";
					when "10001010001111011" => rgb <= "000000";
					when "10001010001111100" => rgb <= "000000";
					when "10001010001111101" => rgb <= "000000";
					when "10001010001111110" => rgb <= "000000";
					when "10001010001111111" => rgb <= "000000";
					when "10001010010000000" => rgb <= "000000";
					when "10001010010000001" => rgb <= "000000";
					when "10001010010000010" => rgb <= "000000";
					when "10001010010000011" => rgb <= "000000";
					when "10001010010000100" => rgb <= "000000";
					when "10001010010000101" => rgb <= "000000";
					when "10001010010000110" => rgb <= "000000";
					when "10001010010000111" => rgb <= "000000";
					when "10001010010001000" => rgb <= "000000";
					when "10001010010001001" => rgb <= "000000";
					when "10001010010001010" => rgb <= "000000";
					when "10001010010001011" => rgb <= "000000";
					when "10001010010001100" => rgb <= "000000";
					when "10001010010001101" => rgb <= "000000";
					when "10001010010001110" => rgb <= "000000";
					when "10001010010001111" => rgb <= "000000";
					when "10001010010010000" => rgb <= "000000";
					when "10001010010010001" => rgb <= "000000";
					when "10001010010010010" => rgb <= "000000";
					when "10001010010010011" => rgb <= "000000";
					when "10001010010010100" => rgb <= "000000";
					when "10001010010010101" => rgb <= "000000";
					when "10001010010010110" => rgb <= "000000";
					when "10001010010010111" => rgb <= "000000";
					when "10001010010011000" => rgb <= "000000";
					when "10001010010011001" => rgb <= "000000";
					when "10001010010011010" => rgb <= "000000";
					when "10001010010011011" => rgb <= "000000";
					when "10001010010011100" => rgb <= "000000";
					when "10001010010011101" => rgb <= "000000";
					when "10001010010011110" => rgb <= "000000";
					when "10001010010011111" => rgb <= "000000";
					when "10001010010100000" => rgb <= "000000";
					when "10001010010100001" => rgb <= "000000";
					when "10001010010100010" => rgb <= "000000";
					when "10001010010100011" => rgb <= "000000";
					when "10001010010100100" => rgb <= "000000";
					when "10001010010100101" => rgb <= "000000";
					when "10001010010100110" => rgb <= "000000";
					when "10001010010100111" => rgb <= "000000";
					when "10001010010101000" => rgb <= "000000";
					when "10001010010101001" => rgb <= "000000";
					when "10001010010101010" => rgb <= "000000";
					when "10001010010101011" => rgb <= "000000";
					when "10001010010101100" => rgb <= "000000";
					when "10001010010101101" => rgb <= "000000";
					when "10001010010101110" => rgb <= "000000";
					when "10001010010101111" => rgb <= "000000";
					when "10001010010110000" => rgb <= "000000";
					when "10001010010110001" => rgb <= "000000";
					when "10001010010110010" => rgb <= "000000";
					when "10001010010110011" => rgb <= "000000";
					when "10001010010110100" => rgb <= "000000";
					when "10001010010110101" => rgb <= "000000";
					when "10001010010110110" => rgb <= "000000";
					when "10001010010110111" => rgb <= "000000";
					when "10001010010111000" => rgb <= "000000";
					when "10001010010111001" => rgb <= "000000";
					when "10001010010111010" => rgb <= "000000";
					when "10001010010111011" => rgb <= "000000";
					when "10001010010111100" => rgb <= "000000";
					when "10001010010111101" => rgb <= "000000";
					when "10001010010111110" => rgb <= "000000";
					when "10001010010111111" => rgb <= "000000";
					when "10001010011000000" => rgb <= "000000";
					when "10001010011000001" => rgb <= "000000";
					when "10001010011000010" => rgb <= "000000";
					when "10001010011000011" => rgb <= "000000";
					when "10001010011000100" => rgb <= "000000";
					when "10001010011000101" => rgb <= "000000";
					when "10001010011000110" => rgb <= "000000";
					when "10001010011000111" => rgb <= "000000";
					when "10001010011001000" => rgb <= "000000";
					when "10001010011001001" => rgb <= "000000";
					when "10001010011001010" => rgb <= "000000";
					when "10001010011001011" => rgb <= "000000";
					when "10001010011001100" => rgb <= "000000";
					when "10001010011001101" => rgb <= "000000";
					when "10001010011001110" => rgb <= "000000";
					when "10001010011001111" => rgb <= "000000";
					when "10001010011010000" => rgb <= "000000";
					when "10001010011010001" => rgb <= "000000";
					when "10001010011010010" => rgb <= "000000";
					when "10001010011010011" => rgb <= "000000";
					when "10001010011010100" => rgb <= "000000";
					when "10001010011010101" => rgb <= "000000";
					when "10001010011010110" => rgb <= "000000";
					when "10001010011010111" => rgb <= "000000";
					when "10001010011011000" => rgb <= "000000";
					when "10001010011011001" => rgb <= "000000";
					when "10001010011011010" => rgb <= "000000";
					when "10001010011011011" => rgb <= "000000";
					when "10001010011011100" => rgb <= "000000";
					when "10001010011011101" => rgb <= "000000";
					when "10001010011011110" => rgb <= "000000";
					when "10001010011011111" => rgb <= "000000";
					when "10001010011100000" => rgb <= "000000";
					when "10001010011100001" => rgb <= "000000";
					when "10001010011100010" => rgb <= "000000";
					when "10001010011100011" => rgb <= "000000";
					when "10001010011100100" => rgb <= "000000";
					when "10001010011100101" => rgb <= "000000";
					when "10001010011100110" => rgb <= "000000";
					when "10001010011100111" => rgb <= "000000";
					when "10001010011101000" => rgb <= "000000";
					when "10001010011101001" => rgb <= "000000";
					when "10001010011101010" => rgb <= "000000";
					when "10001010011101011" => rgb <= "000000";
					when "10001010011101100" => rgb <= "000000";
					when "10001010011101101" => rgb <= "000000";
					when "10001010011101110" => rgb <= "000000";
					when "10001010011101111" => rgb <= "000000";
					when "10001010011110000" => rgb <= "000000";
					when "10001010011110001" => rgb <= "000000";
					when "10001010011110010" => rgb <= "000000";
					when "10001010011110011" => rgb <= "000000";
					when "10001010011110100" => rgb <= "000000";
					when "10001010011110101" => rgb <= "000000";
					when "10001010011110110" => rgb <= "000000";
					when "10001010011110111" => rgb <= "000000";
					when "10001010011111000" => rgb <= "000000";
					when "10001010011111001" => rgb <= "000000";
					when "10001010011111010" => rgb <= "000000";
					when "10001010011111011" => rgb <= "000000";
					when "10001010011111100" => rgb <= "000000";
					when "10001010011111101" => rgb <= "000000";
					when "10001010011111110" => rgb <= "000000";
					when "10001010011111111" => rgb <= "000000";
					when "10001010100000000" => rgb <= "000000";
					when "10001010100000001" => rgb <= "000000";
					when "10001010100000010" => rgb <= "000000";
					when "10001010100000011" => rgb <= "000000";
					when "10001010100000100" => rgb <= "000000";
					when "10001010100000101" => rgb <= "000000";
					when "10001010100000110" => rgb <= "000000";
					when "10001010100000111" => rgb <= "000000";
					when "10001010100001000" => rgb <= "000000";
					when "10001010100001001" => rgb <= "000000";
					when "10001010100001010" => rgb <= "000000";
					when "10001010100001011" => rgb <= "000000";
					when "10001010100001100" => rgb <= "000000";
					when "10001010100001101" => rgb <= "000000";
					when "10001010100001110" => rgb <= "000000";
					when "10001010100001111" => rgb <= "000000";
					when "10001010100010000" => rgb <= "000000";
					when "10001010100010001" => rgb <= "000000";
					when "10001010100010010" => rgb <= "000000";
					when "10001010100010011" => rgb <= "000000";
					when "10001010100010100" => rgb <= "000000";
					when "10001010100010101" => rgb <= "000000";
					when "10001010100010110" => rgb <= "000000";
					when "10001010100010111" => rgb <= "000000";
					when "10001010100011000" => rgb <= "000000";
					when "10001010100011001" => rgb <= "000000";
					when "10001010100011010" => rgb <= "000000";
					when "10001010100011011" => rgb <= "000000";
					when "10001010100011100" => rgb <= "000000";
					when "10001010100011101" => rgb <= "000000";
					when "10001010100011110" => rgb <= "000000";
					when "10001010100011111" => rgb <= "000000";
					when "10001010100100000" => rgb <= "000000";
					when "10001010100100001" => rgb <= "000000";
					when "10001010100100010" => rgb <= "000000";
					when "10001010100100011" => rgb <= "000000";
					when "10001010100100100" => rgb <= "000000";
					when "10001010100100101" => rgb <= "000000";
					when "10001010100100110" => rgb <= "000000";
					when "10001010100100111" => rgb <= "000000";
					when "10001010100101000" => rgb <= "000000";
					when "10001010100101001" => rgb <= "000000";
					when "10001010100101010" => rgb <= "000000";
					when "10001010100101011" => rgb <= "000000";
					when "10001010100101100" => rgb <= "000000";
					when "10001010100101101" => rgb <= "000000";
					when "10001010100101110" => rgb <= "000000";
					when "10001010100101111" => rgb <= "000000";
					when "10001010100110000" => rgb <= "000000";
					when "10001010100110001" => rgb <= "000000";
					when "10001010100110010" => rgb <= "000000";
					when "10001010100110011" => rgb <= "000000";
					when "10001010100110100" => rgb <= "000000";
					when "10001010100110101" => rgb <= "000000";
					when "10001010100110110" => rgb <= "000000";
					when "10001010100110111" => rgb <= "000000";
					when "10001010100111000" => rgb <= "000000";
					when "10001010100111001" => rgb <= "000000";
					when "10001010100111010" => rgb <= "000000";
					when "10001010100111011" => rgb <= "000000";
					when "10001010100111100" => rgb <= "000000";
					when "10001010100111101" => rgb <= "000000";
					when "10001010100111110" => rgb <= "000000";
					when "10001010100111111" => rgb <= "000000";
					when "10001011000000000" => rgb <= "000000";
					when "10001011000000001" => rgb <= "000000";
					when "10001011000000010" => rgb <= "000000";
					when "10001011000000011" => rgb <= "000000";
					when "10001011000000100" => rgb <= "000000";
					when "10001011000000101" => rgb <= "000000";
					when "10001011000000110" => rgb <= "000000";
					when "10001011000000111" => rgb <= "000000";
					when "10001011000001000" => rgb <= "000000";
					when "10001011000001001" => rgb <= "000000";
					when "10001011000001010" => rgb <= "000000";
					when "10001011000001011" => rgb <= "000000";
					when "10001011000001100" => rgb <= "000000";
					when "10001011000001101" => rgb <= "000000";
					when "10001011000001110" => rgb <= "000000";
					when "10001011000001111" => rgb <= "000000";
					when "10001011000010000" => rgb <= "000000";
					when "10001011000010001" => rgb <= "000000";
					when "10001011000010010" => rgb <= "000000";
					when "10001011000010011" => rgb <= "000000";
					when "10001011000010100" => rgb <= "000000";
					when "10001011000010101" => rgb <= "000000";
					when "10001011000010110" => rgb <= "000000";
					when "10001011000010111" => rgb <= "000000";
					when "10001011000011000" => rgb <= "000000";
					when "10001011000011001" => rgb <= "000000";
					when "10001011000011010" => rgb <= "000000";
					when "10001011000011011" => rgb <= "000000";
					when "10001011000011100" => rgb <= "000000";
					when "10001011000011101" => rgb <= "000000";
					when "10001011000011110" => rgb <= "000000";
					when "10001011000011111" => rgb <= "000000";
					when "10001011000100000" => rgb <= "000000";
					when "10001011000100001" => rgb <= "000000";
					when "10001011000100010" => rgb <= "000000";
					when "10001011000100011" => rgb <= "000000";
					when "10001011000100100" => rgb <= "000000";
					when "10001011000100101" => rgb <= "000000";
					when "10001011000100110" => rgb <= "000000";
					when "10001011000100111" => rgb <= "000000";
					when "10001011000101000" => rgb <= "000000";
					when "10001011000101001" => rgb <= "000000";
					when "10001011000101010" => rgb <= "000000";
					when "10001011000101011" => rgb <= "000000";
					when "10001011000101100" => rgb <= "000000";
					when "10001011000101101" => rgb <= "000000";
					when "10001011000101110" => rgb <= "000000";
					when "10001011000101111" => rgb <= "000000";
					when "10001011000110000" => rgb <= "000000";
					when "10001011000110001" => rgb <= "000000";
					when "10001011000110010" => rgb <= "000000";
					when "10001011000110011" => rgb <= "000000";
					when "10001011000110100" => rgb <= "000000";
					when "10001011000110101" => rgb <= "000000";
					when "10001011000110110" => rgb <= "000000";
					when "10001011000110111" => rgb <= "000000";
					when "10001011000111000" => rgb <= "000000";
					when "10001011000111001" => rgb <= "000000";
					when "10001011000111010" => rgb <= "000000";
					when "10001011000111011" => rgb <= "000000";
					when "10001011000111100" => rgb <= "000000";
					when "10001011000111101" => rgb <= "000000";
					when "10001011000111110" => rgb <= "000000";
					when "10001011000111111" => rgb <= "000000";
					when "10001011001000000" => rgb <= "000000";
					when "10001011001000001" => rgb <= "000000";
					when "10001011001000010" => rgb <= "000000";
					when "10001011001000011" => rgb <= "000000";
					when "10001011001000100" => rgb <= "000000";
					when "10001011001000101" => rgb <= "000000";
					when "10001011001000110" => rgb <= "000000";
					when "10001011001000111" => rgb <= "000000";
					when "10001011001001000" => rgb <= "000000";
					when "10001011001001001" => rgb <= "000000";
					when "10001011001001010" => rgb <= "000000";
					when "10001011001001011" => rgb <= "000000";
					when "10001011001001100" => rgb <= "000000";
					when "10001011001001101" => rgb <= "000000";
					when "10001011001001110" => rgb <= "000000";
					when "10001011001001111" => rgb <= "000000";
					when "10001011001010000" => rgb <= "000000";
					when "10001011001010001" => rgb <= "000000";
					when "10001011001010010" => rgb <= "000000";
					when "10001011001010011" => rgb <= "000000";
					when "10001011001010100" => rgb <= "000000";
					when "10001011001010101" => rgb <= "000000";
					when "10001011001010110" => rgb <= "000000";
					when "10001011001010111" => rgb <= "000000";
					when "10001011001011000" => rgb <= "000000";
					when "10001011001011001" => rgb <= "000000";
					when "10001011001011010" => rgb <= "000000";
					when "10001011001011011" => rgb <= "000000";
					when "10001011001011100" => rgb <= "000000";
					when "10001011001011101" => rgb <= "000000";
					when "10001011001011110" => rgb <= "000000";
					when "10001011001011111" => rgb <= "000000";
					when "10001011001100000" => rgb <= "000000";
					when "10001011001100001" => rgb <= "000000";
					when "10001011001100010" => rgb <= "000000";
					when "10001011001100011" => rgb <= "000000";
					when "10001011001100100" => rgb <= "000000";
					when "10001011001100101" => rgb <= "000000";
					when "10001011001100110" => rgb <= "000000";
					when "10001011001100111" => rgb <= "000000";
					when "10001011001101000" => rgb <= "000000";
					when "10001011001101001" => rgb <= "000000";
					when "10001011001101010" => rgb <= "000000";
					when "10001011001101011" => rgb <= "000000";
					when "10001011001101100" => rgb <= "000000";
					when "10001011001101101" => rgb <= "000000";
					when "10001011001101110" => rgb <= "000000";
					when "10001011001101111" => rgb <= "000000";
					when "10001011001110000" => rgb <= "000000";
					when "10001011001110001" => rgb <= "000000";
					when "10001011001110010" => rgb <= "000000";
					when "10001011001110011" => rgb <= "000000";
					when "10001011001110100" => rgb <= "000000";
					when "10001011001110101" => rgb <= "000000";
					when "10001011001110110" => rgb <= "000000";
					when "10001011001110111" => rgb <= "000000";
					when "10001011001111000" => rgb <= "000000";
					when "10001011001111001" => rgb <= "000000";
					when "10001011001111010" => rgb <= "000000";
					when "10001011001111011" => rgb <= "000000";
					when "10001011001111100" => rgb <= "000000";
					when "10001011001111101" => rgb <= "000000";
					when "10001011001111110" => rgb <= "000000";
					when "10001011001111111" => rgb <= "000000";
					when "10001011010000000" => rgb <= "000000";
					when "10001011010000001" => rgb <= "000000";
					when "10001011010000010" => rgb <= "000000";
					when "10001011010000011" => rgb <= "000000";
					when "10001011010000100" => rgb <= "000000";
					when "10001011010000101" => rgb <= "000000";
					when "10001011010000110" => rgb <= "000000";
					when "10001011010000111" => rgb <= "000000";
					when "10001011010001000" => rgb <= "000000";
					when "10001011010001001" => rgb <= "000000";
					when "10001011010001010" => rgb <= "000000";
					when "10001011010001011" => rgb <= "000000";
					when "10001011010001100" => rgb <= "000000";
					when "10001011010001101" => rgb <= "000000";
					when "10001011010001110" => rgb <= "000000";
					when "10001011010001111" => rgb <= "000000";
					when "10001011010010000" => rgb <= "000000";
					when "10001011010010001" => rgb <= "000000";
					when "10001011010010010" => rgb <= "000000";
					when "10001011010010011" => rgb <= "000000";
					when "10001011010010100" => rgb <= "000000";
					when "10001011010010101" => rgb <= "000000";
					when "10001011010010110" => rgb <= "000000";
					when "10001011010010111" => rgb <= "000000";
					when "10001011010011000" => rgb <= "000000";
					when "10001011010011001" => rgb <= "000000";
					when "10001011010011010" => rgb <= "000000";
					when "10001011010011011" => rgb <= "000000";
					when "10001011010011100" => rgb <= "000000";
					when "10001011010011101" => rgb <= "000000";
					when "10001011010011110" => rgb <= "000000";
					when "10001011010011111" => rgb <= "000000";
					when "10001011010100000" => rgb <= "000000";
					when "10001011010100001" => rgb <= "000000";
					when "10001011010100010" => rgb <= "000000";
					when "10001011010100011" => rgb <= "000000";
					when "10001011010100100" => rgb <= "000000";
					when "10001011010100101" => rgb <= "000000";
					when "10001011010100110" => rgb <= "000000";
					when "10001011010100111" => rgb <= "000000";
					when "10001011010101000" => rgb <= "000000";
					when "10001011010101001" => rgb <= "000000";
					when "10001011010101010" => rgb <= "000000";
					when "10001011010101011" => rgb <= "000000";
					when "10001011010101100" => rgb <= "000000";
					when "10001011010101101" => rgb <= "000000";
					when "10001011010101110" => rgb <= "000000";
					when "10001011010101111" => rgb <= "000000";
					when "10001011010110000" => rgb <= "000000";
					when "10001011010110001" => rgb <= "000000";
					when "10001011010110010" => rgb <= "000000";
					when "10001011010110011" => rgb <= "000000";
					when "10001011010110100" => rgb <= "000000";
					when "10001011010110101" => rgb <= "000000";
					when "10001011010110110" => rgb <= "000000";
					when "10001011010110111" => rgb <= "000000";
					when "10001011010111000" => rgb <= "000000";
					when "10001011010111001" => rgb <= "000000";
					when "10001011010111010" => rgb <= "000000";
					when "10001011010111011" => rgb <= "000000";
					when "10001011010111100" => rgb <= "000000";
					when "10001011010111101" => rgb <= "000000";
					when "10001011010111110" => rgb <= "000000";
					when "10001011010111111" => rgb <= "000000";
					when "10001011011000000" => rgb <= "000000";
					when "10001011011000001" => rgb <= "000000";
					when "10001011011000010" => rgb <= "000000";
					when "10001011011000011" => rgb <= "000000";
					when "10001011011000100" => rgb <= "000000";
					when "10001011011000101" => rgb <= "000000";
					when "10001011011000110" => rgb <= "000000";
					when "10001011011000111" => rgb <= "000000";
					when "10001011011001000" => rgb <= "000000";
					when "10001011011001001" => rgb <= "000000";
					when "10001011011001010" => rgb <= "000000";
					when "10001011011001011" => rgb <= "000000";
					when "10001011011001100" => rgb <= "000000";
					when "10001011011001101" => rgb <= "000000";
					when "10001011011001110" => rgb <= "000000";
					when "10001011011001111" => rgb <= "000000";
					when "10001011011010000" => rgb <= "000000";
					when "10001011011010001" => rgb <= "000000";
					when "10001011011010010" => rgb <= "000000";
					when "10001011011010011" => rgb <= "000000";
					when "10001011011010100" => rgb <= "000000";
					when "10001011011010101" => rgb <= "000000";
					when "10001011011010110" => rgb <= "000000";
					when "10001011011010111" => rgb <= "000000";
					when "10001011011011000" => rgb <= "000000";
					when "10001011011011001" => rgb <= "000000";
					when "10001011011011010" => rgb <= "000000";
					when "10001011011011011" => rgb <= "000000";
					when "10001011011011100" => rgb <= "000000";
					when "10001011011011101" => rgb <= "000000";
					when "10001011011011110" => rgb <= "000000";
					when "10001011011011111" => rgb <= "000000";
					when "10001011011100000" => rgb <= "000000";
					when "10001011011100001" => rgb <= "000000";
					when "10001011011100010" => rgb <= "000000";
					when "10001011011100011" => rgb <= "000000";
					when "10001011011100100" => rgb <= "000000";
					when "10001011011100101" => rgb <= "000000";
					when "10001011011100110" => rgb <= "000000";
					when "10001011011100111" => rgb <= "000000";
					when "10001011011101000" => rgb <= "000000";
					when "10001011011101001" => rgb <= "000000";
					when "10001011011101010" => rgb <= "000000";
					when "10001011011101011" => rgb <= "000000";
					when "10001011011101100" => rgb <= "000000";
					when "10001011011101101" => rgb <= "000000";
					when "10001011011101110" => rgb <= "000000";
					when "10001011011101111" => rgb <= "000000";
					when "10001011011110000" => rgb <= "000000";
					when "10001011011110001" => rgb <= "000000";
					when "10001011011110010" => rgb <= "000000";
					when "10001011011110011" => rgb <= "000000";
					when "10001011011110100" => rgb <= "000000";
					when "10001011011110101" => rgb <= "000000";
					when "10001011011110110" => rgb <= "000000";
					when "10001011011110111" => rgb <= "000000";
					when "10001011011111000" => rgb <= "000000";
					when "10001011011111001" => rgb <= "000000";
					when "10001011011111010" => rgb <= "000000";
					when "10001011011111011" => rgb <= "000000";
					when "10001011011111100" => rgb <= "000000";
					when "10001011011111101" => rgb <= "000000";
					when "10001011011111110" => rgb <= "000000";
					when "10001011011111111" => rgb <= "000000";
					when "10001011100000000" => rgb <= "000000";
					when "10001011100000001" => rgb <= "000000";
					when "10001011100000010" => rgb <= "000000";
					when "10001011100000011" => rgb <= "000000";
					when "10001011100000100" => rgb <= "000000";
					when "10001011100000101" => rgb <= "000000";
					when "10001011100000110" => rgb <= "000000";
					when "10001011100000111" => rgb <= "000000";
					when "10001011100001000" => rgb <= "000000";
					when "10001011100001001" => rgb <= "000000";
					when "10001011100001010" => rgb <= "000000";
					when "10001011100001011" => rgb <= "000000";
					when "10001011100001100" => rgb <= "000000";
					when "10001011100001101" => rgb <= "000000";
					when "10001011100001110" => rgb <= "000000";
					when "10001011100001111" => rgb <= "000000";
					when "10001011100010000" => rgb <= "000000";
					when "10001011100010001" => rgb <= "000000";
					when "10001011100010010" => rgb <= "000000";
					when "10001011100010011" => rgb <= "000000";
					when "10001011100010100" => rgb <= "000000";
					when "10001011100010101" => rgb <= "000000";
					when "10001011100010110" => rgb <= "000000";
					when "10001011100010111" => rgb <= "000000";
					when "10001011100011000" => rgb <= "000000";
					when "10001011100011001" => rgb <= "000000";
					when "10001011100011010" => rgb <= "000000";
					when "10001011100011011" => rgb <= "000000";
					when "10001011100011100" => rgb <= "000000";
					when "10001011100011101" => rgb <= "000000";
					when "10001011100011110" => rgb <= "000000";
					when "10001011100011111" => rgb <= "000000";
					when "10001011100100000" => rgb <= "000000";
					when "10001011100100001" => rgb <= "000000";
					when "10001011100100010" => rgb <= "000000";
					when "10001011100100011" => rgb <= "000000";
					when "10001011100100100" => rgb <= "000000";
					when "10001011100100101" => rgb <= "000000";
					when "10001011100100110" => rgb <= "000000";
					when "10001011100100111" => rgb <= "000000";
					when "10001011100101000" => rgb <= "000000";
					when "10001011100101001" => rgb <= "000000";
					when "10001011100101010" => rgb <= "000000";
					when "10001011100101011" => rgb <= "000000";
					when "10001011100101100" => rgb <= "000000";
					when "10001011100101101" => rgb <= "000000";
					when "10001011100101110" => rgb <= "000000";
					when "10001011100101111" => rgb <= "000000";
					when "10001011100110000" => rgb <= "000000";
					when "10001011100110001" => rgb <= "000000";
					when "10001011100110010" => rgb <= "000000";
					when "10001011100110011" => rgb <= "000000";
					when "10001011100110100" => rgb <= "000000";
					when "10001011100110101" => rgb <= "000000";
					when "10001011100110110" => rgb <= "000000";
					when "10001011100110111" => rgb <= "000000";
					when "10001011100111000" => rgb <= "000000";
					when "10001011100111001" => rgb <= "000000";
					when "10001011100111010" => rgb <= "000000";
					when "10001011100111011" => rgb <= "000000";
					when "10001011100111100" => rgb <= "000000";
					when "10001011100111101" => rgb <= "000000";
					when "10001011100111110" => rgb <= "000000";
					when "10001011100111111" => rgb <= "000000";
					when "10001100000000000" => rgb <= "000000";
					when "10001100000000001" => rgb <= "000000";
					when "10001100000000010" => rgb <= "000000";
					when "10001100000000011" => rgb <= "000000";
					when "10001100000000100" => rgb <= "000000";
					when "10001100000000101" => rgb <= "000000";
					when "10001100000000110" => rgb <= "000000";
					when "10001100000000111" => rgb <= "000000";
					when "10001100000001000" => rgb <= "000000";
					when "10001100000001001" => rgb <= "000000";
					when "10001100000001010" => rgb <= "000000";
					when "10001100000001011" => rgb <= "000000";
					when "10001100000001100" => rgb <= "000000";
					when "10001100000001101" => rgb <= "000000";
					when "10001100000001110" => rgb <= "000000";
					when "10001100000001111" => rgb <= "000000";
					when "10001100000010000" => rgb <= "000000";
					when "10001100000010001" => rgb <= "000000";
					when "10001100000010010" => rgb <= "000000";
					when "10001100000010011" => rgb <= "000000";
					when "10001100000010100" => rgb <= "000000";
					when "10001100000010101" => rgb <= "000000";
					when "10001100000010110" => rgb <= "000000";
					when "10001100000010111" => rgb <= "000000";
					when "10001100000011000" => rgb <= "000000";
					when "10001100000011001" => rgb <= "000000";
					when "10001100000011010" => rgb <= "000000";
					when "10001100000011011" => rgb <= "000000";
					when "10001100000011100" => rgb <= "000000";
					when "10001100000011101" => rgb <= "000000";
					when "10001100000011110" => rgb <= "000000";
					when "10001100000011111" => rgb <= "000000";
					when "10001100000100000" => rgb <= "000000";
					when "10001100000100001" => rgb <= "000000";
					when "10001100000100010" => rgb <= "000000";
					when "10001100000100011" => rgb <= "000000";
					when "10001100000100100" => rgb <= "000000";
					when "10001100000100101" => rgb <= "000000";
					when "10001100000100110" => rgb <= "000000";
					when "10001100000100111" => rgb <= "000000";
					when "10001100000101000" => rgb <= "000000";
					when "10001100000101001" => rgb <= "000000";
					when "10001100000101010" => rgb <= "000000";
					when "10001100000101011" => rgb <= "000000";
					when "10001100000101100" => rgb <= "000000";
					when "10001100000101101" => rgb <= "000000";
					when "10001100000101110" => rgb <= "000000";
					when "10001100000101111" => rgb <= "000000";
					when "10001100000110000" => rgb <= "000000";
					when "10001100000110001" => rgb <= "000000";
					when "10001100000110010" => rgb <= "000000";
					when "10001100000110011" => rgb <= "000000";
					when "10001100000110100" => rgb <= "000000";
					when "10001100000110101" => rgb <= "000000";
					when "10001100000110110" => rgb <= "000000";
					when "10001100000110111" => rgb <= "000000";
					when "10001100000111000" => rgb <= "000000";
					when "10001100000111001" => rgb <= "000000";
					when "10001100000111010" => rgb <= "000000";
					when "10001100000111011" => rgb <= "000000";
					when "10001100000111100" => rgb <= "000000";
					when "10001100000111101" => rgb <= "000000";
					when "10001100000111110" => rgb <= "000000";
					when "10001100000111111" => rgb <= "000000";
					when "10001100001000000" => rgb <= "000000";
					when "10001100001000001" => rgb <= "000000";
					when "10001100001000010" => rgb <= "000000";
					when "10001100001000011" => rgb <= "000000";
					when "10001100001000100" => rgb <= "000000";
					when "10001100001000101" => rgb <= "000000";
					when "10001100001000110" => rgb <= "000000";
					when "10001100001000111" => rgb <= "000000";
					when "10001100001001000" => rgb <= "000000";
					when "10001100001001001" => rgb <= "000000";
					when "10001100001001010" => rgb <= "000000";
					when "10001100001001011" => rgb <= "000000";
					when "10001100001001100" => rgb <= "000000";
					when "10001100001001101" => rgb <= "000000";
					when "10001100001001110" => rgb <= "000000";
					when "10001100001001111" => rgb <= "000000";
					when "10001100001010000" => rgb <= "000000";
					when "10001100001010001" => rgb <= "000000";
					when "10001100001010010" => rgb <= "000000";
					when "10001100001010011" => rgb <= "000000";
					when "10001100001010100" => rgb <= "000000";
					when "10001100001010101" => rgb <= "000000";
					when "10001100001010110" => rgb <= "000000";
					when "10001100001010111" => rgb <= "000000";
					when "10001100001011000" => rgb <= "000000";
					when "10001100001011001" => rgb <= "000000";
					when "10001100001011010" => rgb <= "000000";
					when "10001100001011011" => rgb <= "000000";
					when "10001100001011100" => rgb <= "000000";
					when "10001100001011101" => rgb <= "000000";
					when "10001100001011110" => rgb <= "000000";
					when "10001100001011111" => rgb <= "000000";
					when "10001100001100000" => rgb <= "000000";
					when "10001100001100001" => rgb <= "000000";
					when "10001100001100010" => rgb <= "000000";
					when "10001100001100011" => rgb <= "000000";
					when "10001100001100100" => rgb <= "000000";
					when "10001100001100101" => rgb <= "000000";
					when "10001100001100110" => rgb <= "000000";
					when "10001100001100111" => rgb <= "000000";
					when "10001100001101000" => rgb <= "000000";
					when "10001100001101001" => rgb <= "000000";
					when "10001100001101010" => rgb <= "000000";
					when "10001100001101011" => rgb <= "000000";
					when "10001100001101100" => rgb <= "000000";
					when "10001100001101101" => rgb <= "000000";
					when "10001100001101110" => rgb <= "000000";
					when "10001100001101111" => rgb <= "000000";
					when "10001100001110000" => rgb <= "000000";
					when "10001100001110001" => rgb <= "000000";
					when "10001100001110010" => rgb <= "000000";
					when "10001100001110011" => rgb <= "000000";
					when "10001100001110100" => rgb <= "000000";
					when "10001100001110101" => rgb <= "000000";
					when "10001100001110110" => rgb <= "000000";
					when "10001100001110111" => rgb <= "000000";
					when "10001100001111000" => rgb <= "000000";
					when "10001100001111001" => rgb <= "000000";
					when "10001100001111010" => rgb <= "000000";
					when "10001100001111011" => rgb <= "000000";
					when "10001100001111100" => rgb <= "000000";
					when "10001100001111101" => rgb <= "000000";
					when "10001100001111110" => rgb <= "000000";
					when "10001100001111111" => rgb <= "000000";
					when "10001100010000000" => rgb <= "000000";
					when "10001100010000001" => rgb <= "000000";
					when "10001100010000010" => rgb <= "000000";
					when "10001100010000011" => rgb <= "000000";
					when "10001100010000100" => rgb <= "000000";
					when "10001100010000101" => rgb <= "000000";
					when "10001100010000110" => rgb <= "000000";
					when "10001100010000111" => rgb <= "000000";
					when "10001100010001000" => rgb <= "000000";
					when "10001100010001001" => rgb <= "000000";
					when "10001100010001010" => rgb <= "000000";
					when "10001100010001011" => rgb <= "000000";
					when "10001100010001100" => rgb <= "000000";
					when "10001100010001101" => rgb <= "000000";
					when "10001100010001110" => rgb <= "000000";
					when "10001100010001111" => rgb <= "000000";
					when "10001100010010000" => rgb <= "000000";
					when "10001100010010001" => rgb <= "000000";
					when "10001100010010010" => rgb <= "000000";
					when "10001100010010011" => rgb <= "000000";
					when "10001100010010100" => rgb <= "000000";
					when "10001100010010101" => rgb <= "000000";
					when "10001100010010110" => rgb <= "000000";
					when "10001100010010111" => rgb <= "000000";
					when "10001100010011000" => rgb <= "000000";
					when "10001100010011001" => rgb <= "000000";
					when "10001100010011010" => rgb <= "000000";
					when "10001100010011011" => rgb <= "000000";
					when "10001100010011100" => rgb <= "000000";
					when "10001100010011101" => rgb <= "000000";
					when "10001100010011110" => rgb <= "000000";
					when "10001100010011111" => rgb <= "000000";
					when "10001100010100000" => rgb <= "000000";
					when "10001100010100001" => rgb <= "000000";
					when "10001100010100010" => rgb <= "000000";
					when "10001100010100011" => rgb <= "000000";
					when "10001100010100100" => rgb <= "000000";
					when "10001100010100101" => rgb <= "000000";
					when "10001100010100110" => rgb <= "000000";
					when "10001100010100111" => rgb <= "000000";
					when "10001100010101000" => rgb <= "000000";
					when "10001100010101001" => rgb <= "000000";
					when "10001100010101010" => rgb <= "000000";
					when "10001100010101011" => rgb <= "000000";
					when "10001100010101100" => rgb <= "000000";
					when "10001100010101101" => rgb <= "000000";
					when "10001100010101110" => rgb <= "000000";
					when "10001100010101111" => rgb <= "000000";
					when "10001100010110000" => rgb <= "000000";
					when "10001100010110001" => rgb <= "000000";
					when "10001100010110010" => rgb <= "000000";
					when "10001100010110011" => rgb <= "000000";
					when "10001100010110100" => rgb <= "000000";
					when "10001100010110101" => rgb <= "000000";
					when "10001100010110110" => rgb <= "000000";
					when "10001100010110111" => rgb <= "000000";
					when "10001100010111000" => rgb <= "000000";
					when "10001100010111001" => rgb <= "000000";
					when "10001100010111010" => rgb <= "000000";
					when "10001100010111011" => rgb <= "000000";
					when "10001100010111100" => rgb <= "000000";
					when "10001100010111101" => rgb <= "000000";
					when "10001100010111110" => rgb <= "000000";
					when "10001100010111111" => rgb <= "000000";
					when "10001100011000000" => rgb <= "000000";
					when "10001100011000001" => rgb <= "000000";
					when "10001100011000010" => rgb <= "000000";
					when "10001100011000011" => rgb <= "000000";
					when "10001100011000100" => rgb <= "000000";
					when "10001100011000101" => rgb <= "000000";
					when "10001100011000110" => rgb <= "000000";
					when "10001100011000111" => rgb <= "000000";
					when "10001100011001000" => rgb <= "000000";
					when "10001100011001001" => rgb <= "000000";
					when "10001100011001010" => rgb <= "000000";
					when "10001100011001011" => rgb <= "000000";
					when "10001100011001100" => rgb <= "000000";
					when "10001100011001101" => rgb <= "000000";
					when "10001100011001110" => rgb <= "000000";
					when "10001100011001111" => rgb <= "000000";
					when "10001100011010000" => rgb <= "000000";
					when "10001100011010001" => rgb <= "000000";
					when "10001100011010010" => rgb <= "000000";
					when "10001100011010011" => rgb <= "000000";
					when "10001100011010100" => rgb <= "000000";
					when "10001100011010101" => rgb <= "000000";
					when "10001100011010110" => rgb <= "000000";
					when "10001100011010111" => rgb <= "000000";
					when "10001100011011000" => rgb <= "000000";
					when "10001100011011001" => rgb <= "000000";
					when "10001100011011010" => rgb <= "000000";
					when "10001100011011011" => rgb <= "000000";
					when "10001100011011100" => rgb <= "000000";
					when "10001100011011101" => rgb <= "000000";
					when "10001100011011110" => rgb <= "000000";
					when "10001100011011111" => rgb <= "000000";
					when "10001100011100000" => rgb <= "000000";
					when "10001100011100001" => rgb <= "000000";
					when "10001100011100010" => rgb <= "000000";
					when "10001100011100011" => rgb <= "000000";
					when "10001100011100100" => rgb <= "000000";
					when "10001100011100101" => rgb <= "000000";
					when "10001100011100110" => rgb <= "000000";
					when "10001100011100111" => rgb <= "000000";
					when "10001100011101000" => rgb <= "000000";
					when "10001100011101001" => rgb <= "000000";
					when "10001100011101010" => rgb <= "000000";
					when "10001100011101011" => rgb <= "000000";
					when "10001100011101100" => rgb <= "000000";
					when "10001100011101101" => rgb <= "000000";
					when "10001100011101110" => rgb <= "000000";
					when "10001100011101111" => rgb <= "000000";
					when "10001100011110000" => rgb <= "000000";
					when "10001100011110001" => rgb <= "000000";
					when "10001100011110010" => rgb <= "000000";
					when "10001100011110011" => rgb <= "000000";
					when "10001100011110100" => rgb <= "000000";
					when "10001100011110101" => rgb <= "000000";
					when "10001100011110110" => rgb <= "000000";
					when "10001100011110111" => rgb <= "000000";
					when "10001100011111000" => rgb <= "000000";
					when "10001100011111001" => rgb <= "000000";
					when "10001100011111010" => rgb <= "000000";
					when "10001100011111011" => rgb <= "000000";
					when "10001100011111100" => rgb <= "000000";
					when "10001100011111101" => rgb <= "000000";
					when "10001100011111110" => rgb <= "000000";
					when "10001100011111111" => rgb <= "000000";
					when "10001100100000000" => rgb <= "000000";
					when "10001100100000001" => rgb <= "000000";
					when "10001100100000010" => rgb <= "000000";
					when "10001100100000011" => rgb <= "000000";
					when "10001100100000100" => rgb <= "000000";
					when "10001100100000101" => rgb <= "000000";
					when "10001100100000110" => rgb <= "000000";
					when "10001100100000111" => rgb <= "000000";
					when "10001100100001000" => rgb <= "000000";
					when "10001100100001001" => rgb <= "000000";
					when "10001100100001010" => rgb <= "000000";
					when "10001100100001011" => rgb <= "000000";
					when "10001100100001100" => rgb <= "000000";
					when "10001100100001101" => rgb <= "000000";
					when "10001100100001110" => rgb <= "000000";
					when "10001100100001111" => rgb <= "000000";
					when "10001100100010000" => rgb <= "000000";
					when "10001100100010001" => rgb <= "000000";
					when "10001100100010010" => rgb <= "000000";
					when "10001100100010011" => rgb <= "000000";
					when "10001100100010100" => rgb <= "000000";
					when "10001100100010101" => rgb <= "000000";
					when "10001100100010110" => rgb <= "000000";
					when "10001100100010111" => rgb <= "000000";
					when "10001100100011000" => rgb <= "000000";
					when "10001100100011001" => rgb <= "000000";
					when "10001100100011010" => rgb <= "000000";
					when "10001100100011011" => rgb <= "000000";
					when "10001100100011100" => rgb <= "000000";
					when "10001100100011101" => rgb <= "000000";
					when "10001100100011110" => rgb <= "000000";
					when "10001100100011111" => rgb <= "000000";
					when "10001100100100000" => rgb <= "000000";
					when "10001100100100001" => rgb <= "000000";
					when "10001100100100010" => rgb <= "000000";
					when "10001100100100011" => rgb <= "000000";
					when "10001100100100100" => rgb <= "000000";
					when "10001100100100101" => rgb <= "000000";
					when "10001100100100110" => rgb <= "000000";
					when "10001100100100111" => rgb <= "000000";
					when "10001100100101000" => rgb <= "000000";
					when "10001100100101001" => rgb <= "000000";
					when "10001100100101010" => rgb <= "000000";
					when "10001100100101011" => rgb <= "000000";
					when "10001100100101100" => rgb <= "000000";
					when "10001100100101101" => rgb <= "000000";
					when "10001100100101110" => rgb <= "000000";
					when "10001100100101111" => rgb <= "000000";
					when "10001100100110000" => rgb <= "000000";
					when "10001100100110001" => rgb <= "000000";
					when "10001100100110010" => rgb <= "000000";
					when "10001100100110011" => rgb <= "000000";
					when "10001100100110100" => rgb <= "000000";
					when "10001100100110101" => rgb <= "000000";
					when "10001100100110110" => rgb <= "000000";
					when "10001100100110111" => rgb <= "000000";
					when "10001100100111000" => rgb <= "000000";
					when "10001100100111001" => rgb <= "000000";
					when "10001100100111010" => rgb <= "000000";
					when "10001100100111011" => rgb <= "000000";
					when "10001100100111100" => rgb <= "000000";
					when "10001100100111101" => rgb <= "000000";
					when "10001100100111110" => rgb <= "000000";
					when "10001100100111111" => rgb <= "000000";
					when "10001101000000000" => rgb <= "000000";
					when "10001101000000001" => rgb <= "000000";
					when "10001101000000010" => rgb <= "000000";
					when "10001101000000011" => rgb <= "000000";
					when "10001101000000100" => rgb <= "000000";
					when "10001101000000101" => rgb <= "000000";
					when "10001101000000110" => rgb <= "000000";
					when "10001101000000111" => rgb <= "000000";
					when "10001101000001000" => rgb <= "000000";
					when "10001101000001001" => rgb <= "000000";
					when "10001101000001010" => rgb <= "000000";
					when "10001101000001011" => rgb <= "000000";
					when "10001101000001100" => rgb <= "000000";
					when "10001101000001101" => rgb <= "000000";
					when "10001101000001110" => rgb <= "000000";
					when "10001101000001111" => rgb <= "000000";
					when "10001101000010000" => rgb <= "000000";
					when "10001101000010001" => rgb <= "000000";
					when "10001101000010010" => rgb <= "000000";
					when "10001101000010011" => rgb <= "000000";
					when "10001101000010100" => rgb <= "000000";
					when "10001101000010101" => rgb <= "000000";
					when "10001101000010110" => rgb <= "000000";
					when "10001101000010111" => rgb <= "000000";
					when "10001101000011000" => rgb <= "000000";
					when "10001101000011001" => rgb <= "000000";
					when "10001101000011010" => rgb <= "000000";
					when "10001101000011011" => rgb <= "000000";
					when "10001101000011100" => rgb <= "000000";
					when "10001101000011101" => rgb <= "000000";
					when "10001101000011110" => rgb <= "000000";
					when "10001101000011111" => rgb <= "000000";
					when "10001101000100000" => rgb <= "000000";
					when "10001101000100001" => rgb <= "000000";
					when "10001101000100010" => rgb <= "000000";
					when "10001101000100011" => rgb <= "000000";
					when "10001101000100100" => rgb <= "000000";
					when "10001101000100101" => rgb <= "000000";
					when "10001101000100110" => rgb <= "000000";
					when "10001101000100111" => rgb <= "000000";
					when "10001101000101000" => rgb <= "000000";
					when "10001101000101001" => rgb <= "000000";
					when "10001101000101010" => rgb <= "000000";
					when "10001101000101011" => rgb <= "000000";
					when "10001101000101100" => rgb <= "000000";
					when "10001101000101101" => rgb <= "000000";
					when "10001101000101110" => rgb <= "000000";
					when "10001101000101111" => rgb <= "000000";
					when "10001101000110000" => rgb <= "000000";
					when "10001101000110001" => rgb <= "000000";
					when "10001101000110010" => rgb <= "000000";
					when "10001101000110011" => rgb <= "000000";
					when "10001101000110100" => rgb <= "000000";
					when "10001101000110101" => rgb <= "000000";
					when "10001101000110110" => rgb <= "000000";
					when "10001101000110111" => rgb <= "000000";
					when "10001101000111000" => rgb <= "000000";
					when "10001101000111001" => rgb <= "000000";
					when "10001101000111010" => rgb <= "000000";
					when "10001101000111011" => rgb <= "000000";
					when "10001101000111100" => rgb <= "000000";
					when "10001101000111101" => rgb <= "000000";
					when "10001101000111110" => rgb <= "000000";
					when "10001101000111111" => rgb <= "000000";
					when "10001101001000000" => rgb <= "000000";
					when "10001101001000001" => rgb <= "000000";
					when "10001101001000010" => rgb <= "000000";
					when "10001101001000011" => rgb <= "000000";
					when "10001101001000100" => rgb <= "000000";
					when "10001101001000101" => rgb <= "000000";
					when "10001101001000110" => rgb <= "000000";
					when "10001101001000111" => rgb <= "000000";
					when "10001101001001000" => rgb <= "000000";
					when "10001101001001001" => rgb <= "000000";
					when "10001101001001010" => rgb <= "000000";
					when "10001101001001011" => rgb <= "000000";
					when "10001101001001100" => rgb <= "000000";
					when "10001101001001101" => rgb <= "000000";
					when "10001101001001110" => rgb <= "000000";
					when "10001101001001111" => rgb <= "000000";
					when "10001101001010000" => rgb <= "000000";
					when "10001101001010001" => rgb <= "000000";
					when "10001101001010010" => rgb <= "000000";
					when "10001101001010011" => rgb <= "000000";
					when "10001101001010100" => rgb <= "000000";
					when "10001101001010101" => rgb <= "000000";
					when "10001101001010110" => rgb <= "000000";
					when "10001101001010111" => rgb <= "000000";
					when "10001101001011000" => rgb <= "000000";
					when "10001101001011001" => rgb <= "000000";
					when "10001101001011010" => rgb <= "000000";
					when "10001101001011011" => rgb <= "000000";
					when "10001101001011100" => rgb <= "000000";
					when "10001101001011101" => rgb <= "000000";
					when "10001101001011110" => rgb <= "000000";
					when "10001101001011111" => rgb <= "000000";
					when "10001101001100000" => rgb <= "000000";
					when "10001101001100001" => rgb <= "000000";
					when "10001101001100010" => rgb <= "000000";
					when "10001101001100011" => rgb <= "000000";
					when "10001101001100100" => rgb <= "000000";
					when "10001101001100101" => rgb <= "000000";
					when "10001101001100110" => rgb <= "000000";
					when "10001101001100111" => rgb <= "000000";
					when "10001101001101000" => rgb <= "000000";
					when "10001101001101001" => rgb <= "000000";
					when "10001101001101010" => rgb <= "000000";
					when "10001101001101011" => rgb <= "000000";
					when "10001101001101100" => rgb <= "000000";
					when "10001101001101101" => rgb <= "000000";
					when "10001101001101110" => rgb <= "000000";
					when "10001101001101111" => rgb <= "000000";
					when "10001101001110000" => rgb <= "000000";
					when "10001101001110001" => rgb <= "000000";
					when "10001101001110010" => rgb <= "000000";
					when "10001101001110011" => rgb <= "000000";
					when "10001101001110100" => rgb <= "000000";
					when "10001101001110101" => rgb <= "000000";
					when "10001101001110110" => rgb <= "000000";
					when "10001101001110111" => rgb <= "000000";
					when "10001101001111000" => rgb <= "000000";
					when "10001101001111001" => rgb <= "000000";
					when "10001101001111010" => rgb <= "000000";
					when "10001101001111011" => rgb <= "000000";
					when "10001101001111100" => rgb <= "000000";
					when "10001101001111101" => rgb <= "000000";
					when "10001101001111110" => rgb <= "000000";
					when "10001101001111111" => rgb <= "000000";
					when "10001101010000000" => rgb <= "000000";
					when "10001101010000001" => rgb <= "000000";
					when "10001101010000010" => rgb <= "000000";
					when "10001101010000011" => rgb <= "000000";
					when "10001101010000100" => rgb <= "000000";
					when "10001101010000101" => rgb <= "000000";
					when "10001101010000110" => rgb <= "000000";
					when "10001101010000111" => rgb <= "000000";
					when "10001101010001000" => rgb <= "000000";
					when "10001101010001001" => rgb <= "000000";
					when "10001101010001010" => rgb <= "000000";
					when "10001101010001011" => rgb <= "000000";
					when "10001101010001100" => rgb <= "000000";
					when "10001101010001101" => rgb <= "000000";
					when "10001101010001110" => rgb <= "000000";
					when "10001101010001111" => rgb <= "000000";
					when "10001101010010000" => rgb <= "000000";
					when "10001101010010001" => rgb <= "000000";
					when "10001101010010010" => rgb <= "000000";
					when "10001101010010011" => rgb <= "000000";
					when "10001101010010100" => rgb <= "000000";
					when "10001101010010101" => rgb <= "000000";
					when "10001101010010110" => rgb <= "000000";
					when "10001101010010111" => rgb <= "000000";
					when "10001101010011000" => rgb <= "000000";
					when "10001101010011001" => rgb <= "000000";
					when "10001101010011010" => rgb <= "000000";
					when "10001101010011011" => rgb <= "000000";
					when "10001101010011100" => rgb <= "000000";
					when "10001101010011101" => rgb <= "000000";
					when "10001101010011110" => rgb <= "000000";
					when "10001101010011111" => rgb <= "000000";
					when "10001101010100000" => rgb <= "000000";
					when "10001101010100001" => rgb <= "000000";
					when "10001101010100010" => rgb <= "000000";
					when "10001101010100011" => rgb <= "000000";
					when "10001101010100100" => rgb <= "000000";
					when "10001101010100101" => rgb <= "000000";
					when "10001101010100110" => rgb <= "000000";
					when "10001101010100111" => rgb <= "000000";
					when "10001101010101000" => rgb <= "000000";
					when "10001101010101001" => rgb <= "000000";
					when "10001101010101010" => rgb <= "000000";
					when "10001101010101011" => rgb <= "000000";
					when "10001101010101100" => rgb <= "000000";
					when "10001101010101101" => rgb <= "000000";
					when "10001101010101110" => rgb <= "000000";
					when "10001101010101111" => rgb <= "000000";
					when "10001101010110000" => rgb <= "000000";
					when "10001101010110001" => rgb <= "000000";
					when "10001101010110010" => rgb <= "000000";
					when "10001101010110011" => rgb <= "000000";
					when "10001101010110100" => rgb <= "000000";
					when "10001101010110101" => rgb <= "000000";
					when "10001101010110110" => rgb <= "000000";
					when "10001101010110111" => rgb <= "000000";
					when "10001101010111000" => rgb <= "000000";
					when "10001101010111001" => rgb <= "000000";
					when "10001101010111010" => rgb <= "000000";
					when "10001101010111011" => rgb <= "000000";
					when "10001101010111100" => rgb <= "000000";
					when "10001101010111101" => rgb <= "000000";
					when "10001101010111110" => rgb <= "000000";
					when "10001101010111111" => rgb <= "000000";
					when "10001101011000000" => rgb <= "000000";
					when "10001101011000001" => rgb <= "000000";
					when "10001101011000010" => rgb <= "000000";
					when "10001101011000011" => rgb <= "000000";
					when "10001101011000100" => rgb <= "000000";
					when "10001101011000101" => rgb <= "000000";
					when "10001101011000110" => rgb <= "000000";
					when "10001101011000111" => rgb <= "000000";
					when "10001101011001000" => rgb <= "000000";
					when "10001101011001001" => rgb <= "000000";
					when "10001101011001010" => rgb <= "000000";
					when "10001101011001011" => rgb <= "000000";
					when "10001101011001100" => rgb <= "000000";
					when "10001101011001101" => rgb <= "000000";
					when "10001101011001110" => rgb <= "000000";
					when "10001101011001111" => rgb <= "000000";
					when "10001101011010000" => rgb <= "000000";
					when "10001101011010001" => rgb <= "000000";
					when "10001101011010010" => rgb <= "000000";
					when "10001101011010011" => rgb <= "000000";
					when "10001101011010100" => rgb <= "000000";
					when "10001101011010101" => rgb <= "000000";
					when "10001101011010110" => rgb <= "000000";
					when "10001101011010111" => rgb <= "000000";
					when "10001101011011000" => rgb <= "000000";
					when "10001101011011001" => rgb <= "000000";
					when "10001101011011010" => rgb <= "000000";
					when "10001101011011011" => rgb <= "000000";
					when "10001101011011100" => rgb <= "000000";
					when "10001101011011101" => rgb <= "000000";
					when "10001101011011110" => rgb <= "000000";
					when "10001101011011111" => rgb <= "000000";
					when "10001101011100000" => rgb <= "000000";
					when "10001101011100001" => rgb <= "000000";
					when "10001101011100010" => rgb <= "000000";
					when "10001101011100011" => rgb <= "000000";
					when "10001101011100100" => rgb <= "000000";
					when "10001101011100101" => rgb <= "000000";
					when "10001101011100110" => rgb <= "000000";
					when "10001101011100111" => rgb <= "000000";
					when "10001101011101000" => rgb <= "000000";
					when "10001101011101001" => rgb <= "000000";
					when "10001101011101010" => rgb <= "000000";
					when "10001101011101011" => rgb <= "000000";
					when "10001101011101100" => rgb <= "000000";
					when "10001101011101101" => rgb <= "000000";
					when "10001101011101110" => rgb <= "000000";
					when "10001101011101111" => rgb <= "000000";
					when "10001101011110000" => rgb <= "000000";
					when "10001101011110001" => rgb <= "000000";
					when "10001101011110010" => rgb <= "000000";
					when "10001101011110011" => rgb <= "000000";
					when "10001101011110100" => rgb <= "000000";
					when "10001101011110101" => rgb <= "000000";
					when "10001101011110110" => rgb <= "000000";
					when "10001101011110111" => rgb <= "000000";
					when "10001101011111000" => rgb <= "000000";
					when "10001101011111001" => rgb <= "000000";
					when "10001101011111010" => rgb <= "000000";
					when "10001101011111011" => rgb <= "000000";
					when "10001101011111100" => rgb <= "000000";
					when "10001101011111101" => rgb <= "000000";
					when "10001101011111110" => rgb <= "000000";
					when "10001101011111111" => rgb <= "000000";
					when "10001101100000000" => rgb <= "000000";
					when "10001101100000001" => rgb <= "000000";
					when "10001101100000010" => rgb <= "000000";
					when "10001101100000011" => rgb <= "000000";
					when "10001101100000100" => rgb <= "000000";
					when "10001101100000101" => rgb <= "000000";
					when "10001101100000110" => rgb <= "000000";
					when "10001101100000111" => rgb <= "000000";
					when "10001101100001000" => rgb <= "000000";
					when "10001101100001001" => rgb <= "000000";
					when "10001101100001010" => rgb <= "000000";
					when "10001101100001011" => rgb <= "000000";
					when "10001101100001100" => rgb <= "000000";
					when "10001101100001101" => rgb <= "000000";
					when "10001101100001110" => rgb <= "000000";
					when "10001101100001111" => rgb <= "000000";
					when "10001101100010000" => rgb <= "000000";
					when "10001101100010001" => rgb <= "000000";
					when "10001101100010010" => rgb <= "000000";
					when "10001101100010011" => rgb <= "000000";
					when "10001101100010100" => rgb <= "000000";
					when "10001101100010101" => rgb <= "000000";
					when "10001101100010110" => rgb <= "000000";
					when "10001101100010111" => rgb <= "000000";
					when "10001101100011000" => rgb <= "000000";
					when "10001101100011001" => rgb <= "000000";
					when "10001101100011010" => rgb <= "000000";
					when "10001101100011011" => rgb <= "000000";
					when "10001101100011100" => rgb <= "000000";
					when "10001101100011101" => rgb <= "000000";
					when "10001101100011110" => rgb <= "000000";
					when "10001101100011111" => rgb <= "000000";
					when "10001101100100000" => rgb <= "000000";
					when "10001101100100001" => rgb <= "000000";
					when "10001101100100010" => rgb <= "000000";
					when "10001101100100011" => rgb <= "000000";
					when "10001101100100100" => rgb <= "000000";
					when "10001101100100101" => rgb <= "000000";
					when "10001101100100110" => rgb <= "000000";
					when "10001101100100111" => rgb <= "000000";
					when "10001101100101000" => rgb <= "000000";
					when "10001101100101001" => rgb <= "000000";
					when "10001101100101010" => rgb <= "000000";
					when "10001101100101011" => rgb <= "000000";
					when "10001101100101100" => rgb <= "000000";
					when "10001101100101101" => rgb <= "000000";
					when "10001101100101110" => rgb <= "000000";
					when "10001101100101111" => rgb <= "000000";
					when "10001101100110000" => rgb <= "000000";
					when "10001101100110001" => rgb <= "000000";
					when "10001101100110010" => rgb <= "000000";
					when "10001101100110011" => rgb <= "000000";
					when "10001101100110100" => rgb <= "000000";
					when "10001101100110101" => rgb <= "000000";
					when "10001101100110110" => rgb <= "000000";
					when "10001101100110111" => rgb <= "000000";
					when "10001101100111000" => rgb <= "000000";
					when "10001101100111001" => rgb <= "000000";
					when "10001101100111010" => rgb <= "000000";
					when "10001101100111011" => rgb <= "000000";
					when "10001101100111100" => rgb <= "000000";
					when "10001101100111101" => rgb <= "000000";
					when "10001101100111110" => rgb <= "000000";
					when "10001101100111111" => rgb <= "000000";
					when "10001110000000000" => rgb <= "000000";
					when "10001110000000001" => rgb <= "000000";
					when "10001110000000010" => rgb <= "000000";
					when "10001110000000011" => rgb <= "000000";
					when "10001110000000100" => rgb <= "000000";
					when "10001110000000101" => rgb <= "000000";
					when "10001110000000110" => rgb <= "000000";
					when "10001110000000111" => rgb <= "000000";
					when "10001110000001000" => rgb <= "000000";
					when "10001110000001001" => rgb <= "000000";
					when "10001110000001010" => rgb <= "000000";
					when "10001110000001011" => rgb <= "000000";
					when "10001110000001100" => rgb <= "000000";
					when "10001110000001101" => rgb <= "000000";
					when "10001110000001110" => rgb <= "000000";
					when "10001110000001111" => rgb <= "000000";
					when "10001110000010000" => rgb <= "000000";
					when "10001110000010001" => rgb <= "000000";
					when "10001110000010010" => rgb <= "000000";
					when "10001110000010011" => rgb <= "000000";
					when "10001110000010100" => rgb <= "000000";
					when "10001110000010101" => rgb <= "000000";
					when "10001110000010110" => rgb <= "000000";
					when "10001110000010111" => rgb <= "000000";
					when "10001110000011000" => rgb <= "000000";
					when "10001110000011001" => rgb <= "000000";
					when "10001110000011010" => rgb <= "000000";
					when "10001110000011011" => rgb <= "000000";
					when "10001110000011100" => rgb <= "000000";
					when "10001110000011101" => rgb <= "000000";
					when "10001110000011110" => rgb <= "000000";
					when "10001110000011111" => rgb <= "000000";
					when "10001110000100000" => rgb <= "000000";
					when "10001110000100001" => rgb <= "000000";
					when "10001110000100010" => rgb <= "000000";
					when "10001110000100011" => rgb <= "000000";
					when "10001110000100100" => rgb <= "000000";
					when "10001110000100101" => rgb <= "000000";
					when "10001110000100110" => rgb <= "000000";
					when "10001110000100111" => rgb <= "000000";
					when "10001110000101000" => rgb <= "000000";
					when "10001110000101001" => rgb <= "000000";
					when "10001110000101010" => rgb <= "000000";
					when "10001110000101011" => rgb <= "000000";
					when "10001110000101100" => rgb <= "000000";
					when "10001110000101101" => rgb <= "000000";
					when "10001110000101110" => rgb <= "000000";
					when "10001110000101111" => rgb <= "000000";
					when "10001110000110000" => rgb <= "000000";
					when "10001110000110001" => rgb <= "000000";
					when "10001110000110010" => rgb <= "000000";
					when "10001110000110011" => rgb <= "000000";
					when "10001110000110100" => rgb <= "000000";
					when "10001110000110101" => rgb <= "000000";
					when "10001110000110110" => rgb <= "000000";
					when "10001110000110111" => rgb <= "000000";
					when "10001110000111000" => rgb <= "000000";
					when "10001110000111001" => rgb <= "000000";
					when "10001110000111010" => rgb <= "000000";
					when "10001110000111011" => rgb <= "000000";
					when "10001110000111100" => rgb <= "000000";
					when "10001110000111101" => rgb <= "000000";
					when "10001110000111110" => rgb <= "000000";
					when "10001110000111111" => rgb <= "000000";
					when "10001110001000000" => rgb <= "000000";
					when "10001110001000001" => rgb <= "000000";
					when "10001110001000010" => rgb <= "000000";
					when "10001110001000011" => rgb <= "000000";
					when "10001110001000100" => rgb <= "000000";
					when "10001110001000101" => rgb <= "000000";
					when "10001110001000110" => rgb <= "000000";
					when "10001110001000111" => rgb <= "000000";
					when "10001110001001000" => rgb <= "000000";
					when "10001110001001001" => rgb <= "000000";
					when "10001110001001010" => rgb <= "000000";
					when "10001110001001011" => rgb <= "000000";
					when "10001110001001100" => rgb <= "000000";
					when "10001110001001101" => rgb <= "000000";
					when "10001110001001110" => rgb <= "000000";
					when "10001110001001111" => rgb <= "000000";
					when "10001110001010000" => rgb <= "000000";
					when "10001110001010001" => rgb <= "000000";
					when "10001110001010010" => rgb <= "000000";
					when "10001110001010011" => rgb <= "000000";
					when "10001110001010100" => rgb <= "000000";
					when "10001110001010101" => rgb <= "000000";
					when "10001110001010110" => rgb <= "000000";
					when "10001110001010111" => rgb <= "000000";
					when "10001110001011000" => rgb <= "000000";
					when "10001110001011001" => rgb <= "000000";
					when "10001110001011010" => rgb <= "000000";
					when "10001110001011011" => rgb <= "000000";
					when "10001110001011100" => rgb <= "000000";
					when "10001110001011101" => rgb <= "000000";
					when "10001110001011110" => rgb <= "000000";
					when "10001110001011111" => rgb <= "000000";
					when "10001110001100000" => rgb <= "000000";
					when "10001110001100001" => rgb <= "000000";
					when "10001110001100010" => rgb <= "000000";
					when "10001110001100011" => rgb <= "000000";
					when "10001110001100100" => rgb <= "000000";
					when "10001110001100101" => rgb <= "000000";
					when "10001110001100110" => rgb <= "000000";
					when "10001110001100111" => rgb <= "000000";
					when "10001110001101000" => rgb <= "000000";
					when "10001110001101001" => rgb <= "000000";
					when "10001110001101010" => rgb <= "000000";
					when "10001110001101011" => rgb <= "000000";
					when "10001110001101100" => rgb <= "000000";
					when "10001110001101101" => rgb <= "000000";
					when "10001110001101110" => rgb <= "000000";
					when "10001110001101111" => rgb <= "000000";
					when "10001110001110000" => rgb <= "000000";
					when "10001110001110001" => rgb <= "000000";
					when "10001110001110010" => rgb <= "000000";
					when "10001110001110011" => rgb <= "000000";
					when "10001110001110100" => rgb <= "000000";
					when "10001110001110101" => rgb <= "000000";
					when "10001110001110110" => rgb <= "000000";
					when "10001110001110111" => rgb <= "000000";
					when "10001110001111000" => rgb <= "000000";
					when "10001110001111001" => rgb <= "000000";
					when "10001110001111010" => rgb <= "000000";
					when "10001110001111011" => rgb <= "000000";
					when "10001110001111100" => rgb <= "000000";
					when "10001110001111101" => rgb <= "000000";
					when "10001110001111110" => rgb <= "000000";
					when "10001110001111111" => rgb <= "000000";
					when "10001110010000000" => rgb <= "000000";
					when "10001110010000001" => rgb <= "000000";
					when "10001110010000010" => rgb <= "000000";
					when "10001110010000011" => rgb <= "000000";
					when "10001110010000100" => rgb <= "000000";
					when "10001110010000101" => rgb <= "000000";
					when "10001110010000110" => rgb <= "000000";
					when "10001110010000111" => rgb <= "000000";
					when "10001110010001000" => rgb <= "000000";
					when "10001110010001001" => rgb <= "000000";
					when "10001110010001010" => rgb <= "000000";
					when "10001110010001011" => rgb <= "000000";
					when "10001110010001100" => rgb <= "000000";
					when "10001110010001101" => rgb <= "000000";
					when "10001110010001110" => rgb <= "000000";
					when "10001110010001111" => rgb <= "000000";
					when "10001110010010000" => rgb <= "000000";
					when "10001110010010001" => rgb <= "000000";
					when "10001110010010010" => rgb <= "000000";
					when "10001110010010011" => rgb <= "000000";
					when "10001110010010100" => rgb <= "000000";
					when "10001110010010101" => rgb <= "000000";
					when "10001110010010110" => rgb <= "000000";
					when "10001110010010111" => rgb <= "000000";
					when "10001110010011000" => rgb <= "000000";
					when "10001110010011001" => rgb <= "000000";
					when "10001110010011010" => rgb <= "000000";
					when "10001110010011011" => rgb <= "000000";
					when "10001110010011100" => rgb <= "000000";
					when "10001110010011101" => rgb <= "000000";
					when "10001110010011110" => rgb <= "000000";
					when "10001110010011111" => rgb <= "000000";
					when "10001110010100000" => rgb <= "000000";
					when "10001110010100001" => rgb <= "000000";
					when "10001110010100010" => rgb <= "000000";
					when "10001110010100011" => rgb <= "000000";
					when "10001110010100100" => rgb <= "000000";
					when "10001110010100101" => rgb <= "000000";
					when "10001110010100110" => rgb <= "000000";
					when "10001110010100111" => rgb <= "000000";
					when "10001110010101000" => rgb <= "000000";
					when "10001110010101001" => rgb <= "000000";
					when "10001110010101010" => rgb <= "000000";
					when "10001110010101011" => rgb <= "000000";
					when "10001110010101100" => rgb <= "000000";
					when "10001110010101101" => rgb <= "000000";
					when "10001110010101110" => rgb <= "000000";
					when "10001110010101111" => rgb <= "000000";
					when "10001110010110000" => rgb <= "000000";
					when "10001110010110001" => rgb <= "000000";
					when "10001110010110010" => rgb <= "000000";
					when "10001110010110011" => rgb <= "000000";
					when "10001110010110100" => rgb <= "000000";
					when "10001110010110101" => rgb <= "000000";
					when "10001110010110110" => rgb <= "000000";
					when "10001110010110111" => rgb <= "000000";
					when "10001110010111000" => rgb <= "000000";
					when "10001110010111001" => rgb <= "000000";
					when "10001110010111010" => rgb <= "000000";
					when "10001110010111011" => rgb <= "000000";
					when "10001110010111100" => rgb <= "000000";
					when "10001110010111101" => rgb <= "000000";
					when "10001110010111110" => rgb <= "000000";
					when "10001110010111111" => rgb <= "000000";
					when "10001110011000000" => rgb <= "000000";
					when "10001110011000001" => rgb <= "000000";
					when "10001110011000010" => rgb <= "000000";
					when "10001110011000011" => rgb <= "000000";
					when "10001110011000100" => rgb <= "000000";
					when "10001110011000101" => rgb <= "000000";
					when "10001110011000110" => rgb <= "000000";
					when "10001110011000111" => rgb <= "000000";
					when "10001110011001000" => rgb <= "000000";
					when "10001110011001001" => rgb <= "000000";
					when "10001110011001010" => rgb <= "000000";
					when "10001110011001011" => rgb <= "000000";
					when "10001110011001100" => rgb <= "000000";
					when "10001110011001101" => rgb <= "000000";
					when "10001110011001110" => rgb <= "000000";
					when "10001110011001111" => rgb <= "000000";
					when "10001110011010000" => rgb <= "000000";
					when "10001110011010001" => rgb <= "000000";
					when "10001110011010010" => rgb <= "000000";
					when "10001110011010011" => rgb <= "000000";
					when "10001110011010100" => rgb <= "000000";
					when "10001110011010101" => rgb <= "000000";
					when "10001110011010110" => rgb <= "000000";
					when "10001110011010111" => rgb <= "000000";
					when "10001110011011000" => rgb <= "000000";
					when "10001110011011001" => rgb <= "000000";
					when "10001110011011010" => rgb <= "000000";
					when "10001110011011011" => rgb <= "000000";
					when "10001110011011100" => rgb <= "000000";
					when "10001110011011101" => rgb <= "000000";
					when "10001110011011110" => rgb <= "000000";
					when "10001110011011111" => rgb <= "000000";
					when "10001110011100000" => rgb <= "000000";
					when "10001110011100001" => rgb <= "000000";
					when "10001110011100010" => rgb <= "000000";
					when "10001110011100011" => rgb <= "000000";
					when "10001110011100100" => rgb <= "000000";
					when "10001110011100101" => rgb <= "000000";
					when "10001110011100110" => rgb <= "000000";
					when "10001110011100111" => rgb <= "000000";
					when "10001110011101000" => rgb <= "000000";
					when "10001110011101001" => rgb <= "000000";
					when "10001110011101010" => rgb <= "000000";
					when "10001110011101011" => rgb <= "000000";
					when "10001110011101100" => rgb <= "000000";
					when "10001110011101101" => rgb <= "000000";
					when "10001110011101110" => rgb <= "000000";
					when "10001110011101111" => rgb <= "000000";
					when "10001110011110000" => rgb <= "000000";
					when "10001110011110001" => rgb <= "000000";
					when "10001110011110010" => rgb <= "000000";
					when "10001110011110011" => rgb <= "000000";
					when "10001110011110100" => rgb <= "000000";
					when "10001110011110101" => rgb <= "000000";
					when "10001110011110110" => rgb <= "000000";
					when "10001110011110111" => rgb <= "000000";
					when "10001110011111000" => rgb <= "000000";
					when "10001110011111001" => rgb <= "000000";
					when "10001110011111010" => rgb <= "000000";
					when "10001110011111011" => rgb <= "000000";
					when "10001110011111100" => rgb <= "000000";
					when "10001110011111101" => rgb <= "000000";
					when "10001110011111110" => rgb <= "000000";
					when "10001110011111111" => rgb <= "000000";
					when "10001110100000000" => rgb <= "000000";
					when "10001110100000001" => rgb <= "000000";
					when "10001110100000010" => rgb <= "000000";
					when "10001110100000011" => rgb <= "000000";
					when "10001110100000100" => rgb <= "000000";
					when "10001110100000101" => rgb <= "000000";
					when "10001110100000110" => rgb <= "000000";
					when "10001110100000111" => rgb <= "000000";
					when "10001110100001000" => rgb <= "000000";
					when "10001110100001001" => rgb <= "000000";
					when "10001110100001010" => rgb <= "000000";
					when "10001110100001011" => rgb <= "000000";
					when "10001110100001100" => rgb <= "000000";
					when "10001110100001101" => rgb <= "000000";
					when "10001110100001110" => rgb <= "000000";
					when "10001110100001111" => rgb <= "000000";
					when "10001110100010000" => rgb <= "000000";
					when "10001110100010001" => rgb <= "000000";
					when "10001110100010010" => rgb <= "000000";
					when "10001110100010011" => rgb <= "000000";
					when "10001110100010100" => rgb <= "000000";
					when "10001110100010101" => rgb <= "000000";
					when "10001110100010110" => rgb <= "000000";
					when "10001110100010111" => rgb <= "000000";
					when "10001110100011000" => rgb <= "000000";
					when "10001110100011001" => rgb <= "000000";
					when "10001110100011010" => rgb <= "000000";
					when "10001110100011011" => rgb <= "000000";
					when "10001110100011100" => rgb <= "000000";
					when "10001110100011101" => rgb <= "000000";
					when "10001110100011110" => rgb <= "000000";
					when "10001110100011111" => rgb <= "000000";
					when "10001110100100000" => rgb <= "000000";
					when "10001110100100001" => rgb <= "000000";
					when "10001110100100010" => rgb <= "000000";
					when "10001110100100011" => rgb <= "000000";
					when "10001110100100100" => rgb <= "000000";
					when "10001110100100101" => rgb <= "000000";
					when "10001110100100110" => rgb <= "000000";
					when "10001110100100111" => rgb <= "000000";
					when "10001110100101000" => rgb <= "000000";
					when "10001110100101001" => rgb <= "000000";
					when "10001110100101010" => rgb <= "000000";
					when "10001110100101011" => rgb <= "000000";
					when "10001110100101100" => rgb <= "000000";
					when "10001110100101101" => rgb <= "000000";
					when "10001110100101110" => rgb <= "000000";
					when "10001110100101111" => rgb <= "000000";
					when "10001110100110000" => rgb <= "000000";
					when "10001110100110001" => rgb <= "000000";
					when "10001110100110010" => rgb <= "000000";
					when "10001110100110011" => rgb <= "000000";
					when "10001110100110100" => rgb <= "000000";
					when "10001110100110101" => rgb <= "000000";
					when "10001110100110110" => rgb <= "000000";
					when "10001110100110111" => rgb <= "000000";
					when "10001110100111000" => rgb <= "000000";
					when "10001110100111001" => rgb <= "000000";
					when "10001110100111010" => rgb <= "000000";
					when "10001110100111011" => rgb <= "000000";
					when "10001110100111100" => rgb <= "000000";
					when "10001110100111101" => rgb <= "000000";
					when "10001110100111110" => rgb <= "000000";
					when "10001110100111111" => rgb <= "000000";
					when "10001111000000000" => rgb <= "000000";
					when "10001111000000001" => rgb <= "000000";
					when "10001111000000010" => rgb <= "000000";
					when "10001111000000011" => rgb <= "000000";
					when "10001111000000100" => rgb <= "000000";
					when "10001111000000101" => rgb <= "000000";
					when "10001111000000110" => rgb <= "000000";
					when "10001111000000111" => rgb <= "000000";
					when "10001111000001000" => rgb <= "000000";
					when "10001111000001001" => rgb <= "000000";
					when "10001111000001010" => rgb <= "000000";
					when "10001111000001011" => rgb <= "000000";
					when "10001111000001100" => rgb <= "000000";
					when "10001111000001101" => rgb <= "000000";
					when "10001111000001110" => rgb <= "000000";
					when "10001111000001111" => rgb <= "000000";
					when "10001111000010000" => rgb <= "000000";
					when "10001111000010001" => rgb <= "000000";
					when "10001111000010010" => rgb <= "000000";
					when "10001111000010011" => rgb <= "000000";
					when "10001111000010100" => rgb <= "000000";
					when "10001111000010101" => rgb <= "000000";
					when "10001111000010110" => rgb <= "000000";
					when "10001111000010111" => rgb <= "000000";
					when "10001111000011000" => rgb <= "000000";
					when "10001111000011001" => rgb <= "000000";
					when "10001111000011010" => rgb <= "000000";
					when "10001111000011011" => rgb <= "000000";
					when "10001111000011100" => rgb <= "000000";
					when "10001111000011101" => rgb <= "000000";
					when "10001111000011110" => rgb <= "000000";
					when "10001111000011111" => rgb <= "000000";
					when "10001111000100000" => rgb <= "000000";
					when "10001111000100001" => rgb <= "000000";
					when "10001111000100010" => rgb <= "000000";
					when "10001111000100011" => rgb <= "000000";
					when "10001111000100100" => rgb <= "000000";
					when "10001111000100101" => rgb <= "000000";
					when "10001111000100110" => rgb <= "000000";
					when "10001111000100111" => rgb <= "000000";
					when "10001111000101000" => rgb <= "000000";
					when "10001111000101001" => rgb <= "000000";
					when "10001111000101010" => rgb <= "000000";
					when "10001111000101011" => rgb <= "000000";
					when "10001111000101100" => rgb <= "000000";
					when "10001111000101101" => rgb <= "000000";
					when "10001111000101110" => rgb <= "000000";
					when "10001111000101111" => rgb <= "000000";
					when "10001111000110000" => rgb <= "000000";
					when "10001111000110001" => rgb <= "000000";
					when "10001111000110010" => rgb <= "000000";
					when "10001111000110011" => rgb <= "000000";
					when "10001111000110100" => rgb <= "000000";
					when "10001111000110101" => rgb <= "000000";
					when "10001111000110110" => rgb <= "000000";
					when "10001111000110111" => rgb <= "000000";
					when "10001111000111000" => rgb <= "000000";
					when "10001111000111001" => rgb <= "000000";
					when "10001111000111010" => rgb <= "000000";
					when "10001111000111011" => rgb <= "000000";
					when "10001111000111100" => rgb <= "000000";
					when "10001111000111101" => rgb <= "000000";
					when "10001111000111110" => rgb <= "000000";
					when "10001111000111111" => rgb <= "000000";
					when "10001111001000000" => rgb <= "000000";
					when "10001111001000001" => rgb <= "000000";
					when "10001111001000010" => rgb <= "000000";
					when "10001111001000011" => rgb <= "000000";
					when "10001111001000100" => rgb <= "000000";
					when "10001111001000101" => rgb <= "000000";
					when "10001111001000110" => rgb <= "000000";
					when "10001111001000111" => rgb <= "000000";
					when "10001111001001000" => rgb <= "000000";
					when "10001111001001001" => rgb <= "000000";
					when "10001111001001010" => rgb <= "000000";
					when "10001111001001011" => rgb <= "000000";
					when "10001111001001100" => rgb <= "000000";
					when "10001111001001101" => rgb <= "000000";
					when "10001111001001110" => rgb <= "000000";
					when "10001111001001111" => rgb <= "000000";
					when "10001111001010000" => rgb <= "000000";
					when "10001111001010001" => rgb <= "000000";
					when "10001111001010010" => rgb <= "000000";
					when "10001111001010011" => rgb <= "000000";
					when "10001111001010100" => rgb <= "000000";
					when "10001111001010101" => rgb <= "000000";
					when "10001111001010110" => rgb <= "000000";
					when "10001111001010111" => rgb <= "000000";
					when "10001111001011000" => rgb <= "000000";
					when "10001111001011001" => rgb <= "000000";
					when "10001111001011010" => rgb <= "000000";
					when "10001111001011011" => rgb <= "000000";
					when "10001111001011100" => rgb <= "000000";
					when "10001111001011101" => rgb <= "000000";
					when "10001111001011110" => rgb <= "000000";
					when "10001111001011111" => rgb <= "000000";
					when "10001111001100000" => rgb <= "000000";
					when "10001111001100001" => rgb <= "000000";
					when "10001111001100010" => rgb <= "000000";
					when "10001111001100011" => rgb <= "000000";
					when "10001111001100100" => rgb <= "000000";
					when "10001111001100101" => rgb <= "000000";
					when "10001111001100110" => rgb <= "000000";
					when "10001111001100111" => rgb <= "000000";
					when "10001111001101000" => rgb <= "000000";
					when "10001111001101001" => rgb <= "000000";
					when "10001111001101010" => rgb <= "000000";
					when "10001111001101011" => rgb <= "000000";
					when "10001111001101100" => rgb <= "000000";
					when "10001111001101101" => rgb <= "000000";
					when "10001111001101110" => rgb <= "000000";
					when "10001111001101111" => rgb <= "000000";
					when "10001111001110000" => rgb <= "000000";
					when "10001111001110001" => rgb <= "000000";
					when "10001111001110010" => rgb <= "000000";
					when "10001111001110011" => rgb <= "000000";
					when "10001111001110100" => rgb <= "000000";
					when "10001111001110101" => rgb <= "000000";
					when "10001111001110110" => rgb <= "000000";
					when "10001111001110111" => rgb <= "000000";
					when "10001111001111000" => rgb <= "000000";
					when "10001111001111001" => rgb <= "000000";
					when "10001111001111010" => rgb <= "000000";
					when "10001111001111011" => rgb <= "000000";
					when "10001111001111100" => rgb <= "000000";
					when "10001111001111101" => rgb <= "000000";
					when "10001111001111110" => rgb <= "000000";
					when "10001111001111111" => rgb <= "000000";
					when "10001111010000000" => rgb <= "000000";
					when "10001111010000001" => rgb <= "000000";
					when "10001111010000010" => rgb <= "000000";
					when "10001111010000011" => rgb <= "000000";
					when "10001111010000100" => rgb <= "000000";
					when "10001111010000101" => rgb <= "000000";
					when "10001111010000110" => rgb <= "000000";
					when "10001111010000111" => rgb <= "000000";
					when "10001111010001000" => rgb <= "000000";
					when "10001111010001001" => rgb <= "000000";
					when "10001111010001010" => rgb <= "000000";
					when "10001111010001011" => rgb <= "000000";
					when "10001111010001100" => rgb <= "000000";
					when "10001111010001101" => rgb <= "000000";
					when "10001111010001110" => rgb <= "000000";
					when "10001111010001111" => rgb <= "000000";
					when "10001111010010000" => rgb <= "000000";
					when "10001111010010001" => rgb <= "000000";
					when "10001111010010010" => rgb <= "000000";
					when "10001111010010011" => rgb <= "000000";
					when "10001111010010100" => rgb <= "000000";
					when "10001111010010101" => rgb <= "000000";
					when "10001111010010110" => rgb <= "000000";
					when "10001111010010111" => rgb <= "000000";
					when "10001111010011000" => rgb <= "000000";
					when "10001111010011001" => rgb <= "000000";
					when "10001111010011010" => rgb <= "000000";
					when "10001111010011011" => rgb <= "000000";
					when "10001111010011100" => rgb <= "000000";
					when "10001111010011101" => rgb <= "000000";
					when "10001111010011110" => rgb <= "000000";
					when "10001111010011111" => rgb <= "000000";
					when "10001111010100000" => rgb <= "000000";
					when "10001111010100001" => rgb <= "000000";
					when "10001111010100010" => rgb <= "000000";
					when "10001111010100011" => rgb <= "000000";
					when "10001111010100100" => rgb <= "000000";
					when "10001111010100101" => rgb <= "000000";
					when "10001111010100110" => rgb <= "000000";
					when "10001111010100111" => rgb <= "000000";
					when "10001111010101000" => rgb <= "000000";
					when "10001111010101001" => rgb <= "000000";
					when "10001111010101010" => rgb <= "000000";
					when "10001111010101011" => rgb <= "000000";
					when "10001111010101100" => rgb <= "000000";
					when "10001111010101101" => rgb <= "000000";
					when "10001111010101110" => rgb <= "000000";
					when "10001111010101111" => rgb <= "000000";
					when "10001111010110000" => rgb <= "000000";
					when "10001111010110001" => rgb <= "000000";
					when "10001111010110010" => rgb <= "000000";
					when "10001111010110011" => rgb <= "000000";
					when "10001111010110100" => rgb <= "000000";
					when "10001111010110101" => rgb <= "000000";
					when "10001111010110110" => rgb <= "000000";
					when "10001111010110111" => rgb <= "000000";
					when "10001111010111000" => rgb <= "000000";
					when "10001111010111001" => rgb <= "000000";
					when "10001111010111010" => rgb <= "000000";
					when "10001111010111011" => rgb <= "000000";
					when "10001111010111100" => rgb <= "000000";
					when "10001111010111101" => rgb <= "000000";
					when "10001111010111110" => rgb <= "000000";
					when "10001111010111111" => rgb <= "000000";
					when "10001111011000000" => rgb <= "000000";
					when "10001111011000001" => rgb <= "000000";
					when "10001111011000010" => rgb <= "000000";
					when "10001111011000011" => rgb <= "000000";
					when "10001111011000100" => rgb <= "000000";
					when "10001111011000101" => rgb <= "000000";
					when "10001111011000110" => rgb <= "000000";
					when "10001111011000111" => rgb <= "000000";
					when "10001111011001000" => rgb <= "000000";
					when "10001111011001001" => rgb <= "000000";
					when "10001111011001010" => rgb <= "000000";
					when "10001111011001011" => rgb <= "000000";
					when "10001111011001100" => rgb <= "000000";
					when "10001111011001101" => rgb <= "000000";
					when "10001111011001110" => rgb <= "000000";
					when "10001111011001111" => rgb <= "000000";
					when "10001111011010000" => rgb <= "000000";
					when "10001111011010001" => rgb <= "000000";
					when "10001111011010010" => rgb <= "000000";
					when "10001111011010011" => rgb <= "000000";
					when "10001111011010100" => rgb <= "000000";
					when "10001111011010101" => rgb <= "000000";
					when "10001111011010110" => rgb <= "000000";
					when "10001111011010111" => rgb <= "000000";
					when "10001111011011000" => rgb <= "000000";
					when "10001111011011001" => rgb <= "000000";
					when "10001111011011010" => rgb <= "000000";
					when "10001111011011011" => rgb <= "000000";
					when "10001111011011100" => rgb <= "000000";
					when "10001111011011101" => rgb <= "000000";
					when "10001111011011110" => rgb <= "000000";
					when "10001111011011111" => rgb <= "000000";
					when "10001111011100000" => rgb <= "000000";
					when "10001111011100001" => rgb <= "000000";
					when "10001111011100010" => rgb <= "000000";
					when "10001111011100011" => rgb <= "000000";
					when "10001111011100100" => rgb <= "000000";
					when "10001111011100101" => rgb <= "000000";
					when "10001111011100110" => rgb <= "000000";
					when "10001111011100111" => rgb <= "000000";
					when "10001111011101000" => rgb <= "000000";
					when "10001111011101001" => rgb <= "000000";
					when "10001111011101010" => rgb <= "000000";
					when "10001111011101011" => rgb <= "000000";
					when "10001111011101100" => rgb <= "000000";
					when "10001111011101101" => rgb <= "000000";
					when "10001111011101110" => rgb <= "000000";
					when "10001111011101111" => rgb <= "000000";
					when "10001111011110000" => rgb <= "000000";
					when "10001111011110001" => rgb <= "000000";
					when "10001111011110010" => rgb <= "000000";
					when "10001111011110011" => rgb <= "000000";
					when "10001111011110100" => rgb <= "000000";
					when "10001111011110101" => rgb <= "000000";
					when "10001111011110110" => rgb <= "000000";
					when "10001111011110111" => rgb <= "000000";
					when "10001111011111000" => rgb <= "000000";
					when "10001111011111001" => rgb <= "000000";
					when "10001111011111010" => rgb <= "000000";
					when "10001111011111011" => rgb <= "000000";
					when "10001111011111100" => rgb <= "000000";
					when "10001111011111101" => rgb <= "000000";
					when "10001111011111110" => rgb <= "000000";
					when "10001111011111111" => rgb <= "000000";
					when "10001111100000000" => rgb <= "000000";
					when "10001111100000001" => rgb <= "000000";
					when "10001111100000010" => rgb <= "000000";
					when "10001111100000011" => rgb <= "000000";
					when "10001111100000100" => rgb <= "000000";
					when "10001111100000101" => rgb <= "000000";
					when "10001111100000110" => rgb <= "000000";
					when "10001111100000111" => rgb <= "000000";
					when "10001111100001000" => rgb <= "000000";
					when "10001111100001001" => rgb <= "000000";
					when "10001111100001010" => rgb <= "000000";
					when "10001111100001011" => rgb <= "000000";
					when "10001111100001100" => rgb <= "000000";
					when "10001111100001101" => rgb <= "000000";
					when "10001111100001110" => rgb <= "000000";
					when "10001111100001111" => rgb <= "000000";
					when "10001111100010000" => rgb <= "000000";
					when "10001111100010001" => rgb <= "000000";
					when "10001111100010010" => rgb <= "000000";
					when "10001111100010011" => rgb <= "000000";
					when "10001111100010100" => rgb <= "000000";
					when "10001111100010101" => rgb <= "000000";
					when "10001111100010110" => rgb <= "000000";
					when "10001111100010111" => rgb <= "000000";
					when "10001111100011000" => rgb <= "000000";
					when "10001111100011001" => rgb <= "000000";
					when "10001111100011010" => rgb <= "000000";
					when "10001111100011011" => rgb <= "000000";
					when "10001111100011100" => rgb <= "000000";
					when "10001111100011101" => rgb <= "000000";
					when "10001111100011110" => rgb <= "000000";
					when "10001111100011111" => rgb <= "000000";
					when "10001111100100000" => rgb <= "000000";
					when "10001111100100001" => rgb <= "000000";
					when "10001111100100010" => rgb <= "000000";
					when "10001111100100011" => rgb <= "000000";
					when "10001111100100100" => rgb <= "000000";
					when "10001111100100101" => rgb <= "000000";
					when "10001111100100110" => rgb <= "000000";
					when "10001111100100111" => rgb <= "000000";
					when "10001111100101000" => rgb <= "000000";
					when "10001111100101001" => rgb <= "000000";
					when "10001111100101010" => rgb <= "000000";
					when "10001111100101011" => rgb <= "000000";
					when "10001111100101100" => rgb <= "000000";
					when "10001111100101101" => rgb <= "000000";
					when "10001111100101110" => rgb <= "000000";
					when "10001111100101111" => rgb <= "000000";
					when "10001111100110000" => rgb <= "000000";
					when "10001111100110001" => rgb <= "000000";
					when "10001111100110010" => rgb <= "000000";
					when "10001111100110011" => rgb <= "000000";
					when "10001111100110100" => rgb <= "000000";
					when "10001111100110101" => rgb <= "000000";
					when "10001111100110110" => rgb <= "000000";
					when "10001111100110111" => rgb <= "000000";
					when "10001111100111000" => rgb <= "000000";
					when "10001111100111001" => rgb <= "000000";
					when "10001111100111010" => rgb <= "000000";
					when "10001111100111011" => rgb <= "000000";
					when "10001111100111100" => rgb <= "000000";
					when "10001111100111101" => rgb <= "000000";
					when "10001111100111110" => rgb <= "000000";
					when "10001111100111111" => rgb <= "000000";
					when "10010000000000000" => rgb <= "000000";
					when "10010000000000001" => rgb <= "000000";
					when "10010000000000010" => rgb <= "000000";
					when "10010000000000011" => rgb <= "000000";
					when "10010000000000100" => rgb <= "000000";
					when "10010000000000101" => rgb <= "000000";
					when "10010000000000110" => rgb <= "000000";
					when "10010000000000111" => rgb <= "000000";
					when "10010000000001000" => rgb <= "000000";
					when "10010000000001001" => rgb <= "000000";
					when "10010000000001010" => rgb <= "000000";
					when "10010000000001011" => rgb <= "000000";
					when "10010000000001100" => rgb <= "000000";
					when "10010000000001101" => rgb <= "000000";
					when "10010000000001110" => rgb <= "000000";
					when "10010000000001111" => rgb <= "000000";
					when "10010000000010000" => rgb <= "000000";
					when "10010000000010001" => rgb <= "000000";
					when "10010000000010010" => rgb <= "000000";
					when "10010000000010011" => rgb <= "000000";
					when "10010000000010100" => rgb <= "000000";
					when "10010000000010101" => rgb <= "000000";
					when "10010000000010110" => rgb <= "000000";
					when "10010000000010111" => rgb <= "000000";
					when "10010000000011000" => rgb <= "000000";
					when "10010000000011001" => rgb <= "000000";
					when "10010000000011010" => rgb <= "000000";
					when "10010000000011011" => rgb <= "000000";
					when "10010000000011100" => rgb <= "000000";
					when "10010000000011101" => rgb <= "000000";
					when "10010000000011110" => rgb <= "000000";
					when "10010000000011111" => rgb <= "000000";
					when "10010000000100000" => rgb <= "000000";
					when "10010000000100001" => rgb <= "000000";
					when "10010000000100010" => rgb <= "000000";
					when "10010000000100011" => rgb <= "000000";
					when "10010000000100100" => rgb <= "000000";
					when "10010000000100101" => rgb <= "000000";
					when "10010000000100110" => rgb <= "000000";
					when "10010000000100111" => rgb <= "000000";
					when "10010000000101000" => rgb <= "000000";
					when "10010000000101001" => rgb <= "000000";
					when "10010000000101010" => rgb <= "000000";
					when "10010000000101011" => rgb <= "000000";
					when "10010000000101100" => rgb <= "000000";
					when "10010000000101101" => rgb <= "000000";
					when "10010000000101110" => rgb <= "000000";
					when "10010000000101111" => rgb <= "000000";
					when "10010000000110000" => rgb <= "000000";
					when "10010000000110001" => rgb <= "000000";
					when "10010000000110010" => rgb <= "000000";
					when "10010000000110011" => rgb <= "000000";
					when "10010000000110100" => rgb <= "000000";
					when "10010000000110101" => rgb <= "000000";
					when "10010000000110110" => rgb <= "000000";
					when "10010000000110111" => rgb <= "000000";
					when "10010000000111000" => rgb <= "000000";
					when "10010000000111001" => rgb <= "000000";
					when "10010000000111010" => rgb <= "000000";
					when "10010000000111011" => rgb <= "000000";
					when "10010000000111100" => rgb <= "000000";
					when "10010000000111101" => rgb <= "000000";
					when "10010000000111110" => rgb <= "000000";
					when "10010000000111111" => rgb <= "000000";
					when "10010000001000000" => rgb <= "000000";
					when "10010000001000001" => rgb <= "000000";
					when "10010000001000010" => rgb <= "000000";
					when "10010000001000011" => rgb <= "000000";
					when "10010000001000100" => rgb <= "000000";
					when "10010000001000101" => rgb <= "000000";
					when "10010000001000110" => rgb <= "000000";
					when "10010000001000111" => rgb <= "000000";
					when "10010000001001000" => rgb <= "000000";
					when "10010000001001001" => rgb <= "000000";
					when "10010000001001010" => rgb <= "000000";
					when "10010000001001011" => rgb <= "000000";
					when "10010000001001100" => rgb <= "000000";
					when "10010000001001101" => rgb <= "000000";
					when "10010000001001110" => rgb <= "000000";
					when "10010000001001111" => rgb <= "000000";
					when "10010000001010000" => rgb <= "000000";
					when "10010000001010001" => rgb <= "000000";
					when "10010000001010010" => rgb <= "000000";
					when "10010000001010011" => rgb <= "000000";
					when "10010000001010100" => rgb <= "000000";
					when "10010000001010101" => rgb <= "000000";
					when "10010000001010110" => rgb <= "000000";
					when "10010000001010111" => rgb <= "000000";
					when "10010000001011000" => rgb <= "000000";
					when "10010000001011001" => rgb <= "000000";
					when "10010000001011010" => rgb <= "000000";
					when "10010000001011011" => rgb <= "000000";
					when "10010000001011100" => rgb <= "000000";
					when "10010000001011101" => rgb <= "000000";
					when "10010000001011110" => rgb <= "000000";
					when "10010000001011111" => rgb <= "000000";
					when "10010000001100000" => rgb <= "000000";
					when "10010000001100001" => rgb <= "000000";
					when "10010000001100010" => rgb <= "000000";
					when "10010000001100011" => rgb <= "000000";
					when "10010000001100100" => rgb <= "000000";
					when "10010000001100101" => rgb <= "000000";
					when "10010000001100110" => rgb <= "000000";
					when "10010000001100111" => rgb <= "000000";
					when "10010000001101000" => rgb <= "000000";
					when "10010000001101001" => rgb <= "000000";
					when "10010000001101010" => rgb <= "000000";
					when "10010000001101011" => rgb <= "000000";
					when "10010000001101100" => rgb <= "000000";
					when "10010000001101101" => rgb <= "000000";
					when "10010000001101110" => rgb <= "000000";
					when "10010000001101111" => rgb <= "000000";
					when "10010000001110000" => rgb <= "000000";
					when "10010000001110001" => rgb <= "000000";
					when "10010000001110010" => rgb <= "000000";
					when "10010000001110011" => rgb <= "000000";
					when "10010000001110100" => rgb <= "000000";
					when "10010000001110101" => rgb <= "000000";
					when "10010000001110110" => rgb <= "000000";
					when "10010000001110111" => rgb <= "000000";
					when "10010000001111000" => rgb <= "000000";
					when "10010000001111001" => rgb <= "000000";
					when "10010000001111010" => rgb <= "000000";
					when "10010000001111011" => rgb <= "000000";
					when "10010000001111100" => rgb <= "000000";
					when "10010000001111101" => rgb <= "000000";
					when "10010000001111110" => rgb <= "000000";
					when "10010000001111111" => rgb <= "000000";
					when "10010000010000000" => rgb <= "000000";
					when "10010000010000001" => rgb <= "000000";
					when "10010000010000010" => rgb <= "000000";
					when "10010000010000011" => rgb <= "000000";
					when "10010000010000100" => rgb <= "000000";
					when "10010000010000101" => rgb <= "000000";
					when "10010000010000110" => rgb <= "000000";
					when "10010000010000111" => rgb <= "000000";
					when "10010000010001000" => rgb <= "000000";
					when "10010000010001001" => rgb <= "000000";
					when "10010000010001010" => rgb <= "000000";
					when "10010000010001011" => rgb <= "000000";
					when "10010000010001100" => rgb <= "000000";
					when "10010000010001101" => rgb <= "000000";
					when "10010000010001110" => rgb <= "000000";
					when "10010000010001111" => rgb <= "000000";
					when "10010000010010000" => rgb <= "000000";
					when "10010000010010001" => rgb <= "000000";
					when "10010000010010010" => rgb <= "000000";
					when "10010000010010011" => rgb <= "000000";
					when "10010000010010100" => rgb <= "000000";
					when "10010000010010101" => rgb <= "000000";
					when "10010000010010110" => rgb <= "000000";
					when "10010000010010111" => rgb <= "000000";
					when "10010000010011000" => rgb <= "000000";
					when "10010000010011001" => rgb <= "000000";
					when "10010000010011010" => rgb <= "000000";
					when "10010000010011011" => rgb <= "000000";
					when "10010000010011100" => rgb <= "000000";
					when "10010000010011101" => rgb <= "000000";
					when "10010000010011110" => rgb <= "000000";
					when "10010000010011111" => rgb <= "000000";
					when "10010000010100000" => rgb <= "000000";
					when "10010000010100001" => rgb <= "000000";
					when "10010000010100010" => rgb <= "000000";
					when "10010000010100011" => rgb <= "000000";
					when "10010000010100100" => rgb <= "000000";
					when "10010000010100101" => rgb <= "000000";
					when "10010000010100110" => rgb <= "000000";
					when "10010000010100111" => rgb <= "000000";
					when "10010000010101000" => rgb <= "000000";
					when "10010000010101001" => rgb <= "000000";
					when "10010000010101010" => rgb <= "000000";
					when "10010000010101011" => rgb <= "000000";
					when "10010000010101100" => rgb <= "000000";
					when "10010000010101101" => rgb <= "000000";
					when "10010000010101110" => rgb <= "000000";
					when "10010000010101111" => rgb <= "000000";
					when "10010000010110000" => rgb <= "000000";
					when "10010000010110001" => rgb <= "000000";
					when "10010000010110010" => rgb <= "000000";
					when "10010000010110011" => rgb <= "000000";
					when "10010000010110100" => rgb <= "000000";
					when "10010000010110101" => rgb <= "000000";
					when "10010000010110110" => rgb <= "000000";
					when "10010000010110111" => rgb <= "000000";
					when "10010000010111000" => rgb <= "000000";
					when "10010000010111001" => rgb <= "000000";
					when "10010000010111010" => rgb <= "000000";
					when "10010000010111011" => rgb <= "000000";
					when "10010000010111100" => rgb <= "000000";
					when "10010000010111101" => rgb <= "000000";
					when "10010000010111110" => rgb <= "000000";
					when "10010000010111111" => rgb <= "000000";
					when "10010000011000000" => rgb <= "000000";
					when "10010000011000001" => rgb <= "000000";
					when "10010000011000010" => rgb <= "000000";
					when "10010000011000011" => rgb <= "000000";
					when "10010000011000100" => rgb <= "000000";
					when "10010000011000101" => rgb <= "000000";
					when "10010000011000110" => rgb <= "000000";
					when "10010000011000111" => rgb <= "000000";
					when "10010000011001000" => rgb <= "000000";
					when "10010000011001001" => rgb <= "000000";
					when "10010000011001010" => rgb <= "000000";
					when "10010000011001011" => rgb <= "000000";
					when "10010000011001100" => rgb <= "000000";
					when "10010000011001101" => rgb <= "000000";
					when "10010000011001110" => rgb <= "000000";
					when "10010000011001111" => rgb <= "000000";
					when "10010000011010000" => rgb <= "000000";
					when "10010000011010001" => rgb <= "000000";
					when "10010000011010010" => rgb <= "000000";
					when "10010000011010011" => rgb <= "000000";
					when "10010000011010100" => rgb <= "000000";
					when "10010000011010101" => rgb <= "000000";
					when "10010000011010110" => rgb <= "000000";
					when "10010000011010111" => rgb <= "000000";
					when "10010000011011000" => rgb <= "000000";
					when "10010000011011001" => rgb <= "000000";
					when "10010000011011010" => rgb <= "000000";
					when "10010000011011011" => rgb <= "000000";
					when "10010000011011100" => rgb <= "000000";
					when "10010000011011101" => rgb <= "000000";
					when "10010000011011110" => rgb <= "000000";
					when "10010000011011111" => rgb <= "000000";
					when "10010000011100000" => rgb <= "000000";
					when "10010000011100001" => rgb <= "000000";
					when "10010000011100010" => rgb <= "000000";
					when "10010000011100011" => rgb <= "000000";
					when "10010000011100100" => rgb <= "000000";
					when "10010000011100101" => rgb <= "000000";
					when "10010000011100110" => rgb <= "000000";
					when "10010000011100111" => rgb <= "000000";
					when "10010000011101000" => rgb <= "000000";
					when "10010000011101001" => rgb <= "000000";
					when "10010000011101010" => rgb <= "000000";
					when "10010000011101011" => rgb <= "000000";
					when "10010000011101100" => rgb <= "000000";
					when "10010000011101101" => rgb <= "000000";
					when "10010000011101110" => rgb <= "000000";
					when "10010000011101111" => rgb <= "000000";
					when "10010000011110000" => rgb <= "000000";
					when "10010000011110001" => rgb <= "000000";
					when "10010000011110010" => rgb <= "000000";
					when "10010000011110011" => rgb <= "000000";
					when "10010000011110100" => rgb <= "000000";
					when "10010000011110101" => rgb <= "000000";
					when "10010000011110110" => rgb <= "000000";
					when "10010000011110111" => rgb <= "000000";
					when "10010000011111000" => rgb <= "000000";
					when "10010000011111001" => rgb <= "000000";
					when "10010000011111010" => rgb <= "000000";
					when "10010000011111011" => rgb <= "000000";
					when "10010000011111100" => rgb <= "000000";
					when "10010000011111101" => rgb <= "000000";
					when "10010000011111110" => rgb <= "000000";
					when "10010000011111111" => rgb <= "000000";
					when "10010000100000000" => rgb <= "000000";
					when "10010000100000001" => rgb <= "000000";
					when "10010000100000010" => rgb <= "000000";
					when "10010000100000011" => rgb <= "000000";
					when "10010000100000100" => rgb <= "000000";
					when "10010000100000101" => rgb <= "000000";
					when "10010000100000110" => rgb <= "000000";
					when "10010000100000111" => rgb <= "000000";
					when "10010000100001000" => rgb <= "000000";
					when "10010000100001001" => rgb <= "000000";
					when "10010000100001010" => rgb <= "000000";
					when "10010000100001011" => rgb <= "000000";
					when "10010000100001100" => rgb <= "000000";
					when "10010000100001101" => rgb <= "000000";
					when "10010000100001110" => rgb <= "000000";
					when "10010000100001111" => rgb <= "000000";
					when "10010000100010000" => rgb <= "000000";
					when "10010000100010001" => rgb <= "000000";
					when "10010000100010010" => rgb <= "000000";
					when "10010000100010011" => rgb <= "000000";
					when "10010000100010100" => rgb <= "000000";
					when "10010000100010101" => rgb <= "000000";
					when "10010000100010110" => rgb <= "000000";
					when "10010000100010111" => rgb <= "000000";
					when "10010000100011000" => rgb <= "000000";
					when "10010000100011001" => rgb <= "000000";
					when "10010000100011010" => rgb <= "000000";
					when "10010000100011011" => rgb <= "000000";
					when "10010000100011100" => rgb <= "000000";
					when "10010000100011101" => rgb <= "000000";
					when "10010000100011110" => rgb <= "000000";
					when "10010000100011111" => rgb <= "000000";
					when "10010000100100000" => rgb <= "000000";
					when "10010000100100001" => rgb <= "000000";
					when "10010000100100010" => rgb <= "000000";
					when "10010000100100011" => rgb <= "000000";
					when "10010000100100100" => rgb <= "000000";
					when "10010000100100101" => rgb <= "000000";
					when "10010000100100110" => rgb <= "000000";
					when "10010000100100111" => rgb <= "000000";
					when "10010000100101000" => rgb <= "000000";
					when "10010000100101001" => rgb <= "000000";
					when "10010000100101010" => rgb <= "000000";
					when "10010000100101011" => rgb <= "000000";
					when "10010000100101100" => rgb <= "000000";
					when "10010000100101101" => rgb <= "000000";
					when "10010000100101110" => rgb <= "000000";
					when "10010000100101111" => rgb <= "000000";
					when "10010000100110000" => rgb <= "000000";
					when "10010000100110001" => rgb <= "000000";
					when "10010000100110010" => rgb <= "000000";
					when "10010000100110011" => rgb <= "000000";
					when "10010000100110100" => rgb <= "000000";
					when "10010000100110101" => rgb <= "000000";
					when "10010000100110110" => rgb <= "000000";
					when "10010000100110111" => rgb <= "000000";
					when "10010000100111000" => rgb <= "000000";
					when "10010000100111001" => rgb <= "000000";
					when "10010000100111010" => rgb <= "000000";
					when "10010000100111011" => rgb <= "000000";
					when "10010000100111100" => rgb <= "000000";
					when "10010000100111101" => rgb <= "000000";
					when "10010000100111110" => rgb <= "000000";
					when "10010000100111111" => rgb <= "000000";
					when "10010001000000000" => rgb <= "000000";
					when "10010001000000001" => rgb <= "000000";
					when "10010001000000010" => rgb <= "000000";
					when "10010001000000011" => rgb <= "000000";
					when "10010001000000100" => rgb <= "000000";
					when "10010001000000101" => rgb <= "000000";
					when "10010001000000110" => rgb <= "000000";
					when "10010001000000111" => rgb <= "000000";
					when "10010001000001000" => rgb <= "000000";
					when "10010001000001001" => rgb <= "000000";
					when "10010001000001010" => rgb <= "000000";
					when "10010001000001011" => rgb <= "000000";
					when "10010001000001100" => rgb <= "000000";
					when "10010001000001101" => rgb <= "000000";
					when "10010001000001110" => rgb <= "000000";
					when "10010001000001111" => rgb <= "000000";
					when "10010001000010000" => rgb <= "000000";
					when "10010001000010001" => rgb <= "000000";
					when "10010001000010010" => rgb <= "000000";
					when "10010001000010011" => rgb <= "000000";
					when "10010001000010100" => rgb <= "000000";
					when "10010001000010101" => rgb <= "000000";
					when "10010001000010110" => rgb <= "000000";
					when "10010001000010111" => rgb <= "000000";
					when "10010001000011000" => rgb <= "000000";
					when "10010001000011001" => rgb <= "000000";
					when "10010001000011010" => rgb <= "000000";
					when "10010001000011011" => rgb <= "000000";
					when "10010001000011100" => rgb <= "000000";
					when "10010001000011101" => rgb <= "000000";
					when "10010001000011110" => rgb <= "000000";
					when "10010001000011111" => rgb <= "000000";
					when "10010001000100000" => rgb <= "000000";
					when "10010001000100001" => rgb <= "000000";
					when "10010001000100010" => rgb <= "000000";
					when "10010001000100011" => rgb <= "000000";
					when "10010001000100100" => rgb <= "000000";
					when "10010001000100101" => rgb <= "000000";
					when "10010001000100110" => rgb <= "000000";
					when "10010001000100111" => rgb <= "000000";
					when "10010001000101000" => rgb <= "000000";
					when "10010001000101001" => rgb <= "000000";
					when "10010001000101010" => rgb <= "000000";
					when "10010001000101011" => rgb <= "000000";
					when "10010001000101100" => rgb <= "000000";
					when "10010001000101101" => rgb <= "000000";
					when "10010001000101110" => rgb <= "000000";
					when "10010001000101111" => rgb <= "000000";
					when "10010001000110000" => rgb <= "000000";
					when "10010001000110001" => rgb <= "000000";
					when "10010001000110010" => rgb <= "000000";
					when "10010001000110011" => rgb <= "000000";
					when "10010001000110100" => rgb <= "000000";
					when "10010001000110101" => rgb <= "000000";
					when "10010001000110110" => rgb <= "000000";
					when "10010001000110111" => rgb <= "000000";
					when "10010001000111000" => rgb <= "000000";
					when "10010001000111001" => rgb <= "000000";
					when "10010001000111010" => rgb <= "000000";
					when "10010001000111011" => rgb <= "000000";
					when "10010001000111100" => rgb <= "000000";
					when "10010001000111101" => rgb <= "000000";
					when "10010001000111110" => rgb <= "000000";
					when "10010001000111111" => rgb <= "000000";
					when "10010001001000000" => rgb <= "000000";
					when "10010001001000001" => rgb <= "000000";
					when "10010001001000010" => rgb <= "000000";
					when "10010001001000011" => rgb <= "000000";
					when "10010001001000100" => rgb <= "000000";
					when "10010001001000101" => rgb <= "000000";
					when "10010001001000110" => rgb <= "000000";
					when "10010001001000111" => rgb <= "000000";
					when "10010001001001000" => rgb <= "000000";
					when "10010001001001001" => rgb <= "000000";
					when "10010001001001010" => rgb <= "000000";
					when "10010001001001011" => rgb <= "000000";
					when "10010001001001100" => rgb <= "000000";
					when "10010001001001101" => rgb <= "000000";
					when "10010001001001110" => rgb <= "000000";
					when "10010001001001111" => rgb <= "000000";
					when "10010001001010000" => rgb <= "000000";
					when "10010001001010001" => rgb <= "000000";
					when "10010001001010010" => rgb <= "000000";
					when "10010001001010011" => rgb <= "000000";
					when "10010001001010100" => rgb <= "000000";
					when "10010001001010101" => rgb <= "000000";
					when "10010001001010110" => rgb <= "000000";
					when "10010001001010111" => rgb <= "000000";
					when "10010001001011000" => rgb <= "000000";
					when "10010001001011001" => rgb <= "000000";
					when "10010001001011010" => rgb <= "000000";
					when "10010001001011011" => rgb <= "000000";
					when "10010001001011100" => rgb <= "000000";
					when "10010001001011101" => rgb <= "000000";
					when "10010001001011110" => rgb <= "000000";
					when "10010001001011111" => rgb <= "000000";
					when "10010001001100000" => rgb <= "000000";
					when "10010001001100001" => rgb <= "000000";
					when "10010001001100010" => rgb <= "000000";
					when "10010001001100011" => rgb <= "000000";
					when "10010001001100100" => rgb <= "000000";
					when "10010001001100101" => rgb <= "000000";
					when "10010001001100110" => rgb <= "000000";
					when "10010001001100111" => rgb <= "000000";
					when "10010001001101000" => rgb <= "000000";
					when "10010001001101001" => rgb <= "000000";
					when "10010001001101010" => rgb <= "000000";
					when "10010001001101011" => rgb <= "000000";
					when "10010001001101100" => rgb <= "000000";
					when "10010001001101101" => rgb <= "000000";
					when "10010001001101110" => rgb <= "000000";
					when "10010001001101111" => rgb <= "000000";
					when "10010001001110000" => rgb <= "000000";
					when "10010001001110001" => rgb <= "000000";
					when "10010001001110010" => rgb <= "000000";
					when "10010001001110011" => rgb <= "000000";
					when "10010001001110100" => rgb <= "000000";
					when "10010001001110101" => rgb <= "000000";
					when "10010001001110110" => rgb <= "000000";
					when "10010001001110111" => rgb <= "000000";
					when "10010001001111000" => rgb <= "000000";
					when "10010001001111001" => rgb <= "000000";
					when "10010001001111010" => rgb <= "000000";
					when "10010001001111011" => rgb <= "000000";
					when "10010001001111100" => rgb <= "000000";
					when "10010001001111101" => rgb <= "000000";
					when "10010001001111110" => rgb <= "000000";
					when "10010001001111111" => rgb <= "000000";
					when "10010001010000000" => rgb <= "000000";
					when "10010001010000001" => rgb <= "000000";
					when "10010001010000010" => rgb <= "000000";
					when "10010001010000011" => rgb <= "000000";
					when "10010001010000100" => rgb <= "000000";
					when "10010001010000101" => rgb <= "000000";
					when "10010001010000110" => rgb <= "000000";
					when "10010001010000111" => rgb <= "000000";
					when "10010001010001000" => rgb <= "000000";
					when "10010001010001001" => rgb <= "000000";
					when "10010001010001010" => rgb <= "000000";
					when "10010001010001011" => rgb <= "000000";
					when "10010001010001100" => rgb <= "000000";
					when "10010001010001101" => rgb <= "000000";
					when "10010001010001110" => rgb <= "000000";
					when "10010001010001111" => rgb <= "000000";
					when "10010001010010000" => rgb <= "000000";
					when "10010001010010001" => rgb <= "000000";
					when "10010001010010010" => rgb <= "000000";
					when "10010001010010011" => rgb <= "000000";
					when "10010001010010100" => rgb <= "000000";
					when "10010001010010101" => rgb <= "000000";
					when "10010001010010110" => rgb <= "000000";
					when "10010001010010111" => rgb <= "000000";
					when "10010001010011000" => rgb <= "000000";
					when "10010001010011001" => rgb <= "000000";
					when "10010001010011010" => rgb <= "000000";
					when "10010001010011011" => rgb <= "000000";
					when "10010001010011100" => rgb <= "000000";
					when "10010001010011101" => rgb <= "000000";
					when "10010001010011110" => rgb <= "000000";
					when "10010001010011111" => rgb <= "000000";
					when "10010001010100000" => rgb <= "000000";
					when "10010001010100001" => rgb <= "000000";
					when "10010001010100010" => rgb <= "000000";
					when "10010001010100011" => rgb <= "000000";
					when "10010001010100100" => rgb <= "000000";
					when "10010001010100101" => rgb <= "000000";
					when "10010001010100110" => rgb <= "000000";
					when "10010001010100111" => rgb <= "000000";
					when "10010001010101000" => rgb <= "000000";
					when "10010001010101001" => rgb <= "000000";
					when "10010001010101010" => rgb <= "000000";
					when "10010001010101011" => rgb <= "000000";
					when "10010001010101100" => rgb <= "000000";
					when "10010001010101101" => rgb <= "000000";
					when "10010001010101110" => rgb <= "000000";
					when "10010001010101111" => rgb <= "000000";
					when "10010001010110000" => rgb <= "000000";
					when "10010001010110001" => rgb <= "000000";
					when "10010001010110010" => rgb <= "000000";
					when "10010001010110011" => rgb <= "000000";
					when "10010001010110100" => rgb <= "000000";
					when "10010001010110101" => rgb <= "000000";
					when "10010001010110110" => rgb <= "000000";
					when "10010001010110111" => rgb <= "000000";
					when "10010001010111000" => rgb <= "000000";
					when "10010001010111001" => rgb <= "000000";
					when "10010001010111010" => rgb <= "000000";
					when "10010001010111011" => rgb <= "000000";
					when "10010001010111100" => rgb <= "000000";
					when "10010001010111101" => rgb <= "000000";
					when "10010001010111110" => rgb <= "000000";
					when "10010001010111111" => rgb <= "000000";
					when "10010001011000000" => rgb <= "000000";
					when "10010001011000001" => rgb <= "000000";
					when "10010001011000010" => rgb <= "000000";
					when "10010001011000011" => rgb <= "000000";
					when "10010001011000100" => rgb <= "000000";
					when "10010001011000101" => rgb <= "000000";
					when "10010001011000110" => rgb <= "000000";
					when "10010001011000111" => rgb <= "000000";
					when "10010001011001000" => rgb <= "000000";
					when "10010001011001001" => rgb <= "000000";
					when "10010001011001010" => rgb <= "000000";
					when "10010001011001011" => rgb <= "000000";
					when "10010001011001100" => rgb <= "000000";
					when "10010001011001101" => rgb <= "000000";
					when "10010001011001110" => rgb <= "000000";
					when "10010001011001111" => rgb <= "000000";
					when "10010001011010000" => rgb <= "000000";
					when "10010001011010001" => rgb <= "000000";
					when "10010001011010010" => rgb <= "000000";
					when "10010001011010011" => rgb <= "000000";
					when "10010001011010100" => rgb <= "000000";
					when "10010001011010101" => rgb <= "000000";
					when "10010001011010110" => rgb <= "000000";
					when "10010001011010111" => rgb <= "000000";
					when "10010001011011000" => rgb <= "000000";
					when "10010001011011001" => rgb <= "000000";
					when "10010001011011010" => rgb <= "000000";
					when "10010001011011011" => rgb <= "000000";
					when "10010001011011100" => rgb <= "000000";
					when "10010001011011101" => rgb <= "000000";
					when "10010001011011110" => rgb <= "000000";
					when "10010001011011111" => rgb <= "000000";
					when "10010001011100000" => rgb <= "000000";
					when "10010001011100001" => rgb <= "000000";
					when "10010001011100010" => rgb <= "000000";
					when "10010001011100011" => rgb <= "000000";
					when "10010001011100100" => rgb <= "000000";
					when "10010001011100101" => rgb <= "000000";
					when "10010001011100110" => rgb <= "000000";
					when "10010001011100111" => rgb <= "000000";
					when "10010001011101000" => rgb <= "000000";
					when "10010001011101001" => rgb <= "000000";
					when "10010001011101010" => rgb <= "000000";
					when "10010001011101011" => rgb <= "000000";
					when "10010001011101100" => rgb <= "000000";
					when "10010001011101101" => rgb <= "000000";
					when "10010001011101110" => rgb <= "000000";
					when "10010001011101111" => rgb <= "000000";
					when "10010001011110000" => rgb <= "000000";
					when "10010001011110001" => rgb <= "000000";
					when "10010001011110010" => rgb <= "000000";
					when "10010001011110011" => rgb <= "000000";
					when "10010001011110100" => rgb <= "000000";
					when "10010001011110101" => rgb <= "000000";
					when "10010001011110110" => rgb <= "000000";
					when "10010001011110111" => rgb <= "000000";
					when "10010001011111000" => rgb <= "000000";
					when "10010001011111001" => rgb <= "000000";
					when "10010001011111010" => rgb <= "000000";
					when "10010001011111011" => rgb <= "000000";
					when "10010001011111100" => rgb <= "000000";
					when "10010001011111101" => rgb <= "000000";
					when "10010001011111110" => rgb <= "000000";
					when "10010001011111111" => rgb <= "000000";
					when "10010001100000000" => rgb <= "000000";
					when "10010001100000001" => rgb <= "000000";
					when "10010001100000010" => rgb <= "000000";
					when "10010001100000011" => rgb <= "000000";
					when "10010001100000100" => rgb <= "000000";
					when "10010001100000101" => rgb <= "000000";
					when "10010001100000110" => rgb <= "000000";
					when "10010001100000111" => rgb <= "000000";
					when "10010001100001000" => rgb <= "000000";
					when "10010001100001001" => rgb <= "000000";
					when "10010001100001010" => rgb <= "000000";
					when "10010001100001011" => rgb <= "000000";
					when "10010001100001100" => rgb <= "000000";
					when "10010001100001101" => rgb <= "000000";
					when "10010001100001110" => rgb <= "000000";
					when "10010001100001111" => rgb <= "000000";
					when "10010001100010000" => rgb <= "000000";
					when "10010001100010001" => rgb <= "000000";
					when "10010001100010010" => rgb <= "000000";
					when "10010001100010011" => rgb <= "000000";
					when "10010001100010100" => rgb <= "000000";
					when "10010001100010101" => rgb <= "000000";
					when "10010001100010110" => rgb <= "000000";
					when "10010001100010111" => rgb <= "000000";
					when "10010001100011000" => rgb <= "000000";
					when "10010001100011001" => rgb <= "000000";
					when "10010001100011010" => rgb <= "000000";
					when "10010001100011011" => rgb <= "000000";
					when "10010001100011100" => rgb <= "000000";
					when "10010001100011101" => rgb <= "000000";
					when "10010001100011110" => rgb <= "000000";
					when "10010001100011111" => rgb <= "000000";
					when "10010001100100000" => rgb <= "000000";
					when "10010001100100001" => rgb <= "000000";
					when "10010001100100010" => rgb <= "000000";
					when "10010001100100011" => rgb <= "000000";
					when "10010001100100100" => rgb <= "000000";
					when "10010001100100101" => rgb <= "000000";
					when "10010001100100110" => rgb <= "000000";
					when "10010001100100111" => rgb <= "000000";
					when "10010001100101000" => rgb <= "000000";
					when "10010001100101001" => rgb <= "000000";
					when "10010001100101010" => rgb <= "000000";
					when "10010001100101011" => rgb <= "000000";
					when "10010001100101100" => rgb <= "000000";
					when "10010001100101101" => rgb <= "000000";
					when "10010001100101110" => rgb <= "000000";
					when "10010001100101111" => rgb <= "000000";
					when "10010001100110000" => rgb <= "000000";
					when "10010001100110001" => rgb <= "000000";
					when "10010001100110010" => rgb <= "000000";
					when "10010001100110011" => rgb <= "000000";
					when "10010001100110100" => rgb <= "000000";
					when "10010001100110101" => rgb <= "000000";
					when "10010001100110110" => rgb <= "000000";
					when "10010001100110111" => rgb <= "000000";
					when "10010001100111000" => rgb <= "000000";
					when "10010001100111001" => rgb <= "000000";
					when "10010001100111010" => rgb <= "000000";
					when "10010001100111011" => rgb <= "000000";
					when "10010001100111100" => rgb <= "000000";
					when "10010001100111101" => rgb <= "000000";
					when "10010001100111110" => rgb <= "000000";
					when "10010001100111111" => rgb <= "000000";
					when "10010010000000000" => rgb <= "000000";
					when "10010010000000001" => rgb <= "000000";
					when "10010010000000010" => rgb <= "000000";
					when "10010010000000011" => rgb <= "000000";
					when "10010010000000100" => rgb <= "000000";
					when "10010010000000101" => rgb <= "000000";
					when "10010010000000110" => rgb <= "000000";
					when "10010010000000111" => rgb <= "000000";
					when "10010010000001000" => rgb <= "000000";
					when "10010010000001001" => rgb <= "000000";
					when "10010010000001010" => rgb <= "000000";
					when "10010010000001011" => rgb <= "000000";
					when "10010010000001100" => rgb <= "000000";
					when "10010010000001101" => rgb <= "000000";
					when "10010010000001110" => rgb <= "000000";
					when "10010010000001111" => rgb <= "000000";
					when "10010010000010000" => rgb <= "000000";
					when "10010010000010001" => rgb <= "000000";
					when "10010010000010010" => rgb <= "000000";
					when "10010010000010011" => rgb <= "000000";
					when "10010010000010100" => rgb <= "000000";
					when "10010010000010101" => rgb <= "000000";
					when "10010010000010110" => rgb <= "000000";
					when "10010010000010111" => rgb <= "000000";
					when "10010010000011000" => rgb <= "000000";
					when "10010010000011001" => rgb <= "000000";
					when "10010010000011010" => rgb <= "000000";
					when "10010010000011011" => rgb <= "000000";
					when "10010010000011100" => rgb <= "000000";
					when "10010010000011101" => rgb <= "000000";
					when "10010010000011110" => rgb <= "000000";
					when "10010010000011111" => rgb <= "000000";
					when "10010010000100000" => rgb <= "000000";
					when "10010010000100001" => rgb <= "000000";
					when "10010010000100010" => rgb <= "000000";
					when "10010010000100011" => rgb <= "000000";
					when "10010010000100100" => rgb <= "000000";
					when "10010010000100101" => rgb <= "000000";
					when "10010010000100110" => rgb <= "000000";
					when "10010010000100111" => rgb <= "000000";
					when "10010010000101000" => rgb <= "000000";
					when "10010010000101001" => rgb <= "000000";
					when "10010010000101010" => rgb <= "000000";
					when "10010010000101011" => rgb <= "000000";
					when "10010010000101100" => rgb <= "000000";
					when "10010010000101101" => rgb <= "000000";
					when "10010010000101110" => rgb <= "000000";
					when "10010010000101111" => rgb <= "000000";
					when "10010010000110000" => rgb <= "000000";
					when "10010010000110001" => rgb <= "000000";
					when "10010010000110010" => rgb <= "000000";
					when "10010010000110011" => rgb <= "000000";
					when "10010010000110100" => rgb <= "000000";
					when "10010010000110101" => rgb <= "000000";
					when "10010010000110110" => rgb <= "000000";
					when "10010010000110111" => rgb <= "000000";
					when "10010010000111000" => rgb <= "000000";
					when "10010010000111001" => rgb <= "000000";
					when "10010010000111010" => rgb <= "000000";
					when "10010010000111011" => rgb <= "000000";
					when "10010010000111100" => rgb <= "000000";
					when "10010010000111101" => rgb <= "000000";
					when "10010010000111110" => rgb <= "000000";
					when "10010010000111111" => rgb <= "000000";
					when "10010010001000000" => rgb <= "000000";
					when "10010010001000001" => rgb <= "000000";
					when "10010010001000010" => rgb <= "000000";
					when "10010010001000011" => rgb <= "000000";
					when "10010010001000100" => rgb <= "000000";
					when "10010010001000101" => rgb <= "000000";
					when "10010010001000110" => rgb <= "000000";
					when "10010010001000111" => rgb <= "000000";
					when "10010010001001000" => rgb <= "000000";
					when "10010010001001001" => rgb <= "000000";
					when "10010010001001010" => rgb <= "000000";
					when "10010010001001011" => rgb <= "000000";
					when "10010010001001100" => rgb <= "000000";
					when "10010010001001101" => rgb <= "000000";
					when "10010010001001110" => rgb <= "000000";
					when "10010010001001111" => rgb <= "000000";
					when "10010010001010000" => rgb <= "000000";
					when "10010010001010001" => rgb <= "000000";
					when "10010010001010010" => rgb <= "000000";
					when "10010010001010011" => rgb <= "000000";
					when "10010010001010100" => rgb <= "000000";
					when "10010010001010101" => rgb <= "000000";
					when "10010010001010110" => rgb <= "000000";
					when "10010010001010111" => rgb <= "000000";
					when "10010010001011000" => rgb <= "000000";
					when "10010010001011001" => rgb <= "000000";
					when "10010010001011010" => rgb <= "000000";
					when "10010010001011011" => rgb <= "000000";
					when "10010010001011100" => rgb <= "000000";
					when "10010010001011101" => rgb <= "000000";
					when "10010010001011110" => rgb <= "000000";
					when "10010010001011111" => rgb <= "000000";
					when "10010010001100000" => rgb <= "000000";
					when "10010010001100001" => rgb <= "000000";
					when "10010010001100010" => rgb <= "000000";
					when "10010010001100011" => rgb <= "000000";
					when "10010010001100100" => rgb <= "000000";
					when "10010010001100101" => rgb <= "000000";
					when "10010010001100110" => rgb <= "000000";
					when "10010010001100111" => rgb <= "000000";
					when "10010010001101000" => rgb <= "000000";
					when "10010010001101001" => rgb <= "000000";
					when "10010010001101010" => rgb <= "000000";
					when "10010010001101011" => rgb <= "000000";
					when "10010010001101100" => rgb <= "000000";
					when "10010010001101101" => rgb <= "000000";
					when "10010010001101110" => rgb <= "000000";
					when "10010010001101111" => rgb <= "000000";
					when "10010010001110000" => rgb <= "000000";
					when "10010010001110001" => rgb <= "000000";
					when "10010010001110010" => rgb <= "000000";
					when "10010010001110011" => rgb <= "000000";
					when "10010010001110100" => rgb <= "000000";
					when "10010010001110101" => rgb <= "000000";
					when "10010010001110110" => rgb <= "000000";
					when "10010010001110111" => rgb <= "000000";
					when "10010010001111000" => rgb <= "000000";
					when "10010010001111001" => rgb <= "000000";
					when "10010010001111010" => rgb <= "000000";
					when "10010010001111011" => rgb <= "000000";
					when "10010010001111100" => rgb <= "000000";
					when "10010010001111101" => rgb <= "000000";
					when "10010010001111110" => rgb <= "000000";
					when "10010010001111111" => rgb <= "000000";
					when "10010010010000000" => rgb <= "000000";
					when "10010010010000001" => rgb <= "000000";
					when "10010010010000010" => rgb <= "000000";
					when "10010010010000011" => rgb <= "000000";
					when "10010010010000100" => rgb <= "000000";
					when "10010010010000101" => rgb <= "000000";
					when "10010010010000110" => rgb <= "000000";
					when "10010010010000111" => rgb <= "000000";
					when "10010010010001000" => rgb <= "000000";
					when "10010010010001001" => rgb <= "000000";
					when "10010010010001010" => rgb <= "000000";
					when "10010010010001011" => rgb <= "000000";
					when "10010010010001100" => rgb <= "000000";
					when "10010010010001101" => rgb <= "000000";
					when "10010010010001110" => rgb <= "000000";
					when "10010010010001111" => rgb <= "000000";
					when "10010010010010000" => rgb <= "000000";
					when "10010010010010001" => rgb <= "000000";
					when "10010010010010010" => rgb <= "000000";
					when "10010010010010011" => rgb <= "000000";
					when "10010010010010100" => rgb <= "000000";
					when "10010010010010101" => rgb <= "000000";
					when "10010010010010110" => rgb <= "000000";
					when "10010010010010111" => rgb <= "000000";
					when "10010010010011000" => rgb <= "000000";
					when "10010010010011001" => rgb <= "000000";
					when "10010010010011010" => rgb <= "000000";
					when "10010010010011011" => rgb <= "000000";
					when "10010010010011100" => rgb <= "000000";
					when "10010010010011101" => rgb <= "000000";
					when "10010010010011110" => rgb <= "000000";
					when "10010010010011111" => rgb <= "000000";
					when "10010010010100000" => rgb <= "000000";
					when "10010010010100001" => rgb <= "000000";
					when "10010010010100010" => rgb <= "000000";
					when "10010010010100011" => rgb <= "000000";
					when "10010010010100100" => rgb <= "000000";
					when "10010010010100101" => rgb <= "000000";
					when "10010010010100110" => rgb <= "000000";
					when "10010010010100111" => rgb <= "000000";
					when "10010010010101000" => rgb <= "000000";
					when "10010010010101001" => rgb <= "000000";
					when "10010010010101010" => rgb <= "000000";
					when "10010010010101011" => rgb <= "000000";
					when "10010010010101100" => rgb <= "000000";
					when "10010010010101101" => rgb <= "000000";
					when "10010010010101110" => rgb <= "000000";
					when "10010010010101111" => rgb <= "000000";
					when "10010010010110000" => rgb <= "000000";
					when "10010010010110001" => rgb <= "000000";
					when "10010010010110010" => rgb <= "000000";
					when "10010010010110011" => rgb <= "000000";
					when "10010010010110100" => rgb <= "000000";
					when "10010010010110101" => rgb <= "000000";
					when "10010010010110110" => rgb <= "000000";
					when "10010010010110111" => rgb <= "000000";
					when "10010010010111000" => rgb <= "000000";
					when "10010010010111001" => rgb <= "000000";
					when "10010010010111010" => rgb <= "000000";
					when "10010010010111011" => rgb <= "000000";
					when "10010010010111100" => rgb <= "000000";
					when "10010010010111101" => rgb <= "000000";
					when "10010010010111110" => rgb <= "000000";
					when "10010010010111111" => rgb <= "000000";
					when "10010010011000000" => rgb <= "000000";
					when "10010010011000001" => rgb <= "000000";
					when "10010010011000010" => rgb <= "000000";
					when "10010010011000011" => rgb <= "000000";
					when "10010010011000100" => rgb <= "000000";
					when "10010010011000101" => rgb <= "000000";
					when "10010010011000110" => rgb <= "000000";
					when "10010010011000111" => rgb <= "000000";
					when "10010010011001000" => rgb <= "000000";
					when "10010010011001001" => rgb <= "000000";
					when "10010010011001010" => rgb <= "000000";
					when "10010010011001011" => rgb <= "000000";
					when "10010010011001100" => rgb <= "000000";
					when "10010010011001101" => rgb <= "000000";
					when "10010010011001110" => rgb <= "000000";
					when "10010010011001111" => rgb <= "000000";
					when "10010010011010000" => rgb <= "000000";
					when "10010010011010001" => rgb <= "000000";
					when "10010010011010010" => rgb <= "000000";
					when "10010010011010011" => rgb <= "000000";
					when "10010010011010100" => rgb <= "000000";
					when "10010010011010101" => rgb <= "000000";
					when "10010010011010110" => rgb <= "000000";
					when "10010010011010111" => rgb <= "000000";
					when "10010010011011000" => rgb <= "000000";
					when "10010010011011001" => rgb <= "000000";
					when "10010010011011010" => rgb <= "000000";
					when "10010010011011011" => rgb <= "000000";
					when "10010010011011100" => rgb <= "000000";
					when "10010010011011101" => rgb <= "000000";
					when "10010010011011110" => rgb <= "000000";
					when "10010010011011111" => rgb <= "000000";
					when "10010010011100000" => rgb <= "000000";
					when "10010010011100001" => rgb <= "000000";
					when "10010010011100010" => rgb <= "000000";
					when "10010010011100011" => rgb <= "000000";
					when "10010010011100100" => rgb <= "000000";
					when "10010010011100101" => rgb <= "000000";
					when "10010010011100110" => rgb <= "000000";
					when "10010010011100111" => rgb <= "000000";
					when "10010010011101000" => rgb <= "000000";
					when "10010010011101001" => rgb <= "000000";
					when "10010010011101010" => rgb <= "000000";
					when "10010010011101011" => rgb <= "000000";
					when "10010010011101100" => rgb <= "000000";
					when "10010010011101101" => rgb <= "000000";
					when "10010010011101110" => rgb <= "000000";
					when "10010010011101111" => rgb <= "000000";
					when "10010010011110000" => rgb <= "000000";
					when "10010010011110001" => rgb <= "000000";
					when "10010010011110010" => rgb <= "000000";
					when "10010010011110011" => rgb <= "000000";
					when "10010010011110100" => rgb <= "000000";
					when "10010010011110101" => rgb <= "000000";
					when "10010010011110110" => rgb <= "000000";
					when "10010010011110111" => rgb <= "000000";
					when "10010010011111000" => rgb <= "000000";
					when "10010010011111001" => rgb <= "000000";
					when "10010010011111010" => rgb <= "000000";
					when "10010010011111011" => rgb <= "000000";
					when "10010010011111100" => rgb <= "000000";
					when "10010010011111101" => rgb <= "000000";
					when "10010010011111110" => rgb <= "000000";
					when "10010010011111111" => rgb <= "000000";
					when "10010010100000000" => rgb <= "000000";
					when "10010010100000001" => rgb <= "000000";
					when "10010010100000010" => rgb <= "000000";
					when "10010010100000011" => rgb <= "000000";
					when "10010010100000100" => rgb <= "000000";
					when "10010010100000101" => rgb <= "000000";
					when "10010010100000110" => rgb <= "000000";
					when "10010010100000111" => rgb <= "000000";
					when "10010010100001000" => rgb <= "000000";
					when "10010010100001001" => rgb <= "000000";
					when "10010010100001010" => rgb <= "000000";
					when "10010010100001011" => rgb <= "000000";
					when "10010010100001100" => rgb <= "000000";
					when "10010010100001101" => rgb <= "000000";
					when "10010010100001110" => rgb <= "000000";
					when "10010010100001111" => rgb <= "000000";
					when "10010010100010000" => rgb <= "000000";
					when "10010010100010001" => rgb <= "000000";
					when "10010010100010010" => rgb <= "000000";
					when "10010010100010011" => rgb <= "000000";
					when "10010010100010100" => rgb <= "000000";
					when "10010010100010101" => rgb <= "000000";
					when "10010010100010110" => rgb <= "000000";
					when "10010010100010111" => rgb <= "000000";
					when "10010010100011000" => rgb <= "000000";
					when "10010010100011001" => rgb <= "000000";
					when "10010010100011010" => rgb <= "000000";
					when "10010010100011011" => rgb <= "000000";
					when "10010010100011100" => rgb <= "000000";
					when "10010010100011101" => rgb <= "000000";
					when "10010010100011110" => rgb <= "000000";
					when "10010010100011111" => rgb <= "000000";
					when "10010010100100000" => rgb <= "000000";
					when "10010010100100001" => rgb <= "000000";
					when "10010010100100010" => rgb <= "000000";
					when "10010010100100011" => rgb <= "000000";
					when "10010010100100100" => rgb <= "000000";
					when "10010010100100101" => rgb <= "000000";
					when "10010010100100110" => rgb <= "000000";
					when "10010010100100111" => rgb <= "000000";
					when "10010010100101000" => rgb <= "000000";
					when "10010010100101001" => rgb <= "000000";
					when "10010010100101010" => rgb <= "000000";
					when "10010010100101011" => rgb <= "000000";
					when "10010010100101100" => rgb <= "000000";
					when "10010010100101101" => rgb <= "000000";
					when "10010010100101110" => rgb <= "000000";
					when "10010010100101111" => rgb <= "000000";
					when "10010010100110000" => rgb <= "000000";
					when "10010010100110001" => rgb <= "000000";
					when "10010010100110010" => rgb <= "000000";
					when "10010010100110011" => rgb <= "000000";
					when "10010010100110100" => rgb <= "000000";
					when "10010010100110101" => rgb <= "000000";
					when "10010010100110110" => rgb <= "000000";
					when "10010010100110111" => rgb <= "000000";
					when "10010010100111000" => rgb <= "000000";
					when "10010010100111001" => rgb <= "000000";
					when "10010010100111010" => rgb <= "000000";
					when "10010010100111011" => rgb <= "000000";
					when "10010010100111100" => rgb <= "000000";
					when "10010010100111101" => rgb <= "000000";
					when "10010010100111110" => rgb <= "000000";
					when "10010010100111111" => rgb <= "000000";
					when "10010011000000000" => rgb <= "000000";
					when "10010011000000001" => rgb <= "000000";
					when "10010011000000010" => rgb <= "000000";
					when "10010011000000011" => rgb <= "000000";
					when "10010011000000100" => rgb <= "000000";
					when "10010011000000101" => rgb <= "000000";
					when "10010011000000110" => rgb <= "000000";
					when "10010011000000111" => rgb <= "000000";
					when "10010011000001000" => rgb <= "000000";
					when "10010011000001001" => rgb <= "000000";
					when "10010011000001010" => rgb <= "000000";
					when "10010011000001011" => rgb <= "000000";
					when "10010011000001100" => rgb <= "000000";
					when "10010011000001101" => rgb <= "000000";
					when "10010011000001110" => rgb <= "000000";
					when "10010011000001111" => rgb <= "000000";
					when "10010011000010000" => rgb <= "000000";
					when "10010011000010001" => rgb <= "000000";
					when "10010011000010010" => rgb <= "000000";
					when "10010011000010011" => rgb <= "000000";
					when "10010011000010100" => rgb <= "000000";
					when "10010011000010101" => rgb <= "000000";
					when "10010011000010110" => rgb <= "000000";
					when "10010011000010111" => rgb <= "000000";
					when "10010011000011000" => rgb <= "000000";
					when "10010011000011001" => rgb <= "000000";
					when "10010011000011010" => rgb <= "000000";
					when "10010011000011011" => rgb <= "000000";
					when "10010011000011100" => rgb <= "000000";
					when "10010011000011101" => rgb <= "000000";
					when "10010011000011110" => rgb <= "000000";
					when "10010011000011111" => rgb <= "000000";
					when "10010011000100000" => rgb <= "000000";
					when "10010011000100001" => rgb <= "000000";
					when "10010011000100010" => rgb <= "000000";
					when "10010011000100011" => rgb <= "000000";
					when "10010011000100100" => rgb <= "000000";
					when "10010011000100101" => rgb <= "000000";
					when "10010011000100110" => rgb <= "000000";
					when "10010011000100111" => rgb <= "000000";
					when "10010011000101000" => rgb <= "000000";
					when "10010011000101001" => rgb <= "000000";
					when "10010011000101010" => rgb <= "000000";
					when "10010011000101011" => rgb <= "000000";
					when "10010011000101100" => rgb <= "000000";
					when "10010011000101101" => rgb <= "000000";
					when "10010011000101110" => rgb <= "000000";
					when "10010011000101111" => rgb <= "000000";
					when "10010011000110000" => rgb <= "000000";
					when "10010011000110001" => rgb <= "000000";
					when "10010011000110010" => rgb <= "000000";
					when "10010011000110011" => rgb <= "000000";
					when "10010011000110100" => rgb <= "000000";
					when "10010011000110101" => rgb <= "000000";
					when "10010011000110110" => rgb <= "000000";
					when "10010011000110111" => rgb <= "000000";
					when "10010011000111000" => rgb <= "000000";
					when "10010011000111001" => rgb <= "000000";
					when "10010011000111010" => rgb <= "000000";
					when "10010011000111011" => rgb <= "000000";
					when "10010011000111100" => rgb <= "000000";
					when "10010011000111101" => rgb <= "000000";
					when "10010011000111110" => rgb <= "000000";
					when "10010011000111111" => rgb <= "000000";
					when "10010011001000000" => rgb <= "000000";
					when "10010011001000001" => rgb <= "000000";
					when "10010011001000010" => rgb <= "000000";
					when "10010011001000011" => rgb <= "000000";
					when "10010011001000100" => rgb <= "000000";
					when "10010011001000101" => rgb <= "000000";
					when "10010011001000110" => rgb <= "000000";
					when "10010011001000111" => rgb <= "000000";
					when "10010011001001000" => rgb <= "000000";
					when "10010011001001001" => rgb <= "000000";
					when "10010011001001010" => rgb <= "000000";
					when "10010011001001011" => rgb <= "000000";
					when "10010011001001100" => rgb <= "000000";
					when "10010011001001101" => rgb <= "000000";
					when "10010011001001110" => rgb <= "000000";
					when "10010011001001111" => rgb <= "000000";
					when "10010011001010000" => rgb <= "000000";
					when "10010011001010001" => rgb <= "000000";
					when "10010011001010010" => rgb <= "000000";
					when "10010011001010011" => rgb <= "000000";
					when "10010011001010100" => rgb <= "000000";
					when "10010011001010101" => rgb <= "000000";
					when "10010011001010110" => rgb <= "000000";
					when "10010011001010111" => rgb <= "000000";
					when "10010011001011000" => rgb <= "000000";
					when "10010011001011001" => rgb <= "000000";
					when "10010011001011010" => rgb <= "000000";
					when "10010011001011011" => rgb <= "000000";
					when "10010011001011100" => rgb <= "000000";
					when "10010011001011101" => rgb <= "000000";
					when "10010011001011110" => rgb <= "000000";
					when "10010011001011111" => rgb <= "000000";
					when "10010011001100000" => rgb <= "000000";
					when "10010011001100001" => rgb <= "000000";
					when "10010011001100010" => rgb <= "000000";
					when "10010011001100011" => rgb <= "000000";
					when "10010011001100100" => rgb <= "000000";
					when "10010011001100101" => rgb <= "000000";
					when "10010011001100110" => rgb <= "000000";
					when "10010011001100111" => rgb <= "000000";
					when "10010011001101000" => rgb <= "000000";
					when "10010011001101001" => rgb <= "000000";
					when "10010011001101010" => rgb <= "000000";
					when "10010011001101011" => rgb <= "000000";
					when "10010011001101100" => rgb <= "000000";
					when "10010011001101101" => rgb <= "000000";
					when "10010011001101110" => rgb <= "000000";
					when "10010011001101111" => rgb <= "000000";
					when "10010011001110000" => rgb <= "000000";
					when "10010011001110001" => rgb <= "000000";
					when "10010011001110010" => rgb <= "000000";
					when "10010011001110011" => rgb <= "000000";
					when "10010011001110100" => rgb <= "000000";
					when "10010011001110101" => rgb <= "000000";
					when "10010011001110110" => rgb <= "000000";
					when "10010011001110111" => rgb <= "000000";
					when "10010011001111000" => rgb <= "000000";
					when "10010011001111001" => rgb <= "000000";
					when "10010011001111010" => rgb <= "000000";
					when "10010011001111011" => rgb <= "000000";
					when "10010011001111100" => rgb <= "000000";
					when "10010011001111101" => rgb <= "000000";
					when "10010011001111110" => rgb <= "000000";
					when "10010011001111111" => rgb <= "000000";
					when "10010011010000000" => rgb <= "000000";
					when "10010011010000001" => rgb <= "000000";
					when "10010011010000010" => rgb <= "000000";
					when "10010011010000011" => rgb <= "000000";
					when "10010011010000100" => rgb <= "000000";
					when "10010011010000101" => rgb <= "000000";
					when "10010011010000110" => rgb <= "000000";
					when "10010011010000111" => rgb <= "000000";
					when "10010011010001000" => rgb <= "000000";
					when "10010011010001001" => rgb <= "000000";
					when "10010011010001010" => rgb <= "000000";
					when "10010011010001011" => rgb <= "000000";
					when "10010011010001100" => rgb <= "000000";
					when "10010011010001101" => rgb <= "000000";
					when "10010011010001110" => rgb <= "000000";
					when "10010011010001111" => rgb <= "000000";
					when "10010011010010000" => rgb <= "000000";
					when "10010011010010001" => rgb <= "000000";
					when "10010011010010010" => rgb <= "000000";
					when "10010011010010011" => rgb <= "000000";
					when "10010011010010100" => rgb <= "000000";
					when "10010011010010101" => rgb <= "000000";
					when "10010011010010110" => rgb <= "000000";
					when "10010011010010111" => rgb <= "000000";
					when "10010011010011000" => rgb <= "000000";
					when "10010011010011001" => rgb <= "000000";
					when "10010011010011010" => rgb <= "000000";
					when "10010011010011011" => rgb <= "000000";
					when "10010011010011100" => rgb <= "000000";
					when "10010011010011101" => rgb <= "000000";
					when "10010011010011110" => rgb <= "000000";
					when "10010011010011111" => rgb <= "000000";
					when "10010011010100000" => rgb <= "000000";
					when "10010011010100001" => rgb <= "000000";
					when "10010011010100010" => rgb <= "000000";
					when "10010011010100011" => rgb <= "000000";
					when "10010011010100100" => rgb <= "000000";
					when "10010011010100101" => rgb <= "000000";
					when "10010011010100110" => rgb <= "000000";
					when "10010011010100111" => rgb <= "000000";
					when "10010011010101000" => rgb <= "000000";
					when "10010011010101001" => rgb <= "000000";
					when "10010011010101010" => rgb <= "000000";
					when "10010011010101011" => rgb <= "000000";
					when "10010011010101100" => rgb <= "000000";
					when "10010011010101101" => rgb <= "000000";
					when "10010011010101110" => rgb <= "000000";
					when "10010011010101111" => rgb <= "000000";
					when "10010011010110000" => rgb <= "000000";
					when "10010011010110001" => rgb <= "000000";
					when "10010011010110010" => rgb <= "000000";
					when "10010011010110011" => rgb <= "000000";
					when "10010011010110100" => rgb <= "000000";
					when "10010011010110101" => rgb <= "000000";
					when "10010011010110110" => rgb <= "000000";
					when "10010011010110111" => rgb <= "000000";
					when "10010011010111000" => rgb <= "000000";
					when "10010011010111001" => rgb <= "000000";
					when "10010011010111010" => rgb <= "000000";
					when "10010011010111011" => rgb <= "000000";
					when "10010011010111100" => rgb <= "000000";
					when "10010011010111101" => rgb <= "000000";
					when "10010011010111110" => rgb <= "000000";
					when "10010011010111111" => rgb <= "000000";
					when "10010011011000000" => rgb <= "000000";
					when "10010011011000001" => rgb <= "000000";
					when "10010011011000010" => rgb <= "000000";
					when "10010011011000011" => rgb <= "000000";
					when "10010011011000100" => rgb <= "000000";
					when "10010011011000101" => rgb <= "000000";
					when "10010011011000110" => rgb <= "000000";
					when "10010011011000111" => rgb <= "000000";
					when "10010011011001000" => rgb <= "000000";
					when "10010011011001001" => rgb <= "000000";
					when "10010011011001010" => rgb <= "000000";
					when "10010011011001011" => rgb <= "000000";
					when "10010011011001100" => rgb <= "000000";
					when "10010011011001101" => rgb <= "000000";
					when "10010011011001110" => rgb <= "000000";
					when "10010011011001111" => rgb <= "000000";
					when "10010011011010000" => rgb <= "000000";
					when "10010011011010001" => rgb <= "000000";
					when "10010011011010010" => rgb <= "000000";
					when "10010011011010011" => rgb <= "000000";
					when "10010011011010100" => rgb <= "000000";
					when "10010011011010101" => rgb <= "000000";
					when "10010011011010110" => rgb <= "000000";
					when "10010011011010111" => rgb <= "000000";
					when "10010011011011000" => rgb <= "000000";
					when "10010011011011001" => rgb <= "000000";
					when "10010011011011010" => rgb <= "000000";
					when "10010011011011011" => rgb <= "000000";
					when "10010011011011100" => rgb <= "000000";
					when "10010011011011101" => rgb <= "000000";
					when "10010011011011110" => rgb <= "000000";
					when "10010011011011111" => rgb <= "000000";
					when "10010011011100000" => rgb <= "000000";
					when "10010011011100001" => rgb <= "000000";
					when "10010011011100010" => rgb <= "000000";
					when "10010011011100011" => rgb <= "000000";
					when "10010011011100100" => rgb <= "000000";
					when "10010011011100101" => rgb <= "000000";
					when "10010011011100110" => rgb <= "000000";
					when "10010011011100111" => rgb <= "000000";
					when "10010011011101000" => rgb <= "000000";
					when "10010011011101001" => rgb <= "000000";
					when "10010011011101010" => rgb <= "000000";
					when "10010011011101011" => rgb <= "000000";
					when "10010011011101100" => rgb <= "000000";
					when "10010011011101101" => rgb <= "000000";
					when "10010011011101110" => rgb <= "000000";
					when "10010011011101111" => rgb <= "000000";
					when "10010011011110000" => rgb <= "000000";
					when "10010011011110001" => rgb <= "000000";
					when "10010011011110010" => rgb <= "000000";
					when "10010011011110011" => rgb <= "000000";
					when "10010011011110100" => rgb <= "000000";
					when "10010011011110101" => rgb <= "000000";
					when "10010011011110110" => rgb <= "000000";
					when "10010011011110111" => rgb <= "000000";
					when "10010011011111000" => rgb <= "000000";
					when "10010011011111001" => rgb <= "000000";
					when "10010011011111010" => rgb <= "000000";
					when "10010011011111011" => rgb <= "000000";
					when "10010011011111100" => rgb <= "000000";
					when "10010011011111101" => rgb <= "000000";
					when "10010011011111110" => rgb <= "000000";
					when "10010011011111111" => rgb <= "000000";
					when "10010011100000000" => rgb <= "000000";
					when "10010011100000001" => rgb <= "000000";
					when "10010011100000010" => rgb <= "000000";
					when "10010011100000011" => rgb <= "000000";
					when "10010011100000100" => rgb <= "000000";
					when "10010011100000101" => rgb <= "000000";
					when "10010011100000110" => rgb <= "000000";
					when "10010011100000111" => rgb <= "000000";
					when "10010011100001000" => rgb <= "000000";
					when "10010011100001001" => rgb <= "000000";
					when "10010011100001010" => rgb <= "000000";
					when "10010011100001011" => rgb <= "000000";
					when "10010011100001100" => rgb <= "000000";
					when "10010011100001101" => rgb <= "000000";
					when "10010011100001110" => rgb <= "000000";
					when "10010011100001111" => rgb <= "000000";
					when "10010011100010000" => rgb <= "000000";
					when "10010011100010001" => rgb <= "000000";
					when "10010011100010010" => rgb <= "000000";
					when "10010011100010011" => rgb <= "000000";
					when "10010011100010100" => rgb <= "000000";
					when "10010011100010101" => rgb <= "000000";
					when "10010011100010110" => rgb <= "000000";
					when "10010011100010111" => rgb <= "000000";
					when "10010011100011000" => rgb <= "000000";
					when "10010011100011001" => rgb <= "000000";
					when "10010011100011010" => rgb <= "000000";
					when "10010011100011011" => rgb <= "000000";
					when "10010011100011100" => rgb <= "000000";
					when "10010011100011101" => rgb <= "000000";
					when "10010011100011110" => rgb <= "000000";
					when "10010011100011111" => rgb <= "000000";
					when "10010011100100000" => rgb <= "000000";
					when "10010011100100001" => rgb <= "000000";
					when "10010011100100010" => rgb <= "000000";
					when "10010011100100011" => rgb <= "000000";
					when "10010011100100100" => rgb <= "000000";
					when "10010011100100101" => rgb <= "000000";
					when "10010011100100110" => rgb <= "000000";
					when "10010011100100111" => rgb <= "000000";
					when "10010011100101000" => rgb <= "000000";
					when "10010011100101001" => rgb <= "000000";
					when "10010011100101010" => rgb <= "000000";
					when "10010011100101011" => rgb <= "000000";
					when "10010011100101100" => rgb <= "000000";
					when "10010011100101101" => rgb <= "000000";
					when "10010011100101110" => rgb <= "000000";
					when "10010011100101111" => rgb <= "000000";
					when "10010011100110000" => rgb <= "000000";
					when "10010011100110001" => rgb <= "000000";
					when "10010011100110010" => rgb <= "000000";
					when "10010011100110011" => rgb <= "000000";
					when "10010011100110100" => rgb <= "000000";
					when "10010011100110101" => rgb <= "000000";
					when "10010011100110110" => rgb <= "000000";
					when "10010011100110111" => rgb <= "000000";
					when "10010011100111000" => rgb <= "000000";
					when "10010011100111001" => rgb <= "000000";
					when "10010011100111010" => rgb <= "000000";
					when "10010011100111011" => rgb <= "000000";
					when "10010011100111100" => rgb <= "000000";
					when "10010011100111101" => rgb <= "000000";
					when "10010011100111110" => rgb <= "000000";
					when "10010011100111111" => rgb <= "000000";
					when "10010100000000000" => rgb <= "000000";
					when "10010100000000001" => rgb <= "000000";
					when "10010100000000010" => rgb <= "000000";
					when "10010100000000011" => rgb <= "000000";
					when "10010100000000100" => rgb <= "000000";
					when "10010100000000101" => rgb <= "000000";
					when "10010100000000110" => rgb <= "000000";
					when "10010100000000111" => rgb <= "000000";
					when "10010100000001000" => rgb <= "000000";
					when "10010100000001001" => rgb <= "000000";
					when "10010100000001010" => rgb <= "000000";
					when "10010100000001011" => rgb <= "000000";
					when "10010100000001100" => rgb <= "000000";
					when "10010100000001101" => rgb <= "000000";
					when "10010100000001110" => rgb <= "000000";
					when "10010100000001111" => rgb <= "000000";
					when "10010100000010000" => rgb <= "000000";
					when "10010100000010001" => rgb <= "000000";
					when "10010100000010010" => rgb <= "000000";
					when "10010100000010011" => rgb <= "000000";
					when "10010100000010100" => rgb <= "000000";
					when "10010100000010101" => rgb <= "000000";
					when "10010100000010110" => rgb <= "000000";
					when "10010100000010111" => rgb <= "000000";
					when "10010100000011000" => rgb <= "000000";
					when "10010100000011001" => rgb <= "000000";
					when "10010100000011010" => rgb <= "000000";
					when "10010100000011011" => rgb <= "000000";
					when "10010100000011100" => rgb <= "000000";
					when "10010100000011101" => rgb <= "000000";
					when "10010100000011110" => rgb <= "000000";
					when "10010100000011111" => rgb <= "000000";
					when "10010100000100000" => rgb <= "000000";
					when "10010100000100001" => rgb <= "000000";
					when "10010100000100010" => rgb <= "000000";
					when "10010100000100011" => rgb <= "000000";
					when "10010100000100100" => rgb <= "000000";
					when "10010100000100101" => rgb <= "000000";
					when "10010100000100110" => rgb <= "000000";
					when "10010100000100111" => rgb <= "000000";
					when "10010100000101000" => rgb <= "000000";
					when "10010100000101001" => rgb <= "000000";
					when "10010100000101010" => rgb <= "000000";
					when "10010100000101011" => rgb <= "000000";
					when "10010100000101100" => rgb <= "000000";
					when "10010100000101101" => rgb <= "000000";
					when "10010100000101110" => rgb <= "000000";
					when "10010100000101111" => rgb <= "000000";
					when "10010100000110000" => rgb <= "000000";
					when "10010100000110001" => rgb <= "000000";
					when "10010100000110010" => rgb <= "000000";
					when "10010100000110011" => rgb <= "000000";
					when "10010100000110100" => rgb <= "000000";
					when "10010100000110101" => rgb <= "000000";
					when "10010100000110110" => rgb <= "000000";
					when "10010100000110111" => rgb <= "000000";
					when "10010100000111000" => rgb <= "000000";
					when "10010100000111001" => rgb <= "000000";
					when "10010100000111010" => rgb <= "000000";
					when "10010100000111011" => rgb <= "000000";
					when "10010100000111100" => rgb <= "000000";
					when "10010100000111101" => rgb <= "000000";
					when "10010100000111110" => rgb <= "000000";
					when "10010100000111111" => rgb <= "000000";
					when "10010100001000000" => rgb <= "000000";
					when "10010100001000001" => rgb <= "000000";
					when "10010100001000010" => rgb <= "000000";
					when "10010100001000011" => rgb <= "000000";
					when "10010100001000100" => rgb <= "000000";
					when "10010100001000101" => rgb <= "000000";
					when "10010100001000110" => rgb <= "000000";
					when "10010100001000111" => rgb <= "000000";
					when "10010100001001000" => rgb <= "000000";
					when "10010100001001001" => rgb <= "000000";
					when "10010100001001010" => rgb <= "000000";
					when "10010100001001011" => rgb <= "000000";
					when "10010100001001100" => rgb <= "000000";
					when "10010100001001101" => rgb <= "000000";
					when "10010100001001110" => rgb <= "000000";
					when "10010100001001111" => rgb <= "000000";
					when "10010100001010000" => rgb <= "000000";
					when "10010100001010001" => rgb <= "000000";
					when "10010100001010010" => rgb <= "000000";
					when "10010100001010011" => rgb <= "000000";
					when "10010100001010100" => rgb <= "000000";
					when "10010100001010101" => rgb <= "000000";
					when "10010100001010110" => rgb <= "000000";
					when "10010100001010111" => rgb <= "000000";
					when "10010100001011000" => rgb <= "000000";
					when "10010100001011001" => rgb <= "000000";
					when "10010100001011010" => rgb <= "000000";
					when "10010100001011011" => rgb <= "000000";
					when "10010100001011100" => rgb <= "000000";
					when "10010100001011101" => rgb <= "000000";
					when "10010100001011110" => rgb <= "000000";
					when "10010100001011111" => rgb <= "000000";
					when "10010100001100000" => rgb <= "000000";
					when "10010100001100001" => rgb <= "000000";
					when "10010100001100010" => rgb <= "000000";
					when "10010100001100011" => rgb <= "000000";
					when "10010100001100100" => rgb <= "000000";
					when "10010100001100101" => rgb <= "000000";
					when "10010100001100110" => rgb <= "000000";
					when "10010100001100111" => rgb <= "000000";
					when "10010100001101000" => rgb <= "000000";
					when "10010100001101001" => rgb <= "000000";
					when "10010100001101010" => rgb <= "000000";
					when "10010100001101011" => rgb <= "000000";
					when "10010100001101100" => rgb <= "000000";
					when "10010100001101101" => rgb <= "000000";
					when "10010100001101110" => rgb <= "000000";
					when "10010100001101111" => rgb <= "000000";
					when "10010100001110000" => rgb <= "000000";
					when "10010100001110001" => rgb <= "000000";
					when "10010100001110010" => rgb <= "000000";
					when "10010100001110011" => rgb <= "000000";
					when "10010100001110100" => rgb <= "000000";
					when "10010100001110101" => rgb <= "000000";
					when "10010100001110110" => rgb <= "000000";
					when "10010100001110111" => rgb <= "000000";
					when "10010100001111000" => rgb <= "000000";
					when "10010100001111001" => rgb <= "000000";
					when "10010100001111010" => rgb <= "000000";
					when "10010100001111011" => rgb <= "000000";
					when "10010100001111100" => rgb <= "000000";
					when "10010100001111101" => rgb <= "000000";
					when "10010100001111110" => rgb <= "000000";
					when "10010100001111111" => rgb <= "000000";
					when "10010100010000000" => rgb <= "000000";
					when "10010100010000001" => rgb <= "000000";
					when "10010100010000010" => rgb <= "000000";
					when "10010100010000011" => rgb <= "000000";
					when "10010100010000100" => rgb <= "000000";
					when "10010100010000101" => rgb <= "000000";
					when "10010100010000110" => rgb <= "000000";
					when "10010100010000111" => rgb <= "000000";
					when "10010100010001000" => rgb <= "000000";
					when "10010100010001001" => rgb <= "000000";
					when "10010100010001010" => rgb <= "000000";
					when "10010100010001011" => rgb <= "000000";
					when "10010100010001100" => rgb <= "000000";
					when "10010100010001101" => rgb <= "000000";
					when "10010100010001110" => rgb <= "000000";
					when "10010100010001111" => rgb <= "000000";
					when "10010100010010000" => rgb <= "000000";
					when "10010100010010001" => rgb <= "000000";
					when "10010100010010010" => rgb <= "000000";
					when "10010100010010011" => rgb <= "000000";
					when "10010100010010100" => rgb <= "000000";
					when "10010100010010101" => rgb <= "000000";
					when "10010100010010110" => rgb <= "000000";
					when "10010100010010111" => rgb <= "000000";
					when "10010100010011000" => rgb <= "000000";
					when "10010100010011001" => rgb <= "000000";
					when "10010100010011010" => rgb <= "000000";
					when "10010100010011011" => rgb <= "000000";
					when "10010100010011100" => rgb <= "000000";
					when "10010100010011101" => rgb <= "000000";
					when "10010100010011110" => rgb <= "000000";
					when "10010100010011111" => rgb <= "000000";
					when "10010100010100000" => rgb <= "000000";
					when "10010100010100001" => rgb <= "000000";
					when "10010100010100010" => rgb <= "000000";
					when "10010100010100011" => rgb <= "000000";
					when "10010100010100100" => rgb <= "000000";
					when "10010100010100101" => rgb <= "000000";
					when "10010100010100110" => rgb <= "000000";
					when "10010100010100111" => rgb <= "000000";
					when "10010100010101000" => rgb <= "000000";
					when "10010100010101001" => rgb <= "000000";
					when "10010100010101010" => rgb <= "000000";
					when "10010100010101011" => rgb <= "000000";
					when "10010100010101100" => rgb <= "000000";
					when "10010100010101101" => rgb <= "000000";
					when "10010100010101110" => rgb <= "000000";
					when "10010100010101111" => rgb <= "000000";
					when "10010100010110000" => rgb <= "000000";
					when "10010100010110001" => rgb <= "000000";
					when "10010100010110010" => rgb <= "000000";
					when "10010100010110011" => rgb <= "000000";
					when "10010100010110100" => rgb <= "000000";
					when "10010100010110101" => rgb <= "000000";
					when "10010100010110110" => rgb <= "000000";
					when "10010100010110111" => rgb <= "000000";
					when "10010100010111000" => rgb <= "000000";
					when "10010100010111001" => rgb <= "000000";
					when "10010100010111010" => rgb <= "000000";
					when "10010100010111011" => rgb <= "000000";
					when "10010100010111100" => rgb <= "000000";
					when "10010100010111101" => rgb <= "000000";
					when "10010100010111110" => rgb <= "000000";
					when "10010100010111111" => rgb <= "000000";
					when "10010100011000000" => rgb <= "000000";
					when "10010100011000001" => rgb <= "000000";
					when "10010100011000010" => rgb <= "000000";
					when "10010100011000011" => rgb <= "000000";
					when "10010100011000100" => rgb <= "000000";
					when "10010100011000101" => rgb <= "000000";
					when "10010100011000110" => rgb <= "000000";
					when "10010100011000111" => rgb <= "000000";
					when "10010100011001000" => rgb <= "000000";
					when "10010100011001001" => rgb <= "000000";
					when "10010100011001010" => rgb <= "000000";
					when "10010100011001011" => rgb <= "000000";
					when "10010100011001100" => rgb <= "000000";
					when "10010100011001101" => rgb <= "000000";
					when "10010100011001110" => rgb <= "000000";
					when "10010100011001111" => rgb <= "000000";
					when "10010100011010000" => rgb <= "000000";
					when "10010100011010001" => rgb <= "000000";
					when "10010100011010010" => rgb <= "000000";
					when "10010100011010011" => rgb <= "000000";
					when "10010100011010100" => rgb <= "000000";
					when "10010100011010101" => rgb <= "000000";
					when "10010100011010110" => rgb <= "000000";
					when "10010100011010111" => rgb <= "000000";
					when "10010100011011000" => rgb <= "000000";
					when "10010100011011001" => rgb <= "000000";
					when "10010100011011010" => rgb <= "000000";
					when "10010100011011011" => rgb <= "000000";
					when "10010100011011100" => rgb <= "000000";
					when "10010100011011101" => rgb <= "000000";
					when "10010100011011110" => rgb <= "000000";
					when "10010100011011111" => rgb <= "000000";
					when "10010100011100000" => rgb <= "000000";
					when "10010100011100001" => rgb <= "000000";
					when "10010100011100010" => rgb <= "000000";
					when "10010100011100011" => rgb <= "000000";
					when "10010100011100100" => rgb <= "000000";
					when "10010100011100101" => rgb <= "000000";
					when "10010100011100110" => rgb <= "000000";
					when "10010100011100111" => rgb <= "000000";
					when "10010100011101000" => rgb <= "000000";
					when "10010100011101001" => rgb <= "000000";
					when "10010100011101010" => rgb <= "000000";
					when "10010100011101011" => rgb <= "000000";
					when "10010100011101100" => rgb <= "000000";
					when "10010100011101101" => rgb <= "000000";
					when "10010100011101110" => rgb <= "000000";
					when "10010100011101111" => rgb <= "000000";
					when "10010100011110000" => rgb <= "000000";
					when "10010100011110001" => rgb <= "000000";
					when "10010100011110010" => rgb <= "000000";
					when "10010100011110011" => rgb <= "000000";
					when "10010100011110100" => rgb <= "000000";
					when "10010100011110101" => rgb <= "000000";
					when "10010100011110110" => rgb <= "000000";
					when "10010100011110111" => rgb <= "000000";
					when "10010100011111000" => rgb <= "000000";
					when "10010100011111001" => rgb <= "000000";
					when "10010100011111010" => rgb <= "000000";
					when "10010100011111011" => rgb <= "000000";
					when "10010100011111100" => rgb <= "000000";
					when "10010100011111101" => rgb <= "000000";
					when "10010100011111110" => rgb <= "000000";
					when "10010100011111111" => rgb <= "000000";
					when "10010100100000000" => rgb <= "000000";
					when "10010100100000001" => rgb <= "000000";
					when "10010100100000010" => rgb <= "000000";
					when "10010100100000011" => rgb <= "000000";
					when "10010100100000100" => rgb <= "000000";
					when "10010100100000101" => rgb <= "000000";
					when "10010100100000110" => rgb <= "000000";
					when "10010100100000111" => rgb <= "000000";
					when "10010100100001000" => rgb <= "000000";
					when "10010100100001001" => rgb <= "000000";
					when "10010100100001010" => rgb <= "000000";
					when "10010100100001011" => rgb <= "000000";
					when "10010100100001100" => rgb <= "000000";
					when "10010100100001101" => rgb <= "000000";
					when "10010100100001110" => rgb <= "000000";
					when "10010100100001111" => rgb <= "000000";
					when "10010100100010000" => rgb <= "000000";
					when "10010100100010001" => rgb <= "000000";
					when "10010100100010010" => rgb <= "000000";
					when "10010100100010011" => rgb <= "000000";
					when "10010100100010100" => rgb <= "000000";
					when "10010100100010101" => rgb <= "000000";
					when "10010100100010110" => rgb <= "000000";
					when "10010100100010111" => rgb <= "000000";
					when "10010100100011000" => rgb <= "000000";
					when "10010100100011001" => rgb <= "000000";
					when "10010100100011010" => rgb <= "000000";
					when "10010100100011011" => rgb <= "000000";
					when "10010100100011100" => rgb <= "000000";
					when "10010100100011101" => rgb <= "000000";
					when "10010100100011110" => rgb <= "000000";
					when "10010100100011111" => rgb <= "000000";
					when "10010100100100000" => rgb <= "000000";
					when "10010100100100001" => rgb <= "000000";
					when "10010100100100010" => rgb <= "000000";
					when "10010100100100011" => rgb <= "000000";
					when "10010100100100100" => rgb <= "000000";
					when "10010100100100101" => rgb <= "000000";
					when "10010100100100110" => rgb <= "000000";
					when "10010100100100111" => rgb <= "000000";
					when "10010100100101000" => rgb <= "000000";
					when "10010100100101001" => rgb <= "000000";
					when "10010100100101010" => rgb <= "000000";
					when "10010100100101011" => rgb <= "000000";
					when "10010100100101100" => rgb <= "000000";
					when "10010100100101101" => rgb <= "000000";
					when "10010100100101110" => rgb <= "000000";
					when "10010100100101111" => rgb <= "000000";
					when "10010100100110000" => rgb <= "000000";
					when "10010100100110001" => rgb <= "000000";
					when "10010100100110010" => rgb <= "000000";
					when "10010100100110011" => rgb <= "000000";
					when "10010100100110100" => rgb <= "000000";
					when "10010100100110101" => rgb <= "000000";
					when "10010100100110110" => rgb <= "000000";
					when "10010100100110111" => rgb <= "000000";
					when "10010100100111000" => rgb <= "000000";
					when "10010100100111001" => rgb <= "000000";
					when "10010100100111010" => rgb <= "000000";
					when "10010100100111011" => rgb <= "000000";
					when "10010100100111100" => rgb <= "000000";
					when "10010100100111101" => rgb <= "000000";
					when "10010100100111110" => rgb <= "000000";
					when "10010100100111111" => rgb <= "000000";
					when "10010101000000000" => rgb <= "000000";
					when "10010101000000001" => rgb <= "000000";
					when "10010101000000010" => rgb <= "000000";
					when "10010101000000011" => rgb <= "000000";
					when "10010101000000100" => rgb <= "000000";
					when "10010101000000101" => rgb <= "000000";
					when "10010101000000110" => rgb <= "000000";
					when "10010101000000111" => rgb <= "000000";
					when "10010101000001000" => rgb <= "000000";
					when "10010101000001001" => rgb <= "000000";
					when "10010101000001010" => rgb <= "000000";
					when "10010101000001011" => rgb <= "000000";
					when "10010101000001100" => rgb <= "000000";
					when "10010101000001101" => rgb <= "000000";
					when "10010101000001110" => rgb <= "000000";
					when "10010101000001111" => rgb <= "000000";
					when "10010101000010000" => rgb <= "000000";
					when "10010101000010001" => rgb <= "000000";
					when "10010101000010010" => rgb <= "000000";
					when "10010101000010011" => rgb <= "000000";
					when "10010101000010100" => rgb <= "000000";
					when "10010101000010101" => rgb <= "000000";
					when "10010101000010110" => rgb <= "000000";
					when "10010101000010111" => rgb <= "000000";
					when "10010101000011000" => rgb <= "000000";
					when "10010101000011001" => rgb <= "000000";
					when "10010101000011010" => rgb <= "000000";
					when "10010101000011011" => rgb <= "000000";
					when "10010101000011100" => rgb <= "000000";
					when "10010101000011101" => rgb <= "000000";
					when "10010101000011110" => rgb <= "000000";
					when "10010101000011111" => rgb <= "000000";
					when "10010101000100000" => rgb <= "000000";
					when "10010101000100001" => rgb <= "000000";
					when "10010101000100010" => rgb <= "000000";
					when "10010101000100011" => rgb <= "000000";
					when "10010101000100100" => rgb <= "000000";
					when "10010101000100101" => rgb <= "000000";
					when "10010101000100110" => rgb <= "000000";
					when "10010101000100111" => rgb <= "000000";
					when "10010101000101000" => rgb <= "000000";
					when "10010101000101001" => rgb <= "000000";
					when "10010101000101010" => rgb <= "000000";
					when "10010101000101011" => rgb <= "000000";
					when "10010101000101100" => rgb <= "000000";
					when "10010101000101101" => rgb <= "000000";
					when "10010101000101110" => rgb <= "000000";
					when "10010101000101111" => rgb <= "000000";
					when "10010101000110000" => rgb <= "000000";
					when "10010101000110001" => rgb <= "000000";
					when "10010101000110010" => rgb <= "000000";
					when "10010101000110011" => rgb <= "000000";
					when "10010101000110100" => rgb <= "000000";
					when "10010101000110101" => rgb <= "000000";
					when "10010101000110110" => rgb <= "000000";
					when "10010101000110111" => rgb <= "000000";
					when "10010101000111000" => rgb <= "000000";
					when "10010101000111001" => rgb <= "000000";
					when "10010101000111010" => rgb <= "000000";
					when "10010101000111011" => rgb <= "000000";
					when "10010101000111100" => rgb <= "000000";
					when "10010101000111101" => rgb <= "000000";
					when "10010101000111110" => rgb <= "000000";
					when "10010101000111111" => rgb <= "000000";
					when "10010101001000000" => rgb <= "000000";
					when "10010101001000001" => rgb <= "000000";
					when "10010101001000010" => rgb <= "000000";
					when "10010101001000011" => rgb <= "000000";
					when "10010101001000100" => rgb <= "000000";
					when "10010101001000101" => rgb <= "000000";
					when "10010101001000110" => rgb <= "000000";
					when "10010101001000111" => rgb <= "000000";
					when "10010101001001000" => rgb <= "000000";
					when "10010101001001001" => rgb <= "000000";
					when "10010101001001010" => rgb <= "000000";
					when "10010101001001011" => rgb <= "000000";
					when "10010101001001100" => rgb <= "000000";
					when "10010101001001101" => rgb <= "000000";
					when "10010101001001110" => rgb <= "000000";
					when "10010101001001111" => rgb <= "000000";
					when "10010101001010000" => rgb <= "000000";
					when "10010101001010001" => rgb <= "000000";
					when "10010101001010010" => rgb <= "000000";
					when "10010101001010011" => rgb <= "000000";
					when "10010101001010100" => rgb <= "000000";
					when "10010101001010101" => rgb <= "000000";
					when "10010101001010110" => rgb <= "000000";
					when "10010101001010111" => rgb <= "000000";
					when "10010101001011000" => rgb <= "000000";
					when "10010101001011001" => rgb <= "000000";
					when "10010101001011010" => rgb <= "000000";
					when "10010101001011011" => rgb <= "000000";
					when "10010101001011100" => rgb <= "000000";
					when "10010101001011101" => rgb <= "000000";
					when "10010101001011110" => rgb <= "000000";
					when "10010101001011111" => rgb <= "000000";
					when "10010101001100000" => rgb <= "000000";
					when "10010101001100001" => rgb <= "000000";
					when "10010101001100010" => rgb <= "000000";
					when "10010101001100011" => rgb <= "000000";
					when "10010101001100100" => rgb <= "000000";
					when "10010101001100101" => rgb <= "000000";
					when "10010101001100110" => rgb <= "000000";
					when "10010101001100111" => rgb <= "000000";
					when "10010101001101000" => rgb <= "000000";
					when "10010101001101001" => rgb <= "000000";
					when "10010101001101010" => rgb <= "000000";
					when "10010101001101011" => rgb <= "000000";
					when "10010101001101100" => rgb <= "000000";
					when "10010101001101101" => rgb <= "000000";
					when "10010101001101110" => rgb <= "000000";
					when "10010101001101111" => rgb <= "000000";
					when "10010101001110000" => rgb <= "000000";
					when "10010101001110001" => rgb <= "000000";
					when "10010101001110010" => rgb <= "000000";
					when "10010101001110011" => rgb <= "000000";
					when "10010101001110100" => rgb <= "000000";
					when "10010101001110101" => rgb <= "000000";
					when "10010101001110110" => rgb <= "000000";
					when "10010101001110111" => rgb <= "000000";
					when "10010101001111000" => rgb <= "000000";
					when "10010101001111001" => rgb <= "000000";
					when "10010101001111010" => rgb <= "000000";
					when "10010101001111011" => rgb <= "000000";
					when "10010101001111100" => rgb <= "000000";
					when "10010101001111101" => rgb <= "000000";
					when "10010101001111110" => rgb <= "000000";
					when "10010101001111111" => rgb <= "000000";
					when "10010101010000000" => rgb <= "000000";
					when "10010101010000001" => rgb <= "000000";
					when "10010101010000010" => rgb <= "000000";
					when "10010101010000011" => rgb <= "000000";
					when "10010101010000100" => rgb <= "000000";
					when "10010101010000101" => rgb <= "000000";
					when "10010101010000110" => rgb <= "000000";
					when "10010101010000111" => rgb <= "000000";
					when "10010101010001000" => rgb <= "000000";
					when "10010101010001001" => rgb <= "000000";
					when "10010101010001010" => rgb <= "000000";
					when "10010101010001011" => rgb <= "000000";
					when "10010101010001100" => rgb <= "000000";
					when "10010101010001101" => rgb <= "000000";
					when "10010101010001110" => rgb <= "000000";
					when "10010101010001111" => rgb <= "000000";
					when "10010101010010000" => rgb <= "000000";
					when "10010101010010001" => rgb <= "000000";
					when "10010101010010010" => rgb <= "000000";
					when "10010101010010011" => rgb <= "000000";
					when "10010101010010100" => rgb <= "000000";
					when "10010101010010101" => rgb <= "000000";
					when "10010101010010110" => rgb <= "000000";
					when "10010101010010111" => rgb <= "000000";
					when "10010101010011000" => rgb <= "000000";
					when "10010101010011001" => rgb <= "000000";
					when "10010101010011010" => rgb <= "000000";
					when "10010101010011011" => rgb <= "000000";
					when "10010101010011100" => rgb <= "000000";
					when "10010101010011101" => rgb <= "000000";
					when "10010101010011110" => rgb <= "000000";
					when "10010101010011111" => rgb <= "000000";
					when "10010101010100000" => rgb <= "000000";
					when "10010101010100001" => rgb <= "000000";
					when "10010101010100010" => rgb <= "000000";
					when "10010101010100011" => rgb <= "000000";
					when "10010101010100100" => rgb <= "000000";
					when "10010101010100101" => rgb <= "000000";
					when "10010101010100110" => rgb <= "000000";
					when "10010101010100111" => rgb <= "000000";
					when "10010101010101000" => rgb <= "000000";
					when "10010101010101001" => rgb <= "000000";
					when "10010101010101010" => rgb <= "000000";
					when "10010101010101011" => rgb <= "000000";
					when "10010101010101100" => rgb <= "000000";
					when "10010101010101101" => rgb <= "000000";
					when "10010101010101110" => rgb <= "000000";
					when "10010101010101111" => rgb <= "000000";
					when "10010101010110000" => rgb <= "000000";
					when "10010101010110001" => rgb <= "000000";
					when "10010101010110010" => rgb <= "000000";
					when "10010101010110011" => rgb <= "000000";
					when "10010101010110100" => rgb <= "000000";
					when "10010101010110101" => rgb <= "000000";
					when "10010101010110110" => rgb <= "000000";
					when "10010101010110111" => rgb <= "000000";
					when "10010101010111000" => rgb <= "000000";
					when "10010101010111001" => rgb <= "000000";
					when "10010101010111010" => rgb <= "000000";
					when "10010101010111011" => rgb <= "000000";
					when "10010101010111100" => rgb <= "000000";
					when "10010101010111101" => rgb <= "000000";
					when "10010101010111110" => rgb <= "000000";
					when "10010101010111111" => rgb <= "000000";
					when "10010101011000000" => rgb <= "000000";
					when "10010101011000001" => rgb <= "000000";
					when "10010101011000010" => rgb <= "000000";
					when "10010101011000011" => rgb <= "000000";
					when "10010101011000100" => rgb <= "000000";
					when "10010101011000101" => rgb <= "000000";
					when "10010101011000110" => rgb <= "000000";
					when "10010101011000111" => rgb <= "000000";
					when "10010101011001000" => rgb <= "000000";
					when "10010101011001001" => rgb <= "000000";
					when "10010101011001010" => rgb <= "000000";
					when "10010101011001011" => rgb <= "000000";
					when "10010101011001100" => rgb <= "000000";
					when "10010101011001101" => rgb <= "000000";
					when "10010101011001110" => rgb <= "000000";
					when "10010101011001111" => rgb <= "000000";
					when "10010101011010000" => rgb <= "000000";
					when "10010101011010001" => rgb <= "000000";
					when "10010101011010010" => rgb <= "000000";
					when "10010101011010011" => rgb <= "000000";
					when "10010101011010100" => rgb <= "000000";
					when "10010101011010101" => rgb <= "000000";
					when "10010101011010110" => rgb <= "000000";
					when "10010101011010111" => rgb <= "000000";
					when "10010101011011000" => rgb <= "000000";
					when "10010101011011001" => rgb <= "000000";
					when "10010101011011010" => rgb <= "000000";
					when "10010101011011011" => rgb <= "000000";
					when "10010101011011100" => rgb <= "000000";
					when "10010101011011101" => rgb <= "000000";
					when "10010101011011110" => rgb <= "000000";
					when "10010101011011111" => rgb <= "000000";
					when "10010101011100000" => rgb <= "000000";
					when "10010101011100001" => rgb <= "000000";
					when "10010101011100010" => rgb <= "000000";
					when "10010101011100011" => rgb <= "000000";
					when "10010101011100100" => rgb <= "000000";
					when "10010101011100101" => rgb <= "000000";
					when "10010101011100110" => rgb <= "000000";
					when "10010101011100111" => rgb <= "000000";
					when "10010101011101000" => rgb <= "000000";
					when "10010101011101001" => rgb <= "000000";
					when "10010101011101010" => rgb <= "000000";
					when "10010101011101011" => rgb <= "000000";
					when "10010101011101100" => rgb <= "000000";
					when "10010101011101101" => rgb <= "000000";
					when "10010101011101110" => rgb <= "000000";
					when "10010101011101111" => rgb <= "000000";
					when "10010101011110000" => rgb <= "000000";
					when "10010101011110001" => rgb <= "000000";
					when "10010101011110010" => rgb <= "000000";
					when "10010101011110011" => rgb <= "000000";
					when "10010101011110100" => rgb <= "000000";
					when "10010101011110101" => rgb <= "000000";
					when "10010101011110110" => rgb <= "000000";
					when "10010101011110111" => rgb <= "000000";
					when "10010101011111000" => rgb <= "000000";
					when "10010101011111001" => rgb <= "000000";
					when "10010101011111010" => rgb <= "000000";
					when "10010101011111011" => rgb <= "000000";
					when "10010101011111100" => rgb <= "000000";
					when "10010101011111101" => rgb <= "000000";
					when "10010101011111110" => rgb <= "000000";
					when "10010101011111111" => rgb <= "000000";
					when "10010101100000000" => rgb <= "000000";
					when "10010101100000001" => rgb <= "000000";
					when "10010101100000010" => rgb <= "000000";
					when "10010101100000011" => rgb <= "000000";
					when "10010101100000100" => rgb <= "000000";
					when "10010101100000101" => rgb <= "000000";
					when "10010101100000110" => rgb <= "000000";
					when "10010101100000111" => rgb <= "000000";
					when "10010101100001000" => rgb <= "000000";
					when "10010101100001001" => rgb <= "000000";
					when "10010101100001010" => rgb <= "000000";
					when "10010101100001011" => rgb <= "000000";
					when "10010101100001100" => rgb <= "000000";
					when "10010101100001101" => rgb <= "000000";
					when "10010101100001110" => rgb <= "000000";
					when "10010101100001111" => rgb <= "000000";
					when "10010101100010000" => rgb <= "000000";
					when "10010101100010001" => rgb <= "000000";
					when "10010101100010010" => rgb <= "000000";
					when "10010101100010011" => rgb <= "000000";
					when "10010101100010100" => rgb <= "000000";
					when "10010101100010101" => rgb <= "000000";
					when "10010101100010110" => rgb <= "000000";
					when "10010101100010111" => rgb <= "000000";
					when "10010101100011000" => rgb <= "000000";
					when "10010101100011001" => rgb <= "000000";
					when "10010101100011010" => rgb <= "000000";
					when "10010101100011011" => rgb <= "000000";
					when "10010101100011100" => rgb <= "000000";
					when "10010101100011101" => rgb <= "000000";
					when "10010101100011110" => rgb <= "000000";
					when "10010101100011111" => rgb <= "000000";
					when "10010101100100000" => rgb <= "000000";
					when "10010101100100001" => rgb <= "000000";
					when "10010101100100010" => rgb <= "000000";
					when "10010101100100011" => rgb <= "000000";
					when "10010101100100100" => rgb <= "000000";
					when "10010101100100101" => rgb <= "000000";
					when "10010101100100110" => rgb <= "000000";
					when "10010101100100111" => rgb <= "000000";
					when "10010101100101000" => rgb <= "000000";
					when "10010101100101001" => rgb <= "000000";
					when "10010101100101010" => rgb <= "000000";
					when "10010101100101011" => rgb <= "000000";
					when "10010101100101100" => rgb <= "000000";
					when "10010101100101101" => rgb <= "000000";
					when "10010101100101110" => rgb <= "000000";
					when "10010101100101111" => rgb <= "000000";
					when "10010101100110000" => rgb <= "000000";
					when "10010101100110001" => rgb <= "000000";
					when "10010101100110010" => rgb <= "000000";
					when "10010101100110011" => rgb <= "000000";
					when "10010101100110100" => rgb <= "000000";
					when "10010101100110101" => rgb <= "000000";
					when "10010101100110110" => rgb <= "000000";
					when "10010101100110111" => rgb <= "000000";
					when "10010101100111000" => rgb <= "000000";
					when "10010101100111001" => rgb <= "000000";
					when "10010101100111010" => rgb <= "000000";
					when "10010101100111011" => rgb <= "000000";
					when "10010101100111100" => rgb <= "000000";
					when "10010101100111101" => rgb <= "000000";
					when "10010101100111110" => rgb <= "000000";
					when "10010101100111111" => rgb <= "000000";
					when "10010110000000000" => rgb <= "000000";
					when "10010110000000001" => rgb <= "000000";
					when "10010110000000010" => rgb <= "000000";
					when "10010110000000011" => rgb <= "000000";
					when "10010110000000100" => rgb <= "000000";
					when "10010110000000101" => rgb <= "000000";
					when "10010110000000110" => rgb <= "000000";
					when "10010110000000111" => rgb <= "000000";
					when "10010110000001000" => rgb <= "000000";
					when "10010110000001001" => rgb <= "000000";
					when "10010110000001010" => rgb <= "000000";
					when "10010110000001011" => rgb <= "000000";
					when "10010110000001100" => rgb <= "000000";
					when "10010110000001101" => rgb <= "000000";
					when "10010110000001110" => rgb <= "000000";
					when "10010110000001111" => rgb <= "000000";
					when "10010110000010000" => rgb <= "000000";
					when "10010110000010001" => rgb <= "000000";
					when "10010110000010010" => rgb <= "000000";
					when "10010110000010011" => rgb <= "000000";
					when "10010110000010100" => rgb <= "000000";
					when "10010110000010101" => rgb <= "000000";
					when "10010110000010110" => rgb <= "000000";
					when "10010110000010111" => rgb <= "000000";
					when "10010110000011000" => rgb <= "000000";
					when "10010110000011001" => rgb <= "000000";
					when "10010110000011010" => rgb <= "000000";
					when "10010110000011011" => rgb <= "000000";
					when "10010110000011100" => rgb <= "000000";
					when "10010110000011101" => rgb <= "000000";
					when "10010110000011110" => rgb <= "000000";
					when "10010110000011111" => rgb <= "000000";
					when "10010110000100000" => rgb <= "000000";
					when "10010110000100001" => rgb <= "000000";
					when "10010110000100010" => rgb <= "000000";
					when "10010110000100011" => rgb <= "000000";
					when "10010110000100100" => rgb <= "000000";
					when "10010110000100101" => rgb <= "000000";
					when "10010110000100110" => rgb <= "000000";
					when "10010110000100111" => rgb <= "000000";
					when "10010110000101000" => rgb <= "000000";
					when "10010110000101001" => rgb <= "000000";
					when "10010110000101010" => rgb <= "000000";
					when "10010110000101011" => rgb <= "000000";
					when "10010110000101100" => rgb <= "000000";
					when "10010110000101101" => rgb <= "000000";
					when "10010110000101110" => rgb <= "000000";
					when "10010110000101111" => rgb <= "000000";
					when "10010110000110000" => rgb <= "000000";
					when "10010110000110001" => rgb <= "000000";
					when "10010110000110010" => rgb <= "000000";
					when "10010110000110011" => rgb <= "000000";
					when "10010110000110100" => rgb <= "000000";
					when "10010110000110101" => rgb <= "000000";
					when "10010110000110110" => rgb <= "000000";
					when "10010110000110111" => rgb <= "000000";
					when "10010110000111000" => rgb <= "000000";
					when "10010110000111001" => rgb <= "000000";
					when "10010110000111010" => rgb <= "000000";
					when "10010110000111011" => rgb <= "000000";
					when "10010110000111100" => rgb <= "000000";
					when "10010110000111101" => rgb <= "000000";
					when "10010110000111110" => rgb <= "000000";
					when "10010110000111111" => rgb <= "000000";
					when "10010110001000000" => rgb <= "000000";
					when "10010110001000001" => rgb <= "000000";
					when "10010110001000010" => rgb <= "000000";
					when "10010110001000011" => rgb <= "000000";
					when "10010110001000100" => rgb <= "000000";
					when "10010110001000101" => rgb <= "000000";
					when "10010110001000110" => rgb <= "000000";
					when "10010110001000111" => rgb <= "000000";
					when "10010110001001000" => rgb <= "000000";
					when "10010110001001001" => rgb <= "000000";
					when "10010110001001010" => rgb <= "000000";
					when "10010110001001011" => rgb <= "000000";
					when "10010110001001100" => rgb <= "000000";
					when "10010110001001101" => rgb <= "000000";
					when "10010110001001110" => rgb <= "000000";
					when "10010110001001111" => rgb <= "000000";
					when "10010110001010000" => rgb <= "000000";
					when "10010110001010001" => rgb <= "000000";
					when "10010110001010010" => rgb <= "000000";
					when "10010110001010011" => rgb <= "000000";
					when "10010110001010100" => rgb <= "000000";
					when "10010110001010101" => rgb <= "000000";
					when "10010110001010110" => rgb <= "000000";
					when "10010110001010111" => rgb <= "000000";
					when "10010110001011000" => rgb <= "000000";
					when "10010110001011001" => rgb <= "000000";
					when "10010110001011010" => rgb <= "000000";
					when "10010110001011011" => rgb <= "000000";
					when "10010110001011100" => rgb <= "000000";
					when "10010110001011101" => rgb <= "000000";
					when "10010110001011110" => rgb <= "000000";
					when "10010110001011111" => rgb <= "000000";
					when "10010110001100000" => rgb <= "000000";
					when "10010110001100001" => rgb <= "000000";
					when "10010110001100010" => rgb <= "000000";
					when "10010110001100011" => rgb <= "000000";
					when "10010110001100100" => rgb <= "000000";
					when "10010110001100101" => rgb <= "000000";
					when "10010110001100110" => rgb <= "000000";
					when "10010110001100111" => rgb <= "000000";
					when "10010110001101000" => rgb <= "000000";
					when "10010110001101001" => rgb <= "000000";
					when "10010110001101010" => rgb <= "000000";
					when "10010110001101011" => rgb <= "000000";
					when "10010110001101100" => rgb <= "000000";
					when "10010110001101101" => rgb <= "000000";
					when "10010110001101110" => rgb <= "000000";
					when "10010110001101111" => rgb <= "000000";
					when "10010110001110000" => rgb <= "000000";
					when "10010110001110001" => rgb <= "000000";
					when "10010110001110010" => rgb <= "000000";
					when "10010110001110011" => rgb <= "000000";
					when "10010110001110100" => rgb <= "000000";
					when "10010110001110101" => rgb <= "000000";
					when "10010110001110110" => rgb <= "000000";
					when "10010110001110111" => rgb <= "000000";
					when "10010110001111000" => rgb <= "000000";
					when "10010110001111001" => rgb <= "000000";
					when "10010110001111010" => rgb <= "000000";
					when "10010110001111011" => rgb <= "000000";
					when "10010110001111100" => rgb <= "000000";
					when "10010110001111101" => rgb <= "000000";
					when "10010110001111110" => rgb <= "000000";
					when "10010110001111111" => rgb <= "000000";
					when "10010110010000000" => rgb <= "000000";
					when "10010110010000001" => rgb <= "000000";
					when "10010110010000010" => rgb <= "000000";
					when "10010110010000011" => rgb <= "000000";
					when "10010110010000100" => rgb <= "000000";
					when "10010110010000101" => rgb <= "000000";
					when "10010110010000110" => rgb <= "000000";
					when "10010110010000111" => rgb <= "000000";
					when "10010110010001000" => rgb <= "000000";
					when "10010110010001001" => rgb <= "000000";
					when "10010110010001010" => rgb <= "000000";
					when "10010110010001011" => rgb <= "000000";
					when "10010110010001100" => rgb <= "000000";
					when "10010110010001101" => rgb <= "000000";
					when "10010110010001110" => rgb <= "000000";
					when "10010110010001111" => rgb <= "000000";
					when "10010110010010000" => rgb <= "000000";
					when "10010110010010001" => rgb <= "000000";
					when "10010110010010010" => rgb <= "000000";
					when "10010110010010011" => rgb <= "000000";
					when "10010110010010100" => rgb <= "000000";
					when "10010110010010101" => rgb <= "000000";
					when "10010110010010110" => rgb <= "000000";
					when "10010110010010111" => rgb <= "000000";
					when "10010110010011000" => rgb <= "000000";
					when "10010110010011001" => rgb <= "000000";
					when "10010110010011010" => rgb <= "000000";
					when "10010110010011011" => rgb <= "000000";
					when "10010110010011100" => rgb <= "000000";
					when "10010110010011101" => rgb <= "000000";
					when "10010110010011110" => rgb <= "000000";
					when "10010110010011111" => rgb <= "000000";
					when "10010110010100000" => rgb <= "000000";
					when "10010110010100001" => rgb <= "000000";
					when "10010110010100010" => rgb <= "000000";
					when "10010110010100011" => rgb <= "000000";
					when "10010110010100100" => rgb <= "000000";
					when "10010110010100101" => rgb <= "000000";
					when "10010110010100110" => rgb <= "000000";
					when "10010110010100111" => rgb <= "000000";
					when "10010110010101000" => rgb <= "000000";
					when "10010110010101001" => rgb <= "000000";
					when "10010110010101010" => rgb <= "000000";
					when "10010110010101011" => rgb <= "000000";
					when "10010110010101100" => rgb <= "000000";
					when "10010110010101101" => rgb <= "000000";
					when "10010110010101110" => rgb <= "000000";
					when "10010110010101111" => rgb <= "000000";
					when "10010110010110000" => rgb <= "000000";
					when "10010110010110001" => rgb <= "000000";
					when "10010110010110010" => rgb <= "000000";
					when "10010110010110011" => rgb <= "000000";
					when "10010110010110100" => rgb <= "000000";
					when "10010110010110101" => rgb <= "000000";
					when "10010110010110110" => rgb <= "000000";
					when "10010110010110111" => rgb <= "000000";
					when "10010110010111000" => rgb <= "000000";
					when "10010110010111001" => rgb <= "000000";
					when "10010110010111010" => rgb <= "000000";
					when "10010110010111011" => rgb <= "000000";
					when "10010110010111100" => rgb <= "000000";
					when "10010110010111101" => rgb <= "000000";
					when "10010110010111110" => rgb <= "000000";
					when "10010110010111111" => rgb <= "000000";
					when "10010110011000000" => rgb <= "000000";
					when "10010110011000001" => rgb <= "000000";
					when "10010110011000010" => rgb <= "000000";
					when "10010110011000011" => rgb <= "000000";
					when "10010110011000100" => rgb <= "000000";
					when "10010110011000101" => rgb <= "000000";
					when "10010110011000110" => rgb <= "000000";
					when "10010110011000111" => rgb <= "000000";
					when "10010110011001000" => rgb <= "000000";
					when "10010110011001001" => rgb <= "000000";
					when "10010110011001010" => rgb <= "000000";
					when "10010110011001011" => rgb <= "000000";
					when "10010110011001100" => rgb <= "000000";
					when "10010110011001101" => rgb <= "000000";
					when "10010110011001110" => rgb <= "000000";
					when "10010110011001111" => rgb <= "000000";
					when "10010110011010000" => rgb <= "000000";
					when "10010110011010001" => rgb <= "000000";
					when "10010110011010010" => rgb <= "000000";
					when "10010110011010011" => rgb <= "000000";
					when "10010110011010100" => rgb <= "000000";
					when "10010110011010101" => rgb <= "000000";
					when "10010110011010110" => rgb <= "000000";
					when "10010110011010111" => rgb <= "000000";
					when "10010110011011000" => rgb <= "000000";
					when "10010110011011001" => rgb <= "000000";
					when "10010110011011010" => rgb <= "000000";
					when "10010110011011011" => rgb <= "000000";
					when "10010110011011100" => rgb <= "000000";
					when "10010110011011101" => rgb <= "000000";
					when "10010110011011110" => rgb <= "000000";
					when "10010110011011111" => rgb <= "000000";
					when "10010110011100000" => rgb <= "000000";
					when "10010110011100001" => rgb <= "000000";
					when "10010110011100010" => rgb <= "000000";
					when "10010110011100011" => rgb <= "000000";
					when "10010110011100100" => rgb <= "000000";
					when "10010110011100101" => rgb <= "000000";
					when "10010110011100110" => rgb <= "000000";
					when "10010110011100111" => rgb <= "000000";
					when "10010110011101000" => rgb <= "000000";
					when "10010110011101001" => rgb <= "000000";
					when "10010110011101010" => rgb <= "000000";
					when "10010110011101011" => rgb <= "000000";
					when "10010110011101100" => rgb <= "000000";
					when "10010110011101101" => rgb <= "000000";
					when "10010110011101110" => rgb <= "000000";
					when "10010110011101111" => rgb <= "000000";
					when "10010110011110000" => rgb <= "000000";
					when "10010110011110001" => rgb <= "000000";
					when "10010110011110010" => rgb <= "000000";
					when "10010110011110011" => rgb <= "000000";
					when "10010110011110100" => rgb <= "000000";
					when "10010110011110101" => rgb <= "000000";
					when "10010110011110110" => rgb <= "000000";
					when "10010110011110111" => rgb <= "000000";
					when "10010110011111000" => rgb <= "000000";
					when "10010110011111001" => rgb <= "000000";
					when "10010110011111010" => rgb <= "000000";
					when "10010110011111011" => rgb <= "000000";
					when "10010110011111100" => rgb <= "000000";
					when "10010110011111101" => rgb <= "000000";
					when "10010110011111110" => rgb <= "000000";
					when "10010110011111111" => rgb <= "000000";
					when "10010110100000000" => rgb <= "000000";
					when "10010110100000001" => rgb <= "000000";
					when "10010110100000010" => rgb <= "000000";
					when "10010110100000011" => rgb <= "000000";
					when "10010110100000100" => rgb <= "000000";
					when "10010110100000101" => rgb <= "000000";
					when "10010110100000110" => rgb <= "000000";
					when "10010110100000111" => rgb <= "000000";
					when "10010110100001000" => rgb <= "000000";
					when "10010110100001001" => rgb <= "000000";
					when "10010110100001010" => rgb <= "000000";
					when "10010110100001011" => rgb <= "000000";
					when "10010110100001100" => rgb <= "000000";
					when "10010110100001101" => rgb <= "000000";
					when "10010110100001110" => rgb <= "000000";
					when "10010110100001111" => rgb <= "000000";
					when "10010110100010000" => rgb <= "000000";
					when "10010110100010001" => rgb <= "000000";
					when "10010110100010010" => rgb <= "000000";
					when "10010110100010011" => rgb <= "000000";
					when "10010110100010100" => rgb <= "000000";
					when "10010110100010101" => rgb <= "000000";
					when "10010110100010110" => rgb <= "000000";
					when "10010110100010111" => rgb <= "000000";
					when "10010110100011000" => rgb <= "000000";
					when "10010110100011001" => rgb <= "000000";
					when "10010110100011010" => rgb <= "000000";
					when "10010110100011011" => rgb <= "000000";
					when "10010110100011100" => rgb <= "000000";
					when "10010110100011101" => rgb <= "000000";
					when "10010110100011110" => rgb <= "000000";
					when "10010110100011111" => rgb <= "000000";
					when "10010110100100000" => rgb <= "000000";
					when "10010110100100001" => rgb <= "000000";
					when "10010110100100010" => rgb <= "000000";
					when "10010110100100011" => rgb <= "000000";
					when "10010110100100100" => rgb <= "000000";
					when "10010110100100101" => rgb <= "000000";
					when "10010110100100110" => rgb <= "000000";
					when "10010110100100111" => rgb <= "000000";
					when "10010110100101000" => rgb <= "000000";
					when "10010110100101001" => rgb <= "000000";
					when "10010110100101010" => rgb <= "000000";
					when "10010110100101011" => rgb <= "000000";
					when "10010110100101100" => rgb <= "000000";
					when "10010110100101101" => rgb <= "000000";
					when "10010110100101110" => rgb <= "000000";
					when "10010110100101111" => rgb <= "000000";
					when "10010110100110000" => rgb <= "000000";
					when "10010110100110001" => rgb <= "000000";
					when "10010110100110010" => rgb <= "000000";
					when "10010110100110011" => rgb <= "000000";
					when "10010110100110100" => rgb <= "000000";
					when "10010110100110101" => rgb <= "000000";
					when "10010110100110110" => rgb <= "000000";
					when "10010110100110111" => rgb <= "000000";
					when "10010110100111000" => rgb <= "000000";
					when "10010110100111001" => rgb <= "000000";
					when "10010110100111010" => rgb <= "000000";
					when "10010110100111011" => rgb <= "000000";
					when "10010110100111100" => rgb <= "000000";
					when "10010110100111101" => rgb <= "000000";
					when "10010110100111110" => rgb <= "000000";
					when "10010110100111111" => rgb <= "000000";
					when "10010111000000000" => rgb <= "000000";
					when "10010111000000001" => rgb <= "000000";
					when "10010111000000010" => rgb <= "000000";
					when "10010111000000011" => rgb <= "000000";
					when "10010111000000100" => rgb <= "000000";
					when "10010111000000101" => rgb <= "000000";
					when "10010111000000110" => rgb <= "000000";
					when "10010111000000111" => rgb <= "000000";
					when "10010111000001000" => rgb <= "000000";
					when "10010111000001001" => rgb <= "000000";
					when "10010111000001010" => rgb <= "000000";
					when "10010111000001011" => rgb <= "000000";
					when "10010111000001100" => rgb <= "000000";
					when "10010111000001101" => rgb <= "000000";
					when "10010111000001110" => rgb <= "000000";
					when "10010111000001111" => rgb <= "000000";
					when "10010111000010000" => rgb <= "000000";
					when "10010111000010001" => rgb <= "000000";
					when "10010111000010010" => rgb <= "000000";
					when "10010111000010011" => rgb <= "000000";
					when "10010111000010100" => rgb <= "000000";
					when "10010111000010101" => rgb <= "000000";
					when "10010111000010110" => rgb <= "000000";
					when "10010111000010111" => rgb <= "000000";
					when "10010111000011000" => rgb <= "000000";
					when "10010111000011001" => rgb <= "000000";
					when "10010111000011010" => rgb <= "000000";
					when "10010111000011011" => rgb <= "000000";
					when "10010111000011100" => rgb <= "000000";
					when "10010111000011101" => rgb <= "000000";
					when "10010111000011110" => rgb <= "000000";
					when "10010111000011111" => rgb <= "000000";
					when "10010111000100000" => rgb <= "000000";
					when "10010111000100001" => rgb <= "000000";
					when "10010111000100010" => rgb <= "000000";
					when "10010111000100011" => rgb <= "000000";
					when "10010111000100100" => rgb <= "000000";
					when "10010111000100101" => rgb <= "000000";
					when "10010111000100110" => rgb <= "000000";
					when "10010111000100111" => rgb <= "000000";
					when "10010111000101000" => rgb <= "000000";
					when "10010111000101001" => rgb <= "000000";
					when "10010111000101010" => rgb <= "000000";
					when "10010111000101011" => rgb <= "000000";
					when "10010111000101100" => rgb <= "000000";
					when "10010111000101101" => rgb <= "000000";
					when "10010111000101110" => rgb <= "000000";
					when "10010111000101111" => rgb <= "000000";
					when "10010111000110000" => rgb <= "000000";
					when "10010111000110001" => rgb <= "000000";
					when "10010111000110010" => rgb <= "000000";
					when "10010111000110011" => rgb <= "000000";
					when "10010111000110100" => rgb <= "000000";
					when "10010111000110101" => rgb <= "000000";
					when "10010111000110110" => rgb <= "000000";
					when "10010111000110111" => rgb <= "000000";
					when "10010111000111000" => rgb <= "000000";
					when "10010111000111001" => rgb <= "000000";
					when "10010111000111010" => rgb <= "000000";
					when "10010111000111011" => rgb <= "000000";
					when "10010111000111100" => rgb <= "000000";
					when "10010111000111101" => rgb <= "000000";
					when "10010111000111110" => rgb <= "000000";
					when "10010111000111111" => rgb <= "000000";
					when "10010111001000000" => rgb <= "000000";
					when "10010111001000001" => rgb <= "000000";
					when "10010111001000010" => rgb <= "000000";
					when "10010111001000011" => rgb <= "000000";
					when "10010111001000100" => rgb <= "000000";
					when "10010111001000101" => rgb <= "000000";
					when "10010111001000110" => rgb <= "000000";
					when "10010111001000111" => rgb <= "000000";
					when "10010111001001000" => rgb <= "000000";
					when "10010111001001001" => rgb <= "000000";
					when "10010111001001010" => rgb <= "000000";
					when "10010111001001011" => rgb <= "000000";
					when "10010111001001100" => rgb <= "000000";
					when "10010111001001101" => rgb <= "000000";
					when "10010111001001110" => rgb <= "000000";
					when "10010111001001111" => rgb <= "000000";
					when "10010111001010000" => rgb <= "000000";
					when "10010111001010001" => rgb <= "000000";
					when "10010111001010010" => rgb <= "000000";
					when "10010111001010011" => rgb <= "000000";
					when "10010111001010100" => rgb <= "000000";
					when "10010111001010101" => rgb <= "000000";
					when "10010111001010110" => rgb <= "000000";
					when "10010111001010111" => rgb <= "000000";
					when "10010111001011000" => rgb <= "000000";
					when "10010111001011001" => rgb <= "000000";
					when "10010111001011010" => rgb <= "000000";
					when "10010111001011011" => rgb <= "000000";
					when "10010111001011100" => rgb <= "000000";
					when "10010111001011101" => rgb <= "000000";
					when "10010111001011110" => rgb <= "000000";
					when "10010111001011111" => rgb <= "000000";
					when "10010111001100000" => rgb <= "000000";
					when "10010111001100001" => rgb <= "000000";
					when "10010111001100010" => rgb <= "000000";
					when "10010111001100011" => rgb <= "000000";
					when "10010111001100100" => rgb <= "000000";
					when "10010111001100101" => rgb <= "000000";
					when "10010111001100110" => rgb <= "000000";
					when "10010111001100111" => rgb <= "000000";
					when "10010111001101000" => rgb <= "000000";
					when "10010111001101001" => rgb <= "000000";
					when "10010111001101010" => rgb <= "000000";
					when "10010111001101011" => rgb <= "000000";
					when "10010111001101100" => rgb <= "000000";
					when "10010111001101101" => rgb <= "000000";
					when "10010111001101110" => rgb <= "000000";
					when "10010111001101111" => rgb <= "000000";
					when "10010111001110000" => rgb <= "000000";
					when "10010111001110001" => rgb <= "000000";
					when "10010111001110010" => rgb <= "000000";
					when "10010111001110011" => rgb <= "000000";
					when "10010111001110100" => rgb <= "000000";
					when "10010111001110101" => rgb <= "000000";
					when "10010111001110110" => rgb <= "000000";
					when "10010111001110111" => rgb <= "000000";
					when "10010111001111000" => rgb <= "000000";
					when "10010111001111001" => rgb <= "000000";
					when "10010111001111010" => rgb <= "000000";
					when "10010111001111011" => rgb <= "000000";
					when "10010111001111100" => rgb <= "000000";
					when "10010111001111101" => rgb <= "000000";
					when "10010111001111110" => rgb <= "000000";
					when "10010111001111111" => rgb <= "000000";
					when "10010111010000000" => rgb <= "000000";
					when "10010111010000001" => rgb <= "000000";
					when "10010111010000010" => rgb <= "000000";
					when "10010111010000011" => rgb <= "000000";
					when "10010111010000100" => rgb <= "000000";
					when "10010111010000101" => rgb <= "000000";
					when "10010111010000110" => rgb <= "000000";
					when "10010111010000111" => rgb <= "000000";
					when "10010111010001000" => rgb <= "000000";
					when "10010111010001001" => rgb <= "000000";
					when "10010111010001010" => rgb <= "000000";
					when "10010111010001011" => rgb <= "000000";
					when "10010111010001100" => rgb <= "000000";
					when "10010111010001101" => rgb <= "000000";
					when "10010111010001110" => rgb <= "000000";
					when "10010111010001111" => rgb <= "000000";
					when "10010111010010000" => rgb <= "000000";
					when "10010111010010001" => rgb <= "000000";
					when "10010111010010010" => rgb <= "000000";
					when "10010111010010011" => rgb <= "000000";
					when "10010111010010100" => rgb <= "000000";
					when "10010111010010101" => rgb <= "000000";
					when "10010111010010110" => rgb <= "000000";
					when "10010111010010111" => rgb <= "000000";
					when "10010111010011000" => rgb <= "000000";
					when "10010111010011001" => rgb <= "000000";
					when "10010111010011010" => rgb <= "000000";
					when "10010111010011011" => rgb <= "000000";
					when "10010111010011100" => rgb <= "000000";
					when "10010111010011101" => rgb <= "000000";
					when "10010111010011110" => rgb <= "000000";
					when "10010111010011111" => rgb <= "000000";
					when "10010111010100000" => rgb <= "000000";
					when "10010111010100001" => rgb <= "000000";
					when "10010111010100010" => rgb <= "000000";
					when "10010111010100011" => rgb <= "000000";
					when "10010111010100100" => rgb <= "000000";
					when "10010111010100101" => rgb <= "000000";
					when "10010111010100110" => rgb <= "000000";
					when "10010111010100111" => rgb <= "000000";
					when "10010111010101000" => rgb <= "000000";
					when "10010111010101001" => rgb <= "000000";
					when "10010111010101010" => rgb <= "000000";
					when "10010111010101011" => rgb <= "000000";
					when "10010111010101100" => rgb <= "000000";
					when "10010111010101101" => rgb <= "000000";
					when "10010111010101110" => rgb <= "000000";
					when "10010111010101111" => rgb <= "000000";
					when "10010111010110000" => rgb <= "000000";
					when "10010111010110001" => rgb <= "000000";
					when "10010111010110010" => rgb <= "000000";
					when "10010111010110011" => rgb <= "000000";
					when "10010111010110100" => rgb <= "000000";
					when "10010111010110101" => rgb <= "000000";
					when "10010111010110110" => rgb <= "000000";
					when "10010111010110111" => rgb <= "000000";
					when "10010111010111000" => rgb <= "000000";
					when "10010111010111001" => rgb <= "000000";
					when "10010111010111010" => rgb <= "000000";
					when "10010111010111011" => rgb <= "000000";
					when "10010111010111100" => rgb <= "000000";
					when "10010111010111101" => rgb <= "000000";
					when "10010111010111110" => rgb <= "000000";
					when "10010111010111111" => rgb <= "000000";
					when "10010111011000000" => rgb <= "000000";
					when "10010111011000001" => rgb <= "000000";
					when "10010111011000010" => rgb <= "000000";
					when "10010111011000011" => rgb <= "000000";
					when "10010111011000100" => rgb <= "000000";
					when "10010111011000101" => rgb <= "000000";
					when "10010111011000110" => rgb <= "000000";
					when "10010111011000111" => rgb <= "000000";
					when "10010111011001000" => rgb <= "000000";
					when "10010111011001001" => rgb <= "000000";
					when "10010111011001010" => rgb <= "000000";
					when "10010111011001011" => rgb <= "000000";
					when "10010111011001100" => rgb <= "000000";
					when "10010111011001101" => rgb <= "000000";
					when "10010111011001110" => rgb <= "000000";
					when "10010111011001111" => rgb <= "000000";
					when "10010111011010000" => rgb <= "000000";
					when "10010111011010001" => rgb <= "000000";
					when "10010111011010010" => rgb <= "000000";
					when "10010111011010011" => rgb <= "000000";
					when "10010111011010100" => rgb <= "000000";
					when "10010111011010101" => rgb <= "000000";
					when "10010111011010110" => rgb <= "000000";
					when "10010111011010111" => rgb <= "000000";
					when "10010111011011000" => rgb <= "000000";
					when "10010111011011001" => rgb <= "000000";
					when "10010111011011010" => rgb <= "000000";
					when "10010111011011011" => rgb <= "000000";
					when "10010111011011100" => rgb <= "000000";
					when "10010111011011101" => rgb <= "000000";
					when "10010111011011110" => rgb <= "000000";
					when "10010111011011111" => rgb <= "000000";
					when "10010111011100000" => rgb <= "000000";
					when "10010111011100001" => rgb <= "000000";
					when "10010111011100010" => rgb <= "000000";
					when "10010111011100011" => rgb <= "000000";
					when "10010111011100100" => rgb <= "000000";
					when "10010111011100101" => rgb <= "000000";
					when "10010111011100110" => rgb <= "000000";
					when "10010111011100111" => rgb <= "000000";
					when "10010111011101000" => rgb <= "000000";
					when "10010111011101001" => rgb <= "000000";
					when "10010111011101010" => rgb <= "000000";
					when "10010111011101011" => rgb <= "000000";
					when "10010111011101100" => rgb <= "000000";
					when "10010111011101101" => rgb <= "000000";
					when "10010111011101110" => rgb <= "000000";
					when "10010111011101111" => rgb <= "000000";
					when "10010111011110000" => rgb <= "000000";
					when "10010111011110001" => rgb <= "000000";
					when "10010111011110010" => rgb <= "000000";
					when "10010111011110011" => rgb <= "000000";
					when "10010111011110100" => rgb <= "000000";
					when "10010111011110101" => rgb <= "000000";
					when "10010111011110110" => rgb <= "000000";
					when "10010111011110111" => rgb <= "000000";
					when "10010111011111000" => rgb <= "000000";
					when "10010111011111001" => rgb <= "000000";
					when "10010111011111010" => rgb <= "000000";
					when "10010111011111011" => rgb <= "000000";
					when "10010111011111100" => rgb <= "000000";
					when "10010111011111101" => rgb <= "000000";
					when "10010111011111110" => rgb <= "000000";
					when "10010111011111111" => rgb <= "000000";
					when "10010111100000000" => rgb <= "000000";
					when "10010111100000001" => rgb <= "000000";
					when "10010111100000010" => rgb <= "000000";
					when "10010111100000011" => rgb <= "000000";
					when "10010111100000100" => rgb <= "000000";
					when "10010111100000101" => rgb <= "000000";
					when "10010111100000110" => rgb <= "000000";
					when "10010111100000111" => rgb <= "000000";
					when "10010111100001000" => rgb <= "000000";
					when "10010111100001001" => rgb <= "000000";
					when "10010111100001010" => rgb <= "000000";
					when "10010111100001011" => rgb <= "000000";
					when "10010111100001100" => rgb <= "000000";
					when "10010111100001101" => rgb <= "000000";
					when "10010111100001110" => rgb <= "000000";
					when "10010111100001111" => rgb <= "000000";
					when "10010111100010000" => rgb <= "000000";
					when "10010111100010001" => rgb <= "000000";
					when "10010111100010010" => rgb <= "000000";
					when "10010111100010011" => rgb <= "000000";
					when "10010111100010100" => rgb <= "000000";
					when "10010111100010101" => rgb <= "000000";
					when "10010111100010110" => rgb <= "000000";
					when "10010111100010111" => rgb <= "000000";
					when "10010111100011000" => rgb <= "000000";
					when "10010111100011001" => rgb <= "000000";
					when "10010111100011010" => rgb <= "000000";
					when "10010111100011011" => rgb <= "000000";
					when "10010111100011100" => rgb <= "000000";
					when "10010111100011101" => rgb <= "000000";
					when "10010111100011110" => rgb <= "000000";
					when "10010111100011111" => rgb <= "000000";
					when "10010111100100000" => rgb <= "000000";
					when "10010111100100001" => rgb <= "000000";
					when "10010111100100010" => rgb <= "000000";
					when "10010111100100011" => rgb <= "000000";
					when "10010111100100100" => rgb <= "000000";
					when "10010111100100101" => rgb <= "000000";
					when "10010111100100110" => rgb <= "000000";
					when "10010111100100111" => rgb <= "000000";
					when "10010111100101000" => rgb <= "000000";
					when "10010111100101001" => rgb <= "000000";
					when "10010111100101010" => rgb <= "000000";
					when "10010111100101011" => rgb <= "000000";
					when "10010111100101100" => rgb <= "000000";
					when "10010111100101101" => rgb <= "000000";
					when "10010111100101110" => rgb <= "000000";
					when "10010111100101111" => rgb <= "000000";
					when "10010111100110000" => rgb <= "000000";
					when "10010111100110001" => rgb <= "000000";
					when "10010111100110010" => rgb <= "000000";
					when "10010111100110011" => rgb <= "000000";
					when "10010111100110100" => rgb <= "000000";
					when "10010111100110101" => rgb <= "000000";
					when "10010111100110110" => rgb <= "000000";
					when "10010111100110111" => rgb <= "000000";
					when "10010111100111000" => rgb <= "000000";
					when "10010111100111001" => rgb <= "000000";
					when "10010111100111010" => rgb <= "000000";
					when "10010111100111011" => rgb <= "000000";
					when "10010111100111100" => rgb <= "000000";
					when "10010111100111101" => rgb <= "000000";
					when "10010111100111110" => rgb <= "000000";
					when "10010111100111111" => rgb <= "000000";
					when "10011000000000000" => rgb <= "000000";
					when "10011000000000001" => rgb <= "000000";
					when "10011000000000010" => rgb <= "000000";
					when "10011000000000011" => rgb <= "000000";
					when "10011000000000100" => rgb <= "000000";
					when "10011000000000101" => rgb <= "000000";
					when "10011000000000110" => rgb <= "000000";
					when "10011000000000111" => rgb <= "000000";
					when "10011000000001000" => rgb <= "000000";
					when "10011000000001001" => rgb <= "000000";
					when "10011000000001010" => rgb <= "000000";
					when "10011000000001011" => rgb <= "000000";
					when "10011000000001100" => rgb <= "000000";
					when "10011000000001101" => rgb <= "000000";
					when "10011000000001110" => rgb <= "000000";
					when "10011000000001111" => rgb <= "000000";
					when "10011000000010000" => rgb <= "000000";
					when "10011000000010001" => rgb <= "000000";
					when "10011000000010010" => rgb <= "000000";
					when "10011000000010011" => rgb <= "000000";
					when "10011000000010100" => rgb <= "000000";
					when "10011000000010101" => rgb <= "000000";
					when "10011000000010110" => rgb <= "000000";
					when "10011000000010111" => rgb <= "000000";
					when "10011000000011000" => rgb <= "000000";
					when "10011000000011001" => rgb <= "000000";
					when "10011000000011010" => rgb <= "000000";
					when "10011000000011011" => rgb <= "000000";
					when "10011000000011100" => rgb <= "000000";
					when "10011000000011101" => rgb <= "000000";
					when "10011000000011110" => rgb <= "000000";
					when "10011000000011111" => rgb <= "000000";
					when "10011000000100000" => rgb <= "000000";
					when "10011000000100001" => rgb <= "000000";
					when "10011000000100010" => rgb <= "000000";
					when "10011000000100011" => rgb <= "000000";
					when "10011000000100100" => rgb <= "000000";
					when "10011000000100101" => rgb <= "000000";
					when "10011000000100110" => rgb <= "000000";
					when "10011000000100111" => rgb <= "000000";
					when "10011000000101000" => rgb <= "000000";
					when "10011000000101001" => rgb <= "000000";
					when "10011000000101010" => rgb <= "000000";
					when "10011000000101011" => rgb <= "000000";
					when "10011000000101100" => rgb <= "000000";
					when "10011000000101101" => rgb <= "000000";
					when "10011000000101110" => rgb <= "000000";
					when "10011000000101111" => rgb <= "000000";
					when "10011000000110000" => rgb <= "000000";
					when "10011000000110001" => rgb <= "000000";
					when "10011000000110010" => rgb <= "000000";
					when "10011000000110011" => rgb <= "000000";
					when "10011000000110100" => rgb <= "000000";
					when "10011000000110101" => rgb <= "000000";
					when "10011000000110110" => rgb <= "000000";
					when "10011000000110111" => rgb <= "000000";
					when "10011000000111000" => rgb <= "000000";
					when "10011000000111001" => rgb <= "000000";
					when "10011000000111010" => rgb <= "000000";
					when "10011000000111011" => rgb <= "000000";
					when "10011000000111100" => rgb <= "000000";
					when "10011000000111101" => rgb <= "000000";
					when "10011000000111110" => rgb <= "000000";
					when "10011000000111111" => rgb <= "000000";
					when "10011000001000000" => rgb <= "000000";
					when "10011000001000001" => rgb <= "000000";
					when "10011000001000010" => rgb <= "000000";
					when "10011000001000011" => rgb <= "000000";
					when "10011000001000100" => rgb <= "000000";
					when "10011000001000101" => rgb <= "000000";
					when "10011000001000110" => rgb <= "000000";
					when "10011000001000111" => rgb <= "000000";
					when "10011000001001000" => rgb <= "000000";
					when "10011000001001001" => rgb <= "000000";
					when "10011000001001010" => rgb <= "000000";
					when "10011000001001011" => rgb <= "000000";
					when "10011000001001100" => rgb <= "000000";
					when "10011000001001101" => rgb <= "000000";
					when "10011000001001110" => rgb <= "000000";
					when "10011000001001111" => rgb <= "000000";
					when "10011000001010000" => rgb <= "000000";
					when "10011000001010001" => rgb <= "000000";
					when "10011000001010010" => rgb <= "000000";
					when "10011000001010011" => rgb <= "000000";
					when "10011000001010100" => rgb <= "000000";
					when "10011000001010101" => rgb <= "000000";
					when "10011000001010110" => rgb <= "000000";
					when "10011000001010111" => rgb <= "000000";
					when "10011000001011000" => rgb <= "000000";
					when "10011000001011001" => rgb <= "000000";
					when "10011000001011010" => rgb <= "000000";
					when "10011000001011011" => rgb <= "000000";
					when "10011000001011100" => rgb <= "000000";
					when "10011000001011101" => rgb <= "000000";
					when "10011000001011110" => rgb <= "000000";
					when "10011000001011111" => rgb <= "000000";
					when "10011000001100000" => rgb <= "000000";
					when "10011000001100001" => rgb <= "000000";
					when "10011000001100010" => rgb <= "000000";
					when "10011000001100011" => rgb <= "000000";
					when "10011000001100100" => rgb <= "000000";
					when "10011000001100101" => rgb <= "000000";
					when "10011000001100110" => rgb <= "000000";
					when "10011000001100111" => rgb <= "000000";
					when "10011000001101000" => rgb <= "000000";
					when "10011000001101001" => rgb <= "000000";
					when "10011000001101010" => rgb <= "000000";
					when "10011000001101011" => rgb <= "000000";
					when "10011000001101100" => rgb <= "000000";
					when "10011000001101101" => rgb <= "000000";
					when "10011000001101110" => rgb <= "000000";
					when "10011000001101111" => rgb <= "000000";
					when "10011000001110000" => rgb <= "000000";
					when "10011000001110001" => rgb <= "000000";
					when "10011000001110010" => rgb <= "000000";
					when "10011000001110011" => rgb <= "000000";
					when "10011000001110100" => rgb <= "000000";
					when "10011000001110101" => rgb <= "000000";
					when "10011000001110110" => rgb <= "000000";
					when "10011000001110111" => rgb <= "000000";
					when "10011000001111000" => rgb <= "000000";
					when "10011000001111001" => rgb <= "000000";
					when "10011000001111010" => rgb <= "000000";
					when "10011000001111011" => rgb <= "000000";
					when "10011000001111100" => rgb <= "000000";
					when "10011000001111101" => rgb <= "000000";
					when "10011000001111110" => rgb <= "000000";
					when "10011000001111111" => rgb <= "000000";
					when "10011000010000000" => rgb <= "000000";
					when "10011000010000001" => rgb <= "000000";
					when "10011000010000010" => rgb <= "000000";
					when "10011000010000011" => rgb <= "000000";
					when "10011000010000100" => rgb <= "000000";
					when "10011000010000101" => rgb <= "000000";
					when "10011000010000110" => rgb <= "000000";
					when "10011000010000111" => rgb <= "000000";
					when "10011000010001000" => rgb <= "000000";
					when "10011000010001001" => rgb <= "000000";
					when "10011000010001010" => rgb <= "000000";
					when "10011000010001011" => rgb <= "000000";
					when "10011000010001100" => rgb <= "000000";
					when "10011000010001101" => rgb <= "000000";
					when "10011000010001110" => rgb <= "000000";
					when "10011000010001111" => rgb <= "000000";
					when "10011000010010000" => rgb <= "000000";
					when "10011000010010001" => rgb <= "000000";
					when "10011000010010010" => rgb <= "000000";
					when "10011000010010011" => rgb <= "000000";
					when "10011000010010100" => rgb <= "000000";
					when "10011000010010101" => rgb <= "000000";
					when "10011000010010110" => rgb <= "000000";
					when "10011000010010111" => rgb <= "000000";
					when "10011000010011000" => rgb <= "000000";
					when "10011000010011001" => rgb <= "000000";
					when "10011000010011010" => rgb <= "000000";
					when "10011000010011011" => rgb <= "000000";
					when "10011000010011100" => rgb <= "000000";
					when "10011000010011101" => rgb <= "000000";
					when "10011000010011110" => rgb <= "000000";
					when "10011000010011111" => rgb <= "000000";
					when "10011000010100000" => rgb <= "000000";
					when "10011000010100001" => rgb <= "000000";
					when "10011000010100010" => rgb <= "000000";
					when "10011000010100011" => rgb <= "000000";
					when "10011000010100100" => rgb <= "000000";
					when "10011000010100101" => rgb <= "000000";
					when "10011000010100110" => rgb <= "000000";
					when "10011000010100111" => rgb <= "000000";
					when "10011000010101000" => rgb <= "000000";
					when "10011000010101001" => rgb <= "000000";
					when "10011000010101010" => rgb <= "000000";
					when "10011000010101011" => rgb <= "000000";
					when "10011000010101100" => rgb <= "000000";
					when "10011000010101101" => rgb <= "000000";
					when "10011000010101110" => rgb <= "000000";
					when "10011000010101111" => rgb <= "000000";
					when "10011000010110000" => rgb <= "000000";
					when "10011000010110001" => rgb <= "000000";
					when "10011000010110010" => rgb <= "000000";
					when "10011000010110011" => rgb <= "000000";
					when "10011000010110100" => rgb <= "000000";
					when "10011000010110101" => rgb <= "000000";
					when "10011000010110110" => rgb <= "000000";
					when "10011000010110111" => rgb <= "000000";
					when "10011000010111000" => rgb <= "000000";
					when "10011000010111001" => rgb <= "000000";
					when "10011000010111010" => rgb <= "000000";
					when "10011000010111011" => rgb <= "000000";
					when "10011000010111100" => rgb <= "000000";
					when "10011000010111101" => rgb <= "000000";
					when "10011000010111110" => rgb <= "000000";
					when "10011000010111111" => rgb <= "000000";
					when "10011000011000000" => rgb <= "000000";
					when "10011000011000001" => rgb <= "000000";
					when "10011000011000010" => rgb <= "000000";
					when "10011000011000011" => rgb <= "000000";
					when "10011000011000100" => rgb <= "000000";
					when "10011000011000101" => rgb <= "000000";
					when "10011000011000110" => rgb <= "000000";
					when "10011000011000111" => rgb <= "000000";
					when "10011000011001000" => rgb <= "000000";
					when "10011000011001001" => rgb <= "000000";
					when "10011000011001010" => rgb <= "000000";
					when "10011000011001011" => rgb <= "000000";
					when "10011000011001100" => rgb <= "000000";
					when "10011000011001101" => rgb <= "000000";
					when "10011000011001110" => rgb <= "000000";
					when "10011000011001111" => rgb <= "000000";
					when "10011000011010000" => rgb <= "000000";
					when "10011000011010001" => rgb <= "000000";
					when "10011000011010010" => rgb <= "000000";
					when "10011000011010011" => rgb <= "000000";
					when "10011000011010100" => rgb <= "000000";
					when "10011000011010101" => rgb <= "000000";
					when "10011000011010110" => rgb <= "000000";
					when "10011000011010111" => rgb <= "000000";
					when "10011000011011000" => rgb <= "000000";
					when "10011000011011001" => rgb <= "000000";
					when "10011000011011010" => rgb <= "000000";
					when "10011000011011011" => rgb <= "000000";
					when "10011000011011100" => rgb <= "000000";
					when "10011000011011101" => rgb <= "000000";
					when "10011000011011110" => rgb <= "000000";
					when "10011000011011111" => rgb <= "000000";
					when "10011000011100000" => rgb <= "000000";
					when "10011000011100001" => rgb <= "000000";
					when "10011000011100010" => rgb <= "000000";
					when "10011000011100011" => rgb <= "000000";
					when "10011000011100100" => rgb <= "000000";
					when "10011000011100101" => rgb <= "000000";
					when "10011000011100110" => rgb <= "000000";
					when "10011000011100111" => rgb <= "000000";
					when "10011000011101000" => rgb <= "000000";
					when "10011000011101001" => rgb <= "000000";
					when "10011000011101010" => rgb <= "000000";
					when "10011000011101011" => rgb <= "000000";
					when "10011000011101100" => rgb <= "000000";
					when "10011000011101101" => rgb <= "000000";
					when "10011000011101110" => rgb <= "000000";
					when "10011000011101111" => rgb <= "000000";
					when "10011000011110000" => rgb <= "000000";
					when "10011000011110001" => rgb <= "000000";
					when "10011000011110010" => rgb <= "000000";
					when "10011000011110011" => rgb <= "000000";
					when "10011000011110100" => rgb <= "000000";
					when "10011000011110101" => rgb <= "000000";
					when "10011000011110110" => rgb <= "000000";
					when "10011000011110111" => rgb <= "000000";
					when "10011000011111000" => rgb <= "000000";
					when "10011000011111001" => rgb <= "000000";
					when "10011000011111010" => rgb <= "000000";
					when "10011000011111011" => rgb <= "000000";
					when "10011000011111100" => rgb <= "000000";
					when "10011000011111101" => rgb <= "000000";
					when "10011000011111110" => rgb <= "000000";
					when "10011000011111111" => rgb <= "000000";
					when "10011000100000000" => rgb <= "000000";
					when "10011000100000001" => rgb <= "000000";
					when "10011000100000010" => rgb <= "000000";
					when "10011000100000011" => rgb <= "000000";
					when "10011000100000100" => rgb <= "000000";
					when "10011000100000101" => rgb <= "000000";
					when "10011000100000110" => rgb <= "000000";
					when "10011000100000111" => rgb <= "000000";
					when "10011000100001000" => rgb <= "000000";
					when "10011000100001001" => rgb <= "000000";
					when "10011000100001010" => rgb <= "000000";
					when "10011000100001011" => rgb <= "000000";
					when "10011000100001100" => rgb <= "000000";
					when "10011000100001101" => rgb <= "000000";
					when "10011000100001110" => rgb <= "000000";
					when "10011000100001111" => rgb <= "000000";
					when "10011000100010000" => rgb <= "000000";
					when "10011000100010001" => rgb <= "000000";
					when "10011000100010010" => rgb <= "000000";
					when "10011000100010011" => rgb <= "000000";
					when "10011000100010100" => rgb <= "000000";
					when "10011000100010101" => rgb <= "000000";
					when "10011000100010110" => rgb <= "000000";
					when "10011000100010111" => rgb <= "000000";
					when "10011000100011000" => rgb <= "000000";
					when "10011000100011001" => rgb <= "000000";
					when "10011000100011010" => rgb <= "000000";
					when "10011000100011011" => rgb <= "000000";
					when "10011000100011100" => rgb <= "000000";
					when "10011000100011101" => rgb <= "000000";
					when "10011000100011110" => rgb <= "000000";
					when "10011000100011111" => rgb <= "000000";
					when "10011000100100000" => rgb <= "000000";
					when "10011000100100001" => rgb <= "000000";
					when "10011000100100010" => rgb <= "000000";
					when "10011000100100011" => rgb <= "000000";
					when "10011000100100100" => rgb <= "000000";
					when "10011000100100101" => rgb <= "000000";
					when "10011000100100110" => rgb <= "000000";
					when "10011000100100111" => rgb <= "000000";
					when "10011000100101000" => rgb <= "000000";
					when "10011000100101001" => rgb <= "000000";
					when "10011000100101010" => rgb <= "000000";
					when "10011000100101011" => rgb <= "000000";
					when "10011000100101100" => rgb <= "000000";
					when "10011000100101101" => rgb <= "000000";
					when "10011000100101110" => rgb <= "000000";
					when "10011000100101111" => rgb <= "000000";
					when "10011000100110000" => rgb <= "000000";
					when "10011000100110001" => rgb <= "000000";
					when "10011000100110010" => rgb <= "000000";
					when "10011000100110011" => rgb <= "000000";
					when "10011000100110100" => rgb <= "000000";
					when "10011000100110101" => rgb <= "000000";
					when "10011000100110110" => rgb <= "000000";
					when "10011000100110111" => rgb <= "000000";
					when "10011000100111000" => rgb <= "000000";
					when "10011000100111001" => rgb <= "000000";
					when "10011000100111010" => rgb <= "000000";
					when "10011000100111011" => rgb <= "000000";
					when "10011000100111100" => rgb <= "000000";
					when "10011000100111101" => rgb <= "000000";
					when "10011000100111110" => rgb <= "000000";
					when "10011000100111111" => rgb <= "000000";
					when "10011001000000000" => rgb <= "000000";
					when "10011001000000001" => rgb <= "000000";
					when "10011001000000010" => rgb <= "000000";
					when "10011001000000011" => rgb <= "000000";
					when "10011001000000100" => rgb <= "000000";
					when "10011001000000101" => rgb <= "000000";
					when "10011001000000110" => rgb <= "000000";
					when "10011001000000111" => rgb <= "000000";
					when "10011001000001000" => rgb <= "000000";
					when "10011001000001001" => rgb <= "000000";
					when "10011001000001010" => rgb <= "000000";
					when "10011001000001011" => rgb <= "000000";
					when "10011001000001100" => rgb <= "000000";
					when "10011001000001101" => rgb <= "000000";
					when "10011001000001110" => rgb <= "000000";
					when "10011001000001111" => rgb <= "000000";
					when "10011001000010000" => rgb <= "000000";
					when "10011001000010001" => rgb <= "000000";
					when "10011001000010010" => rgb <= "000000";
					when "10011001000010011" => rgb <= "000000";
					when "10011001000010100" => rgb <= "000000";
					when "10011001000010101" => rgb <= "000000";
					when "10011001000010110" => rgb <= "000000";
					when "10011001000010111" => rgb <= "000000";
					when "10011001000011000" => rgb <= "000000";
					when "10011001000011001" => rgb <= "000000";
					when "10011001000011010" => rgb <= "000000";
					when "10011001000011011" => rgb <= "000000";
					when "10011001000011100" => rgb <= "000000";
					when "10011001000011101" => rgb <= "000000";
					when "10011001000011110" => rgb <= "000000";
					when "10011001000011111" => rgb <= "000000";
					when "10011001000100000" => rgb <= "000000";
					when "10011001000100001" => rgb <= "000000";
					when "10011001000100010" => rgb <= "000000";
					when "10011001000100011" => rgb <= "000000";
					when "10011001000100100" => rgb <= "000000";
					when "10011001000100101" => rgb <= "000000";
					when "10011001000100110" => rgb <= "000000";
					when "10011001000100111" => rgb <= "000000";
					when "10011001000101000" => rgb <= "000000";
					when "10011001000101001" => rgb <= "000000";
					when "10011001000101010" => rgb <= "000000";
					when "10011001000101011" => rgb <= "000000";
					when "10011001000101100" => rgb <= "000000";
					when "10011001000101101" => rgb <= "000000";
					when "10011001000101110" => rgb <= "000000";
					when "10011001000101111" => rgb <= "000000";
					when "10011001000110000" => rgb <= "000000";
					when "10011001000110001" => rgb <= "000000";
					when "10011001000110010" => rgb <= "000000";
					when "10011001000110011" => rgb <= "000000";
					when "10011001000110100" => rgb <= "000000";
					when "10011001000110101" => rgb <= "000000";
					when "10011001000110110" => rgb <= "000000";
					when "10011001000110111" => rgb <= "000000";
					when "10011001000111000" => rgb <= "000000";
					when "10011001000111001" => rgb <= "000000";
					when "10011001000111010" => rgb <= "000000";
					when "10011001000111011" => rgb <= "000000";
					when "10011001000111100" => rgb <= "000000";
					when "10011001000111101" => rgb <= "000000";
					when "10011001000111110" => rgb <= "000000";
					when "10011001000111111" => rgb <= "000000";
					when "10011001001000000" => rgb <= "000000";
					when "10011001001000001" => rgb <= "000000";
					when "10011001001000010" => rgb <= "000000";
					when "10011001001000011" => rgb <= "000000";
					when "10011001001000100" => rgb <= "000000";
					when "10011001001000101" => rgb <= "000000";
					when "10011001001000110" => rgb <= "000000";
					when "10011001001000111" => rgb <= "000000";
					when "10011001001001000" => rgb <= "000000";
					when "10011001001001001" => rgb <= "000000";
					when "10011001001001010" => rgb <= "000000";
					when "10011001001001011" => rgb <= "000000";
					when "10011001001001100" => rgb <= "000000";
					when "10011001001001101" => rgb <= "000000";
					when "10011001001001110" => rgb <= "000000";
					when "10011001001001111" => rgb <= "000000";
					when "10011001001010000" => rgb <= "000000";
					when "10011001001010001" => rgb <= "000000";
					when "10011001001010010" => rgb <= "000000";
					when "10011001001010011" => rgb <= "000000";
					when "10011001001010100" => rgb <= "000000";
					when "10011001001010101" => rgb <= "000000";
					when "10011001001010110" => rgb <= "000000";
					when "10011001001010111" => rgb <= "000000";
					when "10011001001011000" => rgb <= "000000";
					when "10011001001011001" => rgb <= "000000";
					when "10011001001011010" => rgb <= "000000";
					when "10011001001011011" => rgb <= "000000";
					when "10011001001011100" => rgb <= "000000";
					when "10011001001011101" => rgb <= "000000";
					when "10011001001011110" => rgb <= "000000";
					when "10011001001011111" => rgb <= "000000";
					when "10011001001100000" => rgb <= "000000";
					when "10011001001100001" => rgb <= "000000";
					when "10011001001100010" => rgb <= "000000";
					when "10011001001100011" => rgb <= "000000";
					when "10011001001100100" => rgb <= "000000";
					when "10011001001100101" => rgb <= "000000";
					when "10011001001100110" => rgb <= "000000";
					when "10011001001100111" => rgb <= "000000";
					when "10011001001101000" => rgb <= "000000";
					when "10011001001101001" => rgb <= "000000";
					when "10011001001101010" => rgb <= "000000";
					when "10011001001101011" => rgb <= "000000";
					when "10011001001101100" => rgb <= "000000";
					when "10011001001101101" => rgb <= "000000";
					when "10011001001101110" => rgb <= "000000";
					when "10011001001101111" => rgb <= "000000";
					when "10011001001110000" => rgb <= "000000";
					when "10011001001110001" => rgb <= "000000";
					when "10011001001110010" => rgb <= "000000";
					when "10011001001110011" => rgb <= "000000";
					when "10011001001110100" => rgb <= "000000";
					when "10011001001110101" => rgb <= "000000";
					when "10011001001110110" => rgb <= "000000";
					when "10011001001110111" => rgb <= "000000";
					when "10011001001111000" => rgb <= "000000";
					when "10011001001111001" => rgb <= "000000";
					when "10011001001111010" => rgb <= "000000";
					when "10011001001111011" => rgb <= "000000";
					when "10011001001111100" => rgb <= "000000";
					when "10011001001111101" => rgb <= "000000";
					when "10011001001111110" => rgb <= "000000";
					when "10011001001111111" => rgb <= "000000";
					when "10011001010000000" => rgb <= "000000";
					when "10011001010000001" => rgb <= "000000";
					when "10011001010000010" => rgb <= "000000";
					when "10011001010000011" => rgb <= "000000";
					when "10011001010000100" => rgb <= "000000";
					when "10011001010000101" => rgb <= "000000";
					when "10011001010000110" => rgb <= "000000";
					when "10011001010000111" => rgb <= "000000";
					when "10011001010001000" => rgb <= "000000";
					when "10011001010001001" => rgb <= "000000";
					when "10011001010001010" => rgb <= "000000";
					when "10011001010001011" => rgb <= "000000";
					when "10011001010001100" => rgb <= "000000";
					when "10011001010001101" => rgb <= "000000";
					when "10011001010001110" => rgb <= "000000";
					when "10011001010001111" => rgb <= "000000";
					when "10011001010010000" => rgb <= "000000";
					when "10011001010010001" => rgb <= "000000";
					when "10011001010010010" => rgb <= "000000";
					when "10011001010010011" => rgb <= "000000";
					when "10011001010010100" => rgb <= "000000";
					when "10011001010010101" => rgb <= "000000";
					when "10011001010010110" => rgb <= "000000";
					when "10011001010010111" => rgb <= "000000";
					when "10011001010011000" => rgb <= "000000";
					when "10011001010011001" => rgb <= "000000";
					when "10011001010011010" => rgb <= "000000";
					when "10011001010011011" => rgb <= "000000";
					when "10011001010011100" => rgb <= "000000";
					when "10011001010011101" => rgb <= "000000";
					when "10011001010011110" => rgb <= "000000";
					when "10011001010011111" => rgb <= "000000";
					when "10011001010100000" => rgb <= "000000";
					when "10011001010100001" => rgb <= "000000";
					when "10011001010100010" => rgb <= "000000";
					when "10011001010100011" => rgb <= "000000";
					when "10011001010100100" => rgb <= "000000";
					when "10011001010100101" => rgb <= "000000";
					when "10011001010100110" => rgb <= "000000";
					when "10011001010100111" => rgb <= "000000";
					when "10011001010101000" => rgb <= "000000";
					when "10011001010101001" => rgb <= "000000";
					when "10011001010101010" => rgb <= "000000";
					when "10011001010101011" => rgb <= "000000";
					when "10011001010101100" => rgb <= "000000";
					when "10011001010101101" => rgb <= "000000";
					when "10011001010101110" => rgb <= "000000";
					when "10011001010101111" => rgb <= "000000";
					when "10011001010110000" => rgb <= "000000";
					when "10011001010110001" => rgb <= "000000";
					when "10011001010110010" => rgb <= "000000";
					when "10011001010110011" => rgb <= "000000";
					when "10011001010110100" => rgb <= "000000";
					when "10011001010110101" => rgb <= "000000";
					when "10011001010110110" => rgb <= "000000";
					when "10011001010110111" => rgb <= "000000";
					when "10011001010111000" => rgb <= "000000";
					when "10011001010111001" => rgb <= "000000";
					when "10011001010111010" => rgb <= "000000";
					when "10011001010111011" => rgb <= "000000";
					when "10011001010111100" => rgb <= "000000";
					when "10011001010111101" => rgb <= "000000";
					when "10011001010111110" => rgb <= "000000";
					when "10011001010111111" => rgb <= "000000";
					when "10011001011000000" => rgb <= "000000";
					when "10011001011000001" => rgb <= "000000";
					when "10011001011000010" => rgb <= "000000";
					when "10011001011000011" => rgb <= "000000";
					when "10011001011000100" => rgb <= "000000";
					when "10011001011000101" => rgb <= "000000";
					when "10011001011000110" => rgb <= "000000";
					when "10011001011000111" => rgb <= "000000";
					when "10011001011001000" => rgb <= "000000";
					when "10011001011001001" => rgb <= "000000";
					when "10011001011001010" => rgb <= "000000";
					when "10011001011001011" => rgb <= "000000";
					when "10011001011001100" => rgb <= "000000";
					when "10011001011001101" => rgb <= "000000";
					when "10011001011001110" => rgb <= "000000";
					when "10011001011001111" => rgb <= "000000";
					when "10011001011010000" => rgb <= "000000";
					when "10011001011010001" => rgb <= "000000";
					when "10011001011010010" => rgb <= "000000";
					when "10011001011010011" => rgb <= "000000";
					when "10011001011010100" => rgb <= "000000";
					when "10011001011010101" => rgb <= "000000";
					when "10011001011010110" => rgb <= "000000";
					when "10011001011010111" => rgb <= "000000";
					when "10011001011011000" => rgb <= "000000";
					when "10011001011011001" => rgb <= "000000";
					when "10011001011011010" => rgb <= "000000";
					when "10011001011011011" => rgb <= "000000";
					when "10011001011011100" => rgb <= "000000";
					when "10011001011011101" => rgb <= "000000";
					when "10011001011011110" => rgb <= "000000";
					when "10011001011011111" => rgb <= "000000";
					when "10011001011100000" => rgb <= "000000";
					when "10011001011100001" => rgb <= "000000";
					when "10011001011100010" => rgb <= "000000";
					when "10011001011100011" => rgb <= "000000";
					when "10011001011100100" => rgb <= "000000";
					when "10011001011100101" => rgb <= "000000";
					when "10011001011100110" => rgb <= "000000";
					when "10011001011100111" => rgb <= "000000";
					when "10011001011101000" => rgb <= "000000";
					when "10011001011101001" => rgb <= "000000";
					when "10011001011101010" => rgb <= "000000";
					when "10011001011101011" => rgb <= "000000";
					when "10011001011101100" => rgb <= "000000";
					when "10011001011101101" => rgb <= "000000";
					when "10011001011101110" => rgb <= "000000";
					when "10011001011101111" => rgb <= "000000";
					when "10011001011110000" => rgb <= "000000";
					when "10011001011110001" => rgb <= "000000";
					when "10011001011110010" => rgb <= "000000";
					when "10011001011110011" => rgb <= "000000";
					when "10011001011110100" => rgb <= "000000";
					when "10011001011110101" => rgb <= "000000";
					when "10011001011110110" => rgb <= "000000";
					when "10011001011110111" => rgb <= "000000";
					when "10011001011111000" => rgb <= "000000";
					when "10011001011111001" => rgb <= "000000";
					when "10011001011111010" => rgb <= "000000";
					when "10011001011111011" => rgb <= "000000";
					when "10011001011111100" => rgb <= "000000";
					when "10011001011111101" => rgb <= "000000";
					when "10011001011111110" => rgb <= "000000";
					when "10011001011111111" => rgb <= "000000";
					when "10011001100000000" => rgb <= "000000";
					when "10011001100000001" => rgb <= "000000";
					when "10011001100000010" => rgb <= "000000";
					when "10011001100000011" => rgb <= "000000";
					when "10011001100000100" => rgb <= "000000";
					when "10011001100000101" => rgb <= "000000";
					when "10011001100000110" => rgb <= "000000";
					when "10011001100000111" => rgb <= "000000";
					when "10011001100001000" => rgb <= "000000";
					when "10011001100001001" => rgb <= "000000";
					when "10011001100001010" => rgb <= "000000";
					when "10011001100001011" => rgb <= "000000";
					when "10011001100001100" => rgb <= "000000";
					when "10011001100001101" => rgb <= "000000";
					when "10011001100001110" => rgb <= "000000";
					when "10011001100001111" => rgb <= "000000";
					when "10011001100010000" => rgb <= "000000";
					when "10011001100010001" => rgb <= "000000";
					when "10011001100010010" => rgb <= "000000";
					when "10011001100010011" => rgb <= "000000";
					when "10011001100010100" => rgb <= "000000";
					when "10011001100010101" => rgb <= "000000";
					when "10011001100010110" => rgb <= "000000";
					when "10011001100010111" => rgb <= "000000";
					when "10011001100011000" => rgb <= "000000";
					when "10011001100011001" => rgb <= "000000";
					when "10011001100011010" => rgb <= "000000";
					when "10011001100011011" => rgb <= "000000";
					when "10011001100011100" => rgb <= "000000";
					when "10011001100011101" => rgb <= "000000";
					when "10011001100011110" => rgb <= "000000";
					when "10011001100011111" => rgb <= "000000";
					when "10011001100100000" => rgb <= "000000";
					when "10011001100100001" => rgb <= "000000";
					when "10011001100100010" => rgb <= "000000";
					when "10011001100100011" => rgb <= "000000";
					when "10011001100100100" => rgb <= "000000";
					when "10011001100100101" => rgb <= "000000";
					when "10011001100100110" => rgb <= "000000";
					when "10011001100100111" => rgb <= "000000";
					when "10011001100101000" => rgb <= "000000";
					when "10011001100101001" => rgb <= "000000";
					when "10011001100101010" => rgb <= "000000";
					when "10011001100101011" => rgb <= "000000";
					when "10011001100101100" => rgb <= "000000";
					when "10011001100101101" => rgb <= "000000";
					when "10011001100101110" => rgb <= "000000";
					when "10011001100101111" => rgb <= "000000";
					when "10011001100110000" => rgb <= "000000";
					when "10011001100110001" => rgb <= "000000";
					when "10011001100110010" => rgb <= "000000";
					when "10011001100110011" => rgb <= "000000";
					when "10011001100110100" => rgb <= "000000";
					when "10011001100110101" => rgb <= "000000";
					when "10011001100110110" => rgb <= "000000";
					when "10011001100110111" => rgb <= "000000";
					when "10011001100111000" => rgb <= "000000";
					when "10011001100111001" => rgb <= "000000";
					when "10011001100111010" => rgb <= "000000";
					when "10011001100111011" => rgb <= "000000";
					when "10011001100111100" => rgb <= "000000";
					when "10011001100111101" => rgb <= "000000";
					when "10011001100111110" => rgb <= "000000";
					when "10011001100111111" => rgb <= "000000";
					when "10011010000000000" => rgb <= "000000";
					when "10011010000000001" => rgb <= "000000";
					when "10011010000000010" => rgb <= "000000";
					when "10011010000000011" => rgb <= "000000";
					when "10011010000000100" => rgb <= "000000";
					when "10011010000000101" => rgb <= "000000";
					when "10011010000000110" => rgb <= "000000";
					when "10011010000000111" => rgb <= "000000";
					when "10011010000001000" => rgb <= "000000";
					when "10011010000001001" => rgb <= "000000";
					when "10011010000001010" => rgb <= "000000";
					when "10011010000001011" => rgb <= "000000";
					when "10011010000001100" => rgb <= "000000";
					when "10011010000001101" => rgb <= "000000";
					when "10011010000001110" => rgb <= "000000";
					when "10011010000001111" => rgb <= "000000";
					when "10011010000010000" => rgb <= "000000";
					when "10011010000010001" => rgb <= "000000";
					when "10011010000010010" => rgb <= "000000";
					when "10011010000010011" => rgb <= "000000";
					when "10011010000010100" => rgb <= "000000";
					when "10011010000010101" => rgb <= "000000";
					when "10011010000010110" => rgb <= "000000";
					when "10011010000010111" => rgb <= "000000";
					when "10011010000011000" => rgb <= "000000";
					when "10011010000011001" => rgb <= "000000";
					when "10011010000011010" => rgb <= "000000";
					when "10011010000011011" => rgb <= "000000";
					when "10011010000011100" => rgb <= "000000";
					when "10011010000011101" => rgb <= "000000";
					when "10011010000011110" => rgb <= "000000";
					when "10011010000011111" => rgb <= "000000";
					when "10011010000100000" => rgb <= "000000";
					when "10011010000100001" => rgb <= "000000";
					when "10011010000100010" => rgb <= "000000";
					when "10011010000100011" => rgb <= "000000";
					when "10011010000100100" => rgb <= "000000";
					when "10011010000100101" => rgb <= "000000";
					when "10011010000100110" => rgb <= "000000";
					when "10011010000100111" => rgb <= "000000";
					when "10011010000101000" => rgb <= "000000";
					when "10011010000101001" => rgb <= "000000";
					when "10011010000101010" => rgb <= "000000";
					when "10011010000101011" => rgb <= "000000";
					when "10011010000101100" => rgb <= "000000";
					when "10011010000101101" => rgb <= "000000";
					when "10011010000101110" => rgb <= "000000";
					when "10011010000101111" => rgb <= "000000";
					when "10011010000110000" => rgb <= "000000";
					when "10011010000110001" => rgb <= "000000";
					when "10011010000110010" => rgb <= "000000";
					when "10011010000110011" => rgb <= "000000";
					when "10011010000110100" => rgb <= "000000";
					when "10011010000110101" => rgb <= "000000";
					when "10011010000110110" => rgb <= "000000";
					when "10011010000110111" => rgb <= "000000";
					when "10011010000111000" => rgb <= "000000";
					when "10011010000111001" => rgb <= "000000";
					when "10011010000111010" => rgb <= "000000";
					when "10011010000111011" => rgb <= "000000";
					when "10011010000111100" => rgb <= "000000";
					when "10011010000111101" => rgb <= "000000";
					when "10011010000111110" => rgb <= "000000";
					when "10011010000111111" => rgb <= "000000";
					when "10011010001000000" => rgb <= "000000";
					when "10011010001000001" => rgb <= "000000";
					when "10011010001000010" => rgb <= "000000";
					when "10011010001000011" => rgb <= "000000";
					when "10011010001000100" => rgb <= "000000";
					when "10011010001000101" => rgb <= "000000";
					when "10011010001000110" => rgb <= "000000";
					when "10011010001000111" => rgb <= "000000";
					when "10011010001001000" => rgb <= "000000";
					when "10011010001001001" => rgb <= "000000";
					when "10011010001001010" => rgb <= "000000";
					when "10011010001001011" => rgb <= "000000";
					when "10011010001001100" => rgb <= "000000";
					when "10011010001001101" => rgb <= "000000";
					when "10011010001001110" => rgb <= "000000";
					when "10011010001001111" => rgb <= "000000";
					when "10011010001010000" => rgb <= "000000";
					when "10011010001010001" => rgb <= "000000";
					when "10011010001010010" => rgb <= "000000";
					when "10011010001010011" => rgb <= "000000";
					when "10011010001010100" => rgb <= "000000";
					when "10011010001010101" => rgb <= "000000";
					when "10011010001010110" => rgb <= "000000";
					when "10011010001010111" => rgb <= "000000";
					when "10011010001011000" => rgb <= "000000";
					when "10011010001011001" => rgb <= "000000";
					when "10011010001011010" => rgb <= "000000";
					when "10011010001011011" => rgb <= "000000";
					when "10011010001011100" => rgb <= "000000";
					when "10011010001011101" => rgb <= "000000";
					when "10011010001011110" => rgb <= "000000";
					when "10011010001011111" => rgb <= "000000";
					when "10011010001100000" => rgb <= "000000";
					when "10011010001100001" => rgb <= "000000";
					when "10011010001100010" => rgb <= "000000";
					when "10011010001100011" => rgb <= "000000";
					when "10011010001100100" => rgb <= "000000";
					when "10011010001100101" => rgb <= "000000";
					when "10011010001100110" => rgb <= "000000";
					when "10011010001100111" => rgb <= "000000";
					when "10011010001101000" => rgb <= "000000";
					when "10011010001101001" => rgb <= "000000";
					when "10011010001101010" => rgb <= "000000";
					when "10011010001101011" => rgb <= "000000";
					when "10011010001101100" => rgb <= "000000";
					when "10011010001101101" => rgb <= "000000";
					when "10011010001101110" => rgb <= "000000";
					when "10011010001101111" => rgb <= "000000";
					when "10011010001110000" => rgb <= "000000";
					when "10011010001110001" => rgb <= "000000";
					when "10011010001110010" => rgb <= "000000";
					when "10011010001110011" => rgb <= "000000";
					when "10011010001110100" => rgb <= "000000";
					when "10011010001110101" => rgb <= "000000";
					when "10011010001110110" => rgb <= "000000";
					when "10011010001110111" => rgb <= "000000";
					when "10011010001111000" => rgb <= "000000";
					when "10011010001111001" => rgb <= "000000";
					when "10011010001111010" => rgb <= "000000";
					when "10011010001111011" => rgb <= "000000";
					when "10011010001111100" => rgb <= "000000";
					when "10011010001111101" => rgb <= "000000";
					when "10011010001111110" => rgb <= "000000";
					when "10011010001111111" => rgb <= "000000";
					when "10011010010000000" => rgb <= "000000";
					when "10011010010000001" => rgb <= "000000";
					when "10011010010000010" => rgb <= "000000";
					when "10011010010000011" => rgb <= "000000";
					when "10011010010000100" => rgb <= "000000";
					when "10011010010000101" => rgb <= "000000";
					when "10011010010000110" => rgb <= "000000";
					when "10011010010000111" => rgb <= "000000";
					when "10011010010001000" => rgb <= "000000";
					when "10011010010001001" => rgb <= "000000";
					when "10011010010001010" => rgb <= "000000";
					when "10011010010001011" => rgb <= "000000";
					when "10011010010001100" => rgb <= "000000";
					when "10011010010001101" => rgb <= "000000";
					when "10011010010001110" => rgb <= "000000";
					when "10011010010001111" => rgb <= "000000";
					when "10011010010010000" => rgb <= "000000";
					when "10011010010010001" => rgb <= "000000";
					when "10011010010010010" => rgb <= "000000";
					when "10011010010010011" => rgb <= "000000";
					when "10011010010010100" => rgb <= "000000";
					when "10011010010010101" => rgb <= "000000";
					when "10011010010010110" => rgb <= "000000";
					when "10011010010010111" => rgb <= "000000";
					when "10011010010011000" => rgb <= "000000";
					when "10011010010011001" => rgb <= "000000";
					when "10011010010011010" => rgb <= "000000";
					when "10011010010011011" => rgb <= "000000";
					when "10011010010011100" => rgb <= "000000";
					when "10011010010011101" => rgb <= "000000";
					when "10011010010011110" => rgb <= "000000";
					when "10011010010011111" => rgb <= "000000";
					when "10011010010100000" => rgb <= "000000";
					when "10011010010100001" => rgb <= "000000";
					when "10011010010100010" => rgb <= "000000";
					when "10011010010100011" => rgb <= "000000";
					when "10011010010100100" => rgb <= "000000";
					when "10011010010100101" => rgb <= "000000";
					when "10011010010100110" => rgb <= "000000";
					when "10011010010100111" => rgb <= "000000";
					when "10011010010101000" => rgb <= "000000";
					when "10011010010101001" => rgb <= "000000";
					when "10011010010101010" => rgb <= "000000";
					when "10011010010101011" => rgb <= "000000";
					when "10011010010101100" => rgb <= "000000";
					when "10011010010101101" => rgb <= "000000";
					when "10011010010101110" => rgb <= "000000";
					when "10011010010101111" => rgb <= "000000";
					when "10011010010110000" => rgb <= "000000";
					when "10011010010110001" => rgb <= "000000";
					when "10011010010110010" => rgb <= "000000";
					when "10011010010110011" => rgb <= "000000";
					when "10011010010110100" => rgb <= "000000";
					when "10011010010110101" => rgb <= "000000";
					when "10011010010110110" => rgb <= "000000";
					when "10011010010110111" => rgb <= "000000";
					when "10011010010111000" => rgb <= "000000";
					when "10011010010111001" => rgb <= "000000";
					when "10011010010111010" => rgb <= "000000";
					when "10011010010111011" => rgb <= "000000";
					when "10011010010111100" => rgb <= "000000";
					when "10011010010111101" => rgb <= "000000";
					when "10011010010111110" => rgb <= "000000";
					when "10011010010111111" => rgb <= "000000";
					when "10011010011000000" => rgb <= "000000";
					when "10011010011000001" => rgb <= "000000";
					when "10011010011000010" => rgb <= "000000";
					when "10011010011000011" => rgb <= "000000";
					when "10011010011000100" => rgb <= "000000";
					when "10011010011000101" => rgb <= "000000";
					when "10011010011000110" => rgb <= "000000";
					when "10011010011000111" => rgb <= "000000";
					when "10011010011001000" => rgb <= "000000";
					when "10011010011001001" => rgb <= "000000";
					when "10011010011001010" => rgb <= "000000";
					when "10011010011001011" => rgb <= "000000";
					when "10011010011001100" => rgb <= "000000";
					when "10011010011001101" => rgb <= "000000";
					when "10011010011001110" => rgb <= "000000";
					when "10011010011001111" => rgb <= "000000";
					when "10011010011010000" => rgb <= "000000";
					when "10011010011010001" => rgb <= "000000";
					when "10011010011010010" => rgb <= "000000";
					when "10011010011010011" => rgb <= "000000";
					when "10011010011010100" => rgb <= "000000";
					when "10011010011010101" => rgb <= "000000";
					when "10011010011010110" => rgb <= "000000";
					when "10011010011010111" => rgb <= "000000";
					when "10011010011011000" => rgb <= "000000";
					when "10011010011011001" => rgb <= "000000";
					when "10011010011011010" => rgb <= "000000";
					when "10011010011011011" => rgb <= "000000";
					when "10011010011011100" => rgb <= "000000";
					when "10011010011011101" => rgb <= "000000";
					when "10011010011011110" => rgb <= "000000";
					when "10011010011011111" => rgb <= "000000";
					when "10011010011100000" => rgb <= "000000";
					when "10011010011100001" => rgb <= "000000";
					when "10011010011100010" => rgb <= "000000";
					when "10011010011100011" => rgb <= "000000";
					when "10011010011100100" => rgb <= "000000";
					when "10011010011100101" => rgb <= "000000";
					when "10011010011100110" => rgb <= "000000";
					when "10011010011100111" => rgb <= "000000";
					when "10011010011101000" => rgb <= "000000";
					when "10011010011101001" => rgb <= "000000";
					when "10011010011101010" => rgb <= "000000";
					when "10011010011101011" => rgb <= "000000";
					when "10011010011101100" => rgb <= "000000";
					when "10011010011101101" => rgb <= "000000";
					when "10011010011101110" => rgb <= "000000";
					when "10011010011101111" => rgb <= "000000";
					when "10011010011110000" => rgb <= "000000";
					when "10011010011110001" => rgb <= "000000";
					when "10011010011110010" => rgb <= "000000";
					when "10011010011110011" => rgb <= "000000";
					when "10011010011110100" => rgb <= "000000";
					when "10011010011110101" => rgb <= "000000";
					when "10011010011110110" => rgb <= "000000";
					when "10011010011110111" => rgb <= "000000";
					when "10011010011111000" => rgb <= "000000";
					when "10011010011111001" => rgb <= "000000";
					when "10011010011111010" => rgb <= "000000";
					when "10011010011111011" => rgb <= "000000";
					when "10011010011111100" => rgb <= "000000";
					when "10011010011111101" => rgb <= "000000";
					when "10011010011111110" => rgb <= "000000";
					when "10011010011111111" => rgb <= "000000";
					when "10011010100000000" => rgb <= "000000";
					when "10011010100000001" => rgb <= "000000";
					when "10011010100000010" => rgb <= "000000";
					when "10011010100000011" => rgb <= "000000";
					when "10011010100000100" => rgb <= "000000";
					when "10011010100000101" => rgb <= "000000";
					when "10011010100000110" => rgb <= "000000";
					when "10011010100000111" => rgb <= "000000";
					when "10011010100001000" => rgb <= "000000";
					when "10011010100001001" => rgb <= "000000";
					when "10011010100001010" => rgb <= "000000";
					when "10011010100001011" => rgb <= "000000";
					when "10011010100001100" => rgb <= "000000";
					when "10011010100001101" => rgb <= "000000";
					when "10011010100001110" => rgb <= "000000";
					when "10011010100001111" => rgb <= "000000";
					when "10011010100010000" => rgb <= "000000";
					when "10011010100010001" => rgb <= "000000";
					when "10011010100010010" => rgb <= "000000";
					when "10011010100010011" => rgb <= "000000";
					when "10011010100010100" => rgb <= "000000";
					when "10011010100010101" => rgb <= "000000";
					when "10011010100010110" => rgb <= "000000";
					when "10011010100010111" => rgb <= "000000";
					when "10011010100011000" => rgb <= "000000";
					when "10011010100011001" => rgb <= "000000";
					when "10011010100011010" => rgb <= "000000";
					when "10011010100011011" => rgb <= "000000";
					when "10011010100011100" => rgb <= "000000";
					when "10011010100011101" => rgb <= "000000";
					when "10011010100011110" => rgb <= "000000";
					when "10011010100011111" => rgb <= "000000";
					when "10011010100100000" => rgb <= "000000";
					when "10011010100100001" => rgb <= "000000";
					when "10011010100100010" => rgb <= "000000";
					when "10011010100100011" => rgb <= "000000";
					when "10011010100100100" => rgb <= "000000";
					when "10011010100100101" => rgb <= "000000";
					when "10011010100100110" => rgb <= "000000";
					when "10011010100100111" => rgb <= "000000";
					when "10011010100101000" => rgb <= "000000";
					when "10011010100101001" => rgb <= "000000";
					when "10011010100101010" => rgb <= "000000";
					when "10011010100101011" => rgb <= "000000";
					when "10011010100101100" => rgb <= "000000";
					when "10011010100101101" => rgb <= "000000";
					when "10011010100101110" => rgb <= "000000";
					when "10011010100101111" => rgb <= "000000";
					when "10011010100110000" => rgb <= "000000";
					when "10011010100110001" => rgb <= "000000";
					when "10011010100110010" => rgb <= "000000";
					when "10011010100110011" => rgb <= "000000";
					when "10011010100110100" => rgb <= "000000";
					when "10011010100110101" => rgb <= "000000";
					when "10011010100110110" => rgb <= "000000";
					when "10011010100110111" => rgb <= "000000";
					when "10011010100111000" => rgb <= "000000";
					when "10011010100111001" => rgb <= "000000";
					when "10011010100111010" => rgb <= "000000";
					when "10011010100111011" => rgb <= "000000";
					when "10011010100111100" => rgb <= "000000";
					when "10011010100111101" => rgb <= "000000";
					when "10011010100111110" => rgb <= "000000";
					when "10011010100111111" => rgb <= "000000";
					when "10011011000000000" => rgb <= "000000";
					when "10011011000000001" => rgb <= "000000";
					when "10011011000000010" => rgb <= "000000";
					when "10011011000000011" => rgb <= "000000";
					when "10011011000000100" => rgb <= "000000";
					when "10011011000000101" => rgb <= "000000";
					when "10011011000000110" => rgb <= "000000";
					when "10011011000000111" => rgb <= "000000";
					when "10011011000001000" => rgb <= "000000";
					when "10011011000001001" => rgb <= "000000";
					when "10011011000001010" => rgb <= "000000";
					when "10011011000001011" => rgb <= "000000";
					when "10011011000001100" => rgb <= "000000";
					when "10011011000001101" => rgb <= "000000";
					when "10011011000001110" => rgb <= "000000";
					when "10011011000001111" => rgb <= "000000";
					when "10011011000010000" => rgb <= "000000";
					when "10011011000010001" => rgb <= "000000";
					when "10011011000010010" => rgb <= "000000";
					when "10011011000010011" => rgb <= "000000";
					when "10011011000010100" => rgb <= "000000";
					when "10011011000010101" => rgb <= "000000";
					when "10011011000010110" => rgb <= "000000";
					when "10011011000010111" => rgb <= "000000";
					when "10011011000011000" => rgb <= "000000";
					when "10011011000011001" => rgb <= "000000";
					when "10011011000011010" => rgb <= "000000";
					when "10011011000011011" => rgb <= "000000";
					when "10011011000011100" => rgb <= "000000";
					when "10011011000011101" => rgb <= "000000";
					when "10011011000011110" => rgb <= "000000";
					when "10011011000011111" => rgb <= "000000";
					when "10011011000100000" => rgb <= "000000";
					when "10011011000100001" => rgb <= "000000";
					when "10011011000100010" => rgb <= "000000";
					when "10011011000100011" => rgb <= "000000";
					when "10011011000100100" => rgb <= "000000";
					when "10011011000100101" => rgb <= "000000";
					when "10011011000100110" => rgb <= "000000";
					when "10011011000100111" => rgb <= "000000";
					when "10011011000101000" => rgb <= "000000";
					when "10011011000101001" => rgb <= "000000";
					when "10011011000101010" => rgb <= "000000";
					when "10011011000101011" => rgb <= "000000";
					when "10011011000101100" => rgb <= "000000";
					when "10011011000101101" => rgb <= "000000";
					when "10011011000101110" => rgb <= "000000";
					when "10011011000101111" => rgb <= "000000";
					when "10011011000110000" => rgb <= "000000";
					when "10011011000110001" => rgb <= "000000";
					when "10011011000110010" => rgb <= "000000";
					when "10011011000110011" => rgb <= "000000";
					when "10011011000110100" => rgb <= "000000";
					when "10011011000110101" => rgb <= "000000";
					when "10011011000110110" => rgb <= "000000";
					when "10011011000110111" => rgb <= "000000";
					when "10011011000111000" => rgb <= "000000";
					when "10011011000111001" => rgb <= "000000";
					when "10011011000111010" => rgb <= "000000";
					when "10011011000111011" => rgb <= "000000";
					when "10011011000111100" => rgb <= "000000";
					when "10011011000111101" => rgb <= "000000";
					when "10011011000111110" => rgb <= "000000";
					when "10011011000111111" => rgb <= "000000";
					when "10011011001000000" => rgb <= "000000";
					when "10011011001000001" => rgb <= "000000";
					when "10011011001000010" => rgb <= "000000";
					when "10011011001000011" => rgb <= "000000";
					when "10011011001000100" => rgb <= "000000";
					when "10011011001000101" => rgb <= "000000";
					when "10011011001000110" => rgb <= "000000";
					when "10011011001000111" => rgb <= "000000";
					when "10011011001001000" => rgb <= "000000";
					when "10011011001001001" => rgb <= "000000";
					when "10011011001001010" => rgb <= "000000";
					when "10011011001001011" => rgb <= "000000";
					when "10011011001001100" => rgb <= "000000";
					when "10011011001001101" => rgb <= "000000";
					when "10011011001001110" => rgb <= "000000";
					when "10011011001001111" => rgb <= "000000";
					when "10011011001010000" => rgb <= "000000";
					when "10011011001010001" => rgb <= "000000";
					when "10011011001010010" => rgb <= "000000";
					when "10011011001010011" => rgb <= "000000";
					when "10011011001010100" => rgb <= "000000";
					when "10011011001010101" => rgb <= "000000";
					when "10011011001010110" => rgb <= "000000";
					when "10011011001010111" => rgb <= "000000";
					when "10011011001011000" => rgb <= "000000";
					when "10011011001011001" => rgb <= "000000";
					when "10011011001011010" => rgb <= "000000";
					when "10011011001011011" => rgb <= "000000";
					when "10011011001011100" => rgb <= "000000";
					when "10011011001011101" => rgb <= "000000";
					when "10011011001011110" => rgb <= "000000";
					when "10011011001011111" => rgb <= "000000";
					when "10011011001100000" => rgb <= "000000";
					when "10011011001100001" => rgb <= "000000";
					when "10011011001100010" => rgb <= "000000";
					when "10011011001100011" => rgb <= "000000";
					when "10011011001100100" => rgb <= "000000";
					when "10011011001100101" => rgb <= "000000";
					when "10011011001100110" => rgb <= "000000";
					when "10011011001100111" => rgb <= "000000";
					when "10011011001101000" => rgb <= "000000";
					when "10011011001101001" => rgb <= "000000";
					when "10011011001101010" => rgb <= "000000";
					when "10011011001101011" => rgb <= "000000";
					when "10011011001101100" => rgb <= "000000";
					when "10011011001101101" => rgb <= "000000";
					when "10011011001101110" => rgb <= "000000";
					when "10011011001101111" => rgb <= "000000";
					when "10011011001110000" => rgb <= "000000";
					when "10011011001110001" => rgb <= "000000";
					when "10011011001110010" => rgb <= "000000";
					when "10011011001110011" => rgb <= "000000";
					when "10011011001110100" => rgb <= "000000";
					when "10011011001110101" => rgb <= "000000";
					when "10011011001110110" => rgb <= "000000";
					when "10011011001110111" => rgb <= "000000";
					when "10011011001111000" => rgb <= "000000";
					when "10011011001111001" => rgb <= "000000";
					when "10011011001111010" => rgb <= "000000";
					when "10011011001111011" => rgb <= "000000";
					when "10011011001111100" => rgb <= "000000";
					when "10011011001111101" => rgb <= "000000";
					when "10011011001111110" => rgb <= "000000";
					when "10011011001111111" => rgb <= "000000";
					when "10011011010000000" => rgb <= "000000";
					when "10011011010000001" => rgb <= "000000";
					when "10011011010000010" => rgb <= "000000";
					when "10011011010000011" => rgb <= "000000";
					when "10011011010000100" => rgb <= "000000";
					when "10011011010000101" => rgb <= "000000";
					when "10011011010000110" => rgb <= "000000";
					when "10011011010000111" => rgb <= "000000";
					when "10011011010001000" => rgb <= "000000";
					when "10011011010001001" => rgb <= "000000";
					when "10011011010001010" => rgb <= "000000";
					when "10011011010001011" => rgb <= "000000";
					when "10011011010001100" => rgb <= "000000";
					when "10011011010001101" => rgb <= "000000";
					when "10011011010001110" => rgb <= "000000";
					when "10011011010001111" => rgb <= "000000";
					when "10011011010010000" => rgb <= "000000";
					when "10011011010010001" => rgb <= "000000";
					when "10011011010010010" => rgb <= "000000";
					when "10011011010010011" => rgb <= "000000";
					when "10011011010010100" => rgb <= "000000";
					when "10011011010010101" => rgb <= "000000";
					when "10011011010010110" => rgb <= "000000";
					when "10011011010010111" => rgb <= "000000";
					when "10011011010011000" => rgb <= "000000";
					when "10011011010011001" => rgb <= "000000";
					when "10011011010011010" => rgb <= "000000";
					when "10011011010011011" => rgb <= "000000";
					when "10011011010011100" => rgb <= "000000";
					when "10011011010011101" => rgb <= "000000";
					when "10011011010011110" => rgb <= "000000";
					when "10011011010011111" => rgb <= "000000";
					when "10011011010100000" => rgb <= "000000";
					when "10011011010100001" => rgb <= "000000";
					when "10011011010100010" => rgb <= "000000";
					when "10011011010100011" => rgb <= "000000";
					when "10011011010100100" => rgb <= "000000";
					when "10011011010100101" => rgb <= "000000";
					when "10011011010100110" => rgb <= "000000";
					when "10011011010100111" => rgb <= "000000";
					when "10011011010101000" => rgb <= "000000";
					when "10011011010101001" => rgb <= "000000";
					when "10011011010101010" => rgb <= "000000";
					when "10011011010101011" => rgb <= "000000";
					when "10011011010101100" => rgb <= "000000";
					when "10011011010101101" => rgb <= "000000";
					when "10011011010101110" => rgb <= "000000";
					when "10011011010101111" => rgb <= "000000";
					when "10011011010110000" => rgb <= "000000";
					when "10011011010110001" => rgb <= "000000";
					when "10011011010110010" => rgb <= "000000";
					when "10011011010110011" => rgb <= "000000";
					when "10011011010110100" => rgb <= "000000";
					when "10011011010110101" => rgb <= "000000";
					when "10011011010110110" => rgb <= "000000";
					when "10011011010110111" => rgb <= "000000";
					when "10011011010111000" => rgb <= "000000";
					when "10011011010111001" => rgb <= "000000";
					when "10011011010111010" => rgb <= "000000";
					when "10011011010111011" => rgb <= "000000";
					when "10011011010111100" => rgb <= "000000";
					when "10011011010111101" => rgb <= "000000";
					when "10011011010111110" => rgb <= "000000";
					when "10011011010111111" => rgb <= "000000";
					when "10011011011000000" => rgb <= "000000";
					when "10011011011000001" => rgb <= "000000";
					when "10011011011000010" => rgb <= "000000";
					when "10011011011000011" => rgb <= "000000";
					when "10011011011000100" => rgb <= "000000";
					when "10011011011000101" => rgb <= "000000";
					when "10011011011000110" => rgb <= "000000";
					when "10011011011000111" => rgb <= "000000";
					when "10011011011001000" => rgb <= "000000";
					when "10011011011001001" => rgb <= "000000";
					when "10011011011001010" => rgb <= "000000";
					when "10011011011001011" => rgb <= "000000";
					when "10011011011001100" => rgb <= "000000";
					when "10011011011001101" => rgb <= "000000";
					when "10011011011001110" => rgb <= "000000";
					when "10011011011001111" => rgb <= "000000";
					when "10011011011010000" => rgb <= "000000";
					when "10011011011010001" => rgb <= "000000";
					when "10011011011010010" => rgb <= "000000";
					when "10011011011010011" => rgb <= "000000";
					when "10011011011010100" => rgb <= "000000";
					when "10011011011010101" => rgb <= "000000";
					when "10011011011010110" => rgb <= "000000";
					when "10011011011010111" => rgb <= "000000";
					when "10011011011011000" => rgb <= "000000";
					when "10011011011011001" => rgb <= "000000";
					when "10011011011011010" => rgb <= "000000";
					when "10011011011011011" => rgb <= "000000";
					when "10011011011011100" => rgb <= "000000";
					when "10011011011011101" => rgb <= "000000";
					when "10011011011011110" => rgb <= "000000";
					when "10011011011011111" => rgb <= "000000";
					when "10011011011100000" => rgb <= "000000";
					when "10011011011100001" => rgb <= "000000";
					when "10011011011100010" => rgb <= "000000";
					when "10011011011100011" => rgb <= "000000";
					when "10011011011100100" => rgb <= "000000";
					when "10011011011100101" => rgb <= "000000";
					when "10011011011100110" => rgb <= "000000";
					when "10011011011100111" => rgb <= "000000";
					when "10011011011101000" => rgb <= "000000";
					when "10011011011101001" => rgb <= "000000";
					when "10011011011101010" => rgb <= "000000";
					when "10011011011101011" => rgb <= "000000";
					when "10011011011101100" => rgb <= "000000";
					when "10011011011101101" => rgb <= "000000";
					when "10011011011101110" => rgb <= "000000";
					when "10011011011101111" => rgb <= "000000";
					when "10011011011110000" => rgb <= "000000";
					when "10011011011110001" => rgb <= "000000";
					when "10011011011110010" => rgb <= "000000";
					when "10011011011110011" => rgb <= "000000";
					when "10011011011110100" => rgb <= "000000";
					when "10011011011110101" => rgb <= "000000";
					when "10011011011110110" => rgb <= "000000";
					when "10011011011110111" => rgb <= "000000";
					when "10011011011111000" => rgb <= "000000";
					when "10011011011111001" => rgb <= "000000";
					when "10011011011111010" => rgb <= "000000";
					when "10011011011111011" => rgb <= "000000";
					when "10011011011111100" => rgb <= "000000";
					when "10011011011111101" => rgb <= "000000";
					when "10011011011111110" => rgb <= "000000";
					when "10011011011111111" => rgb <= "000000";
					when "10011011100000000" => rgb <= "000000";
					when "10011011100000001" => rgb <= "000000";
					when "10011011100000010" => rgb <= "000000";
					when "10011011100000011" => rgb <= "000000";
					when "10011011100000100" => rgb <= "000000";
					when "10011011100000101" => rgb <= "000000";
					when "10011011100000110" => rgb <= "000000";
					when "10011011100000111" => rgb <= "000000";
					when "10011011100001000" => rgb <= "000000";
					when "10011011100001001" => rgb <= "000000";
					when "10011011100001010" => rgb <= "000000";
					when "10011011100001011" => rgb <= "000000";
					when "10011011100001100" => rgb <= "000000";
					when "10011011100001101" => rgb <= "000000";
					when "10011011100001110" => rgb <= "000000";
					when "10011011100001111" => rgb <= "000000";
					when "10011011100010000" => rgb <= "000000";
					when "10011011100010001" => rgb <= "000000";
					when "10011011100010010" => rgb <= "000000";
					when "10011011100010011" => rgb <= "000000";
					when "10011011100010100" => rgb <= "000000";
					when "10011011100010101" => rgb <= "000000";
					when "10011011100010110" => rgb <= "000000";
					when "10011011100010111" => rgb <= "000000";
					when "10011011100011000" => rgb <= "000000";
					when "10011011100011001" => rgb <= "000000";
					when "10011011100011010" => rgb <= "000000";
					when "10011011100011011" => rgb <= "000000";
					when "10011011100011100" => rgb <= "000000";
					when "10011011100011101" => rgb <= "000000";
					when "10011011100011110" => rgb <= "000000";
					when "10011011100011111" => rgb <= "000000";
					when "10011011100100000" => rgb <= "000000";
					when "10011011100100001" => rgb <= "000000";
					when "10011011100100010" => rgb <= "000000";
					when "10011011100100011" => rgb <= "000000";
					when "10011011100100100" => rgb <= "000000";
					when "10011011100100101" => rgb <= "000000";
					when "10011011100100110" => rgb <= "000000";
					when "10011011100100111" => rgb <= "000000";
					when "10011011100101000" => rgb <= "000000";
					when "10011011100101001" => rgb <= "000000";
					when "10011011100101010" => rgb <= "000000";
					when "10011011100101011" => rgb <= "000000";
					when "10011011100101100" => rgb <= "000000";
					when "10011011100101101" => rgb <= "000000";
					when "10011011100101110" => rgb <= "000000";
					when "10011011100101111" => rgb <= "000000";
					when "10011011100110000" => rgb <= "000000";
					when "10011011100110001" => rgb <= "000000";
					when "10011011100110010" => rgb <= "000000";
					when "10011011100110011" => rgb <= "000000";
					when "10011011100110100" => rgb <= "000000";
					when "10011011100110101" => rgb <= "000000";
					when "10011011100110110" => rgb <= "000000";
					when "10011011100110111" => rgb <= "000000";
					when "10011011100111000" => rgb <= "000000";
					when "10011011100111001" => rgb <= "000000";
					when "10011011100111010" => rgb <= "000000";
					when "10011011100111011" => rgb <= "000000";
					when "10011011100111100" => rgb <= "000000";
					when "10011011100111101" => rgb <= "000000";
					when "10011011100111110" => rgb <= "000000";
					when "10011011100111111" => rgb <= "000000";
					when "10011100000000000" => rgb <= "000000";
					when "10011100000000001" => rgb <= "000000";
					when "10011100000000010" => rgb <= "000000";
					when "10011100000000011" => rgb <= "000000";
					when "10011100000000100" => rgb <= "000000";
					when "10011100000000101" => rgb <= "000000";
					when "10011100000000110" => rgb <= "000000";
					when "10011100000000111" => rgb <= "000000";
					when "10011100000001000" => rgb <= "000000";
					when "10011100000001001" => rgb <= "000000";
					when "10011100000001010" => rgb <= "000000";
					when "10011100000001011" => rgb <= "000000";
					when "10011100000001100" => rgb <= "000000";
					when "10011100000001101" => rgb <= "000000";
					when "10011100000001110" => rgb <= "000000";
					when "10011100000001111" => rgb <= "000000";
					when "10011100000010000" => rgb <= "000000";
					when "10011100000010001" => rgb <= "000000";
					when "10011100000010010" => rgb <= "000000";
					when "10011100000010011" => rgb <= "000000";
					when "10011100000010100" => rgb <= "000000";
					when "10011100000010101" => rgb <= "000000";
					when "10011100000010110" => rgb <= "000000";
					when "10011100000010111" => rgb <= "000000";
					when "10011100000011000" => rgb <= "000000";
					when "10011100000011001" => rgb <= "000000";
					when "10011100000011010" => rgb <= "000000";
					when "10011100000011011" => rgb <= "000000";
					when "10011100000011100" => rgb <= "000000";
					when "10011100000011101" => rgb <= "000000";
					when "10011100000011110" => rgb <= "000000";
					when "10011100000011111" => rgb <= "000000";
					when "10011100000100000" => rgb <= "000000";
					when "10011100000100001" => rgb <= "000000";
					when "10011100000100010" => rgb <= "000000";
					when "10011100000100011" => rgb <= "000000";
					when "10011100000100100" => rgb <= "000000";
					when "10011100000100101" => rgb <= "000000";
					when "10011100000100110" => rgb <= "000000";
					when "10011100000100111" => rgb <= "000000";
					when "10011100000101000" => rgb <= "000000";
					when "10011100000101001" => rgb <= "000000";
					when "10011100000101010" => rgb <= "000000";
					when "10011100000101011" => rgb <= "000000";
					when "10011100000101100" => rgb <= "000000";
					when "10011100000101101" => rgb <= "000000";
					when "10011100000101110" => rgb <= "000000";
					when "10011100000101111" => rgb <= "000000";
					when "10011100000110000" => rgb <= "000000";
					when "10011100000110001" => rgb <= "000000";
					when "10011100000110010" => rgb <= "000000";
					when "10011100000110011" => rgb <= "000000";
					when "10011100000110100" => rgb <= "000000";
					when "10011100000110101" => rgb <= "000000";
					when "10011100000110110" => rgb <= "000000";
					when "10011100000110111" => rgb <= "000000";
					when "10011100000111000" => rgb <= "000000";
					when "10011100000111001" => rgb <= "000000";
					when "10011100000111010" => rgb <= "000000";
					when "10011100000111011" => rgb <= "000000";
					when "10011100000111100" => rgb <= "000000";
					when "10011100000111101" => rgb <= "000000";
					when "10011100000111110" => rgb <= "000000";
					when "10011100000111111" => rgb <= "000000";
					when "10011100001000000" => rgb <= "000000";
					when "10011100001000001" => rgb <= "000000";
					when "10011100001000010" => rgb <= "000000";
					when "10011100001000011" => rgb <= "000000";
					when "10011100001000100" => rgb <= "000000";
					when "10011100001000101" => rgb <= "000000";
					when "10011100001000110" => rgb <= "000000";
					when "10011100001000111" => rgb <= "000000";
					when "10011100001001000" => rgb <= "000000";
					when "10011100001001001" => rgb <= "000000";
					when "10011100001001010" => rgb <= "000000";
					when "10011100001001011" => rgb <= "000000";
					when "10011100001001100" => rgb <= "000000";
					when "10011100001001101" => rgb <= "000000";
					when "10011100001001110" => rgb <= "000000";
					when "10011100001001111" => rgb <= "000000";
					when "10011100001010000" => rgb <= "000000";
					when "10011100001010001" => rgb <= "000000";
					when "10011100001010010" => rgb <= "000000";
					when "10011100001010011" => rgb <= "000000";
					when "10011100001010100" => rgb <= "000000";
					when "10011100001010101" => rgb <= "000000";
					when "10011100001010110" => rgb <= "000000";
					when "10011100001010111" => rgb <= "000000";
					when "10011100001011000" => rgb <= "000000";
					when "10011100001011001" => rgb <= "000000";
					when "10011100001011010" => rgb <= "000000";
					when "10011100001011011" => rgb <= "000000";
					when "10011100001011100" => rgb <= "000000";
					when "10011100001011101" => rgb <= "000000";
					when "10011100001011110" => rgb <= "000000";
					when "10011100001011111" => rgb <= "000000";
					when "10011100001100000" => rgb <= "000000";
					when "10011100001100001" => rgb <= "000000";
					when "10011100001100010" => rgb <= "000000";
					when "10011100001100011" => rgb <= "000000";
					when "10011100001100100" => rgb <= "000000";
					when "10011100001100101" => rgb <= "000000";
					when "10011100001100110" => rgb <= "000000";
					when "10011100001100111" => rgb <= "000000";
					when "10011100001101000" => rgb <= "000000";
					when "10011100001101001" => rgb <= "000000";
					when "10011100001101010" => rgb <= "000000";
					when "10011100001101011" => rgb <= "000000";
					when "10011100001101100" => rgb <= "000000";
					when "10011100001101101" => rgb <= "000000";
					when "10011100001101110" => rgb <= "000000";
					when "10011100001101111" => rgb <= "000000";
					when "10011100001110000" => rgb <= "000000";
					when "10011100001110001" => rgb <= "000000";
					when "10011100001110010" => rgb <= "000000";
					when "10011100001110011" => rgb <= "000000";
					when "10011100001110100" => rgb <= "000000";
					when "10011100001110101" => rgb <= "000000";
					when "10011100001110110" => rgb <= "000000";
					when "10011100001110111" => rgb <= "000000";
					when "10011100001111000" => rgb <= "000000";
					when "10011100001111001" => rgb <= "000000";
					when "10011100001111010" => rgb <= "000000";
					when "10011100001111011" => rgb <= "000000";
					when "10011100001111100" => rgb <= "000000";
					when "10011100001111101" => rgb <= "000000";
					when "10011100001111110" => rgb <= "000000";
					when "10011100001111111" => rgb <= "000000";
					when "10011100010000000" => rgb <= "000000";
					when "10011100010000001" => rgb <= "000000";
					when "10011100010000010" => rgb <= "000000";
					when "10011100010000011" => rgb <= "000000";
					when "10011100010000100" => rgb <= "000000";
					when "10011100010000101" => rgb <= "000000";
					when "10011100010000110" => rgb <= "000000";
					when "10011100010000111" => rgb <= "000000";
					when "10011100010001000" => rgb <= "000000";
					when "10011100010001001" => rgb <= "000000";
					when "10011100010001010" => rgb <= "000000";
					when "10011100010001011" => rgb <= "000000";
					when "10011100010001100" => rgb <= "000000";
					when "10011100010001101" => rgb <= "000000";
					when "10011100010001110" => rgb <= "000000";
					when "10011100010001111" => rgb <= "000000";
					when "10011100010010000" => rgb <= "000000";
					when "10011100010010001" => rgb <= "000000";
					when "10011100010010010" => rgb <= "000000";
					when "10011100010010011" => rgb <= "000000";
					when "10011100010010100" => rgb <= "000000";
					when "10011100010010101" => rgb <= "000000";
					when "10011100010010110" => rgb <= "000000";
					when "10011100010010111" => rgb <= "000000";
					when "10011100010011000" => rgb <= "000000";
					when "10011100010011001" => rgb <= "000000";
					when "10011100010011010" => rgb <= "000000";
					when "10011100010011011" => rgb <= "000000";
					when "10011100010011100" => rgb <= "000000";
					when "10011100010011101" => rgb <= "000000";
					when "10011100010011110" => rgb <= "000000";
					when "10011100010011111" => rgb <= "000000";
					when "10011100010100000" => rgb <= "000000";
					when "10011100010100001" => rgb <= "000000";
					when "10011100010100010" => rgb <= "000000";
					when "10011100010100011" => rgb <= "000000";
					when "10011100010100100" => rgb <= "000000";
					when "10011100010100101" => rgb <= "000000";
					when "10011100010100110" => rgb <= "000000";
					when "10011100010100111" => rgb <= "000000";
					when "10011100010101000" => rgb <= "000000";
					when "10011100010101001" => rgb <= "000000";
					when "10011100010101010" => rgb <= "000000";
					when "10011100010101011" => rgb <= "000000";
					when "10011100010101100" => rgb <= "000000";
					when "10011100010101101" => rgb <= "000000";
					when "10011100010101110" => rgb <= "000000";
					when "10011100010101111" => rgb <= "000000";
					when "10011100010110000" => rgb <= "000000";
					when "10011100010110001" => rgb <= "000000";
					when "10011100010110010" => rgb <= "000000";
					when "10011100010110011" => rgb <= "000000";
					when "10011100010110100" => rgb <= "000000";
					when "10011100010110101" => rgb <= "000000";
					when "10011100010110110" => rgb <= "000000";
					when "10011100010110111" => rgb <= "000000";
					when "10011100010111000" => rgb <= "000000";
					when "10011100010111001" => rgb <= "000000";
					when "10011100010111010" => rgb <= "000000";
					when "10011100010111011" => rgb <= "000000";
					when "10011100010111100" => rgb <= "000000";
					when "10011100010111101" => rgb <= "000000";
					when "10011100010111110" => rgb <= "000000";
					when "10011100010111111" => rgb <= "000000";
					when "10011100011000000" => rgb <= "000000";
					when "10011100011000001" => rgb <= "000000";
					when "10011100011000010" => rgb <= "000000";
					when "10011100011000011" => rgb <= "000000";
					when "10011100011000100" => rgb <= "000000";
					when "10011100011000101" => rgb <= "000000";
					when "10011100011000110" => rgb <= "000000";
					when "10011100011000111" => rgb <= "000000";
					when "10011100011001000" => rgb <= "000000";
					when "10011100011001001" => rgb <= "000000";
					when "10011100011001010" => rgb <= "000000";
					when "10011100011001011" => rgb <= "000000";
					when "10011100011001100" => rgb <= "000000";
					when "10011100011001101" => rgb <= "000000";
					when "10011100011001110" => rgb <= "000000";
					when "10011100011001111" => rgb <= "000000";
					when "10011100011010000" => rgb <= "000000";
					when "10011100011010001" => rgb <= "000000";
					when "10011100011010010" => rgb <= "000000";
					when "10011100011010011" => rgb <= "000000";
					when "10011100011010100" => rgb <= "000000";
					when "10011100011010101" => rgb <= "000000";
					when "10011100011010110" => rgb <= "000000";
					when "10011100011010111" => rgb <= "000000";
					when "10011100011011000" => rgb <= "000000";
					when "10011100011011001" => rgb <= "000000";
					when "10011100011011010" => rgb <= "000000";
					when "10011100011011011" => rgb <= "000000";
					when "10011100011011100" => rgb <= "000000";
					when "10011100011011101" => rgb <= "000000";
					when "10011100011011110" => rgb <= "000000";
					when "10011100011011111" => rgb <= "000000";
					when "10011100011100000" => rgb <= "000000";
					when "10011100011100001" => rgb <= "000000";
					when "10011100011100010" => rgb <= "000000";
					when "10011100011100011" => rgb <= "000000";
					when "10011100011100100" => rgb <= "000000";
					when "10011100011100101" => rgb <= "000000";
					when "10011100011100110" => rgb <= "000000";
					when "10011100011100111" => rgb <= "000000";
					when "10011100011101000" => rgb <= "000000";
					when "10011100011101001" => rgb <= "000000";
					when "10011100011101010" => rgb <= "000000";
					when "10011100011101011" => rgb <= "000000";
					when "10011100011101100" => rgb <= "000000";
					when "10011100011101101" => rgb <= "000000";
					when "10011100011101110" => rgb <= "000000";
					when "10011100011101111" => rgb <= "000000";
					when "10011100011110000" => rgb <= "000000";
					when "10011100011110001" => rgb <= "000000";
					when "10011100011110010" => rgb <= "000000";
					when "10011100011110011" => rgb <= "000000";
					when "10011100011110100" => rgb <= "000000";
					when "10011100011110101" => rgb <= "000000";
					when "10011100011110110" => rgb <= "000000";
					when "10011100011110111" => rgb <= "000000";
					when "10011100011111000" => rgb <= "000000";
					when "10011100011111001" => rgb <= "000000";
					when "10011100011111010" => rgb <= "000000";
					when "10011100011111011" => rgb <= "000000";
					when "10011100011111100" => rgb <= "000000";
					when "10011100011111101" => rgb <= "000000";
					when "10011100011111110" => rgb <= "000000";
					when "10011100011111111" => rgb <= "000000";
					when "10011100100000000" => rgb <= "000000";
					when "10011100100000001" => rgb <= "000000";
					when "10011100100000010" => rgb <= "000000";
					when "10011100100000011" => rgb <= "000000";
					when "10011100100000100" => rgb <= "000000";
					when "10011100100000101" => rgb <= "000000";
					when "10011100100000110" => rgb <= "000000";
					when "10011100100000111" => rgb <= "000000";
					when "10011100100001000" => rgb <= "000000";
					when "10011100100001001" => rgb <= "000000";
					when "10011100100001010" => rgb <= "000000";
					when "10011100100001011" => rgb <= "000000";
					when "10011100100001100" => rgb <= "000000";
					when "10011100100001101" => rgb <= "000000";
					when "10011100100001110" => rgb <= "000000";
					when "10011100100001111" => rgb <= "000000";
					when "10011100100010000" => rgb <= "000000";
					when "10011100100010001" => rgb <= "000000";
					when "10011100100010010" => rgb <= "000000";
					when "10011100100010011" => rgb <= "000000";
					when "10011100100010100" => rgb <= "000000";
					when "10011100100010101" => rgb <= "000000";
					when "10011100100010110" => rgb <= "000000";
					when "10011100100010111" => rgb <= "000000";
					when "10011100100011000" => rgb <= "000000";
					when "10011100100011001" => rgb <= "000000";
					when "10011100100011010" => rgb <= "000000";
					when "10011100100011011" => rgb <= "000000";
					when "10011100100011100" => rgb <= "000000";
					when "10011100100011101" => rgb <= "000000";
					when "10011100100011110" => rgb <= "000000";
					when "10011100100011111" => rgb <= "000000";
					when "10011100100100000" => rgb <= "000000";
					when "10011100100100001" => rgb <= "000000";
					when "10011100100100010" => rgb <= "000000";
					when "10011100100100011" => rgb <= "000000";
					when "10011100100100100" => rgb <= "000000";
					when "10011100100100101" => rgb <= "000000";
					when "10011100100100110" => rgb <= "000000";
					when "10011100100100111" => rgb <= "000000";
					when "10011100100101000" => rgb <= "000000";
					when "10011100100101001" => rgb <= "000000";
					when "10011100100101010" => rgb <= "000000";
					when "10011100100101011" => rgb <= "000000";
					when "10011100100101100" => rgb <= "000000";
					when "10011100100101101" => rgb <= "000000";
					when "10011100100101110" => rgb <= "000000";
					when "10011100100101111" => rgb <= "000000";
					when "10011100100110000" => rgb <= "000000";
					when "10011100100110001" => rgb <= "000000";
					when "10011100100110010" => rgb <= "000000";
					when "10011100100110011" => rgb <= "000000";
					when "10011100100110100" => rgb <= "000000";
					when "10011100100110101" => rgb <= "000000";
					when "10011100100110110" => rgb <= "000000";
					when "10011100100110111" => rgb <= "000000";
					when "10011100100111000" => rgb <= "000000";
					when "10011100100111001" => rgb <= "000000";
					when "10011100100111010" => rgb <= "000000";
					when "10011100100111011" => rgb <= "000000";
					when "10011100100111100" => rgb <= "000000";
					when "10011100100111101" => rgb <= "000000";
					when "10011100100111110" => rgb <= "000000";
					when "10011100100111111" => rgb <= "000000";
					when "10011101000000000" => rgb <= "000000";
					when "10011101000000001" => rgb <= "000000";
					when "10011101000000010" => rgb <= "000000";
					when "10011101000000011" => rgb <= "000000";
					when "10011101000000100" => rgb <= "000000";
					when "10011101000000101" => rgb <= "000000";
					when "10011101000000110" => rgb <= "000000";
					when "10011101000000111" => rgb <= "000000";
					when "10011101000001000" => rgb <= "000000";
					when "10011101000001001" => rgb <= "000000";
					when "10011101000001010" => rgb <= "000000";
					when "10011101000001011" => rgb <= "000000";
					when "10011101000001100" => rgb <= "000000";
					when "10011101000001101" => rgb <= "000000";
					when "10011101000001110" => rgb <= "000000";
					when "10011101000001111" => rgb <= "000000";
					when "10011101000010000" => rgb <= "000000";
					when "10011101000010001" => rgb <= "000000";
					when "10011101000010010" => rgb <= "000000";
					when "10011101000010011" => rgb <= "000000";
					when "10011101000010100" => rgb <= "000000";
					when "10011101000010101" => rgb <= "000000";
					when "10011101000010110" => rgb <= "000000";
					when "10011101000010111" => rgb <= "000000";
					when "10011101000011000" => rgb <= "000000";
					when "10011101000011001" => rgb <= "000000";
					when "10011101000011010" => rgb <= "000000";
					when "10011101000011011" => rgb <= "000000";
					when "10011101000011100" => rgb <= "000000";
					when "10011101000011101" => rgb <= "000000";
					when "10011101000011110" => rgb <= "000000";
					when "10011101000011111" => rgb <= "000000";
					when "10011101000100000" => rgb <= "000000";
					when "10011101000100001" => rgb <= "000000";
					when "10011101000100010" => rgb <= "000000";
					when "10011101000100011" => rgb <= "000000";
					when "10011101000100100" => rgb <= "000000";
					when "10011101000100101" => rgb <= "000000";
					when "10011101000100110" => rgb <= "000000";
					when "10011101000100111" => rgb <= "000000";
					when "10011101000101000" => rgb <= "000000";
					when "10011101000101001" => rgb <= "000000";
					when "10011101000101010" => rgb <= "000000";
					when "10011101000101011" => rgb <= "000000";
					when "10011101000101100" => rgb <= "000000";
					when "10011101000101101" => rgb <= "000000";
					when "10011101000101110" => rgb <= "000000";
					when "10011101000101111" => rgb <= "000000";
					when "10011101000110000" => rgb <= "000000";
					when "10011101000110001" => rgb <= "000000";
					when "10011101000110010" => rgb <= "000000";
					when "10011101000110011" => rgb <= "000000";
					when "10011101000110100" => rgb <= "000000";
					when "10011101000110101" => rgb <= "000000";
					when "10011101000110110" => rgb <= "000000";
					when "10011101000110111" => rgb <= "000000";
					when "10011101000111000" => rgb <= "000000";
					when "10011101000111001" => rgb <= "000000";
					when "10011101000111010" => rgb <= "000000";
					when "10011101000111011" => rgb <= "000000";
					when "10011101000111100" => rgb <= "000000";
					when "10011101000111101" => rgb <= "000000";
					when "10011101000111110" => rgb <= "000000";
					when "10011101000111111" => rgb <= "000000";
					when "10011101001000000" => rgb <= "000000";
					when "10011101001000001" => rgb <= "000000";
					when "10011101001000010" => rgb <= "000000";
					when "10011101001000011" => rgb <= "000000";
					when "10011101001000100" => rgb <= "000000";
					when "10011101001000101" => rgb <= "000000";
					when "10011101001000110" => rgb <= "000000";
					when "10011101001000111" => rgb <= "000000";
					when "10011101001001000" => rgb <= "000000";
					when "10011101001001001" => rgb <= "000000";
					when "10011101001001010" => rgb <= "000000";
					when "10011101001001011" => rgb <= "000000";
					when "10011101001001100" => rgb <= "000000";
					when "10011101001001101" => rgb <= "000000";
					when "10011101001001110" => rgb <= "000000";
					when "10011101001001111" => rgb <= "000000";
					when "10011101001010000" => rgb <= "000000";
					when "10011101001010001" => rgb <= "000000";
					when "10011101001010010" => rgb <= "000000";
					when "10011101001010011" => rgb <= "000000";
					when "10011101001010100" => rgb <= "000000";
					when "10011101001010101" => rgb <= "000000";
					when "10011101001010110" => rgb <= "000000";
					when "10011101001010111" => rgb <= "000000";
					when "10011101001011000" => rgb <= "000000";
					when "10011101001011001" => rgb <= "000000";
					when "10011101001011010" => rgb <= "000000";
					when "10011101001011011" => rgb <= "000000";
					when "10011101001011100" => rgb <= "000000";
					when "10011101001011101" => rgb <= "000000";
					when "10011101001011110" => rgb <= "000000";
					when "10011101001011111" => rgb <= "000000";
					when "10011101001100000" => rgb <= "000000";
					when "10011101001100001" => rgb <= "000000";
					when "10011101001100010" => rgb <= "000000";
					when "10011101001100011" => rgb <= "000000";
					when "10011101001100100" => rgb <= "000000";
					when "10011101001100101" => rgb <= "000000";
					when "10011101001100110" => rgb <= "000000";
					when "10011101001100111" => rgb <= "000000";
					when "10011101001101000" => rgb <= "000000";
					when "10011101001101001" => rgb <= "000000";
					when "10011101001101010" => rgb <= "000000";
					when "10011101001101011" => rgb <= "000000";
					when "10011101001101100" => rgb <= "000000";
					when "10011101001101101" => rgb <= "000000";
					when "10011101001101110" => rgb <= "000000";
					when "10011101001101111" => rgb <= "000000";
					when "10011101001110000" => rgb <= "000000";
					when "10011101001110001" => rgb <= "000000";
					when "10011101001110010" => rgb <= "000000";
					when "10011101001110011" => rgb <= "000000";
					when "10011101001110100" => rgb <= "000000";
					when "10011101001110101" => rgb <= "000000";
					when "10011101001110110" => rgb <= "000000";
					when "10011101001110111" => rgb <= "000000";
					when "10011101001111000" => rgb <= "000000";
					when "10011101001111001" => rgb <= "000000";
					when "10011101001111010" => rgb <= "000000";
					when "10011101001111011" => rgb <= "000000";
					when "10011101001111100" => rgb <= "000000";
					when "10011101001111101" => rgb <= "000000";
					when "10011101001111110" => rgb <= "000000";
					when "10011101001111111" => rgb <= "000000";
					when "10011101010000000" => rgb <= "000000";
					when "10011101010000001" => rgb <= "000000";
					when "10011101010000010" => rgb <= "000000";
					when "10011101010000011" => rgb <= "000000";
					when "10011101010000100" => rgb <= "000000";
					when "10011101010000101" => rgb <= "000000";
					when "10011101010000110" => rgb <= "000000";
					when "10011101010000111" => rgb <= "000000";
					when "10011101010001000" => rgb <= "000000";
					when "10011101010001001" => rgb <= "000000";
					when "10011101010001010" => rgb <= "000000";
					when "10011101010001011" => rgb <= "000000";
					when "10011101010001100" => rgb <= "000000";
					when "10011101010001101" => rgb <= "000000";
					when "10011101010001110" => rgb <= "000000";
					when "10011101010001111" => rgb <= "000000";
					when "10011101010010000" => rgb <= "000000";
					when "10011101010010001" => rgb <= "000000";
					when "10011101010010010" => rgb <= "000000";
					when "10011101010010011" => rgb <= "000000";
					when "10011101010010100" => rgb <= "000000";
					when "10011101010010101" => rgb <= "000000";
					when "10011101010010110" => rgb <= "000000";
					when "10011101010010111" => rgb <= "000000";
					when "10011101010011000" => rgb <= "000000";
					when "10011101010011001" => rgb <= "000000";
					when "10011101010011010" => rgb <= "000000";
					when "10011101010011011" => rgb <= "000000";
					when "10011101010011100" => rgb <= "000000";
					when "10011101010011101" => rgb <= "000000";
					when "10011101010011110" => rgb <= "000000";
					when "10011101010011111" => rgb <= "000000";
					when "10011101010100000" => rgb <= "000000";
					when "10011101010100001" => rgb <= "000000";
					when "10011101010100010" => rgb <= "000000";
					when "10011101010100011" => rgb <= "000000";
					when "10011101010100100" => rgb <= "000000";
					when "10011101010100101" => rgb <= "000000";
					when "10011101010100110" => rgb <= "000000";
					when "10011101010100111" => rgb <= "000000";
					when "10011101010101000" => rgb <= "000000";
					when "10011101010101001" => rgb <= "000000";
					when "10011101010101010" => rgb <= "000000";
					when "10011101010101011" => rgb <= "000000";
					when "10011101010101100" => rgb <= "000000";
					when "10011101010101101" => rgb <= "000000";
					when "10011101010101110" => rgb <= "000000";
					when "10011101010101111" => rgb <= "000000";
					when "10011101010110000" => rgb <= "000000";
					when "10011101010110001" => rgb <= "000000";
					when "10011101010110010" => rgb <= "000000";
					when "10011101010110011" => rgb <= "000000";
					when "10011101010110100" => rgb <= "000000";
					when "10011101010110101" => rgb <= "000000";
					when "10011101010110110" => rgb <= "000000";
					when "10011101010110111" => rgb <= "000000";
					when "10011101010111000" => rgb <= "000000";
					when "10011101010111001" => rgb <= "000000";
					when "10011101010111010" => rgb <= "000000";
					when "10011101010111011" => rgb <= "000000";
					when "10011101010111100" => rgb <= "000000";
					when "10011101010111101" => rgb <= "000000";
					when "10011101010111110" => rgb <= "000000";
					when "10011101010111111" => rgb <= "000000";
					when "10011101011000000" => rgb <= "000000";
					when "10011101011000001" => rgb <= "000000";
					when "10011101011000010" => rgb <= "000000";
					when "10011101011000011" => rgb <= "000000";
					when "10011101011000100" => rgb <= "000000";
					when "10011101011000101" => rgb <= "000000";
					when "10011101011000110" => rgb <= "000000";
					when "10011101011000111" => rgb <= "000000";
					when "10011101011001000" => rgb <= "000000";
					when "10011101011001001" => rgb <= "000000";
					when "10011101011001010" => rgb <= "000000";
					when "10011101011001011" => rgb <= "000000";
					when "10011101011001100" => rgb <= "000000";
					when "10011101011001101" => rgb <= "000000";
					when "10011101011001110" => rgb <= "000000";
					when "10011101011001111" => rgb <= "000000";
					when "10011101011010000" => rgb <= "000000";
					when "10011101011010001" => rgb <= "000000";
					when "10011101011010010" => rgb <= "000000";
					when "10011101011010011" => rgb <= "000000";
					when "10011101011010100" => rgb <= "000000";
					when "10011101011010101" => rgb <= "000000";
					when "10011101011010110" => rgb <= "000000";
					when "10011101011010111" => rgb <= "000000";
					when "10011101011011000" => rgb <= "000000";
					when "10011101011011001" => rgb <= "000000";
					when "10011101011011010" => rgb <= "000000";
					when "10011101011011011" => rgb <= "000000";
					when "10011101011011100" => rgb <= "000000";
					when "10011101011011101" => rgb <= "000000";
					when "10011101011011110" => rgb <= "000000";
					when "10011101011011111" => rgb <= "000000";
					when "10011101011100000" => rgb <= "000000";
					when "10011101011100001" => rgb <= "000000";
					when "10011101011100010" => rgb <= "000000";
					when "10011101011100011" => rgb <= "000000";
					when "10011101011100100" => rgb <= "000000";
					when "10011101011100101" => rgb <= "000000";
					when "10011101011100110" => rgb <= "000000";
					when "10011101011100111" => rgb <= "000000";
					when "10011101011101000" => rgb <= "000000";
					when "10011101011101001" => rgb <= "000000";
					when "10011101011101010" => rgb <= "000000";
					when "10011101011101011" => rgb <= "000000";
					when "10011101011101100" => rgb <= "000000";
					when "10011101011101101" => rgb <= "000000";
					when "10011101011101110" => rgb <= "000000";
					when "10011101011101111" => rgb <= "000000";
					when "10011101011110000" => rgb <= "000000";
					when "10011101011110001" => rgb <= "000000";
					when "10011101011110010" => rgb <= "000000";
					when "10011101011110011" => rgb <= "000000";
					when "10011101011110100" => rgb <= "000000";
					when "10011101011110101" => rgb <= "000000";
					when "10011101011110110" => rgb <= "000000";
					when "10011101011110111" => rgb <= "000000";
					when "10011101011111000" => rgb <= "000000";
					when "10011101011111001" => rgb <= "000000";
					when "10011101011111010" => rgb <= "000000";
					when "10011101011111011" => rgb <= "000000";
					when "10011101011111100" => rgb <= "000000";
					when "10011101011111101" => rgb <= "000000";
					when "10011101011111110" => rgb <= "000000";
					when "10011101011111111" => rgb <= "000000";
					when "10011101100000000" => rgb <= "000000";
					when "10011101100000001" => rgb <= "000000";
					when "10011101100000010" => rgb <= "000000";
					when "10011101100000011" => rgb <= "000000";
					when "10011101100000100" => rgb <= "000000";
					when "10011101100000101" => rgb <= "000000";
					when "10011101100000110" => rgb <= "000000";
					when "10011101100000111" => rgb <= "000000";
					when "10011101100001000" => rgb <= "000000";
					when "10011101100001001" => rgb <= "000000";
					when "10011101100001010" => rgb <= "000000";
					when "10011101100001011" => rgb <= "000000";
					when "10011101100001100" => rgb <= "000000";
					when "10011101100001101" => rgb <= "000000";
					when "10011101100001110" => rgb <= "000000";
					when "10011101100001111" => rgb <= "000000";
					when "10011101100010000" => rgb <= "000000";
					when "10011101100010001" => rgb <= "000000";
					when "10011101100010010" => rgb <= "000000";
					when "10011101100010011" => rgb <= "000000";
					when "10011101100010100" => rgb <= "000000";
					when "10011101100010101" => rgb <= "000000";
					when "10011101100010110" => rgb <= "000000";
					when "10011101100010111" => rgb <= "000000";
					when "10011101100011000" => rgb <= "000000";
					when "10011101100011001" => rgb <= "000000";
					when "10011101100011010" => rgb <= "000000";
					when "10011101100011011" => rgb <= "000000";
					when "10011101100011100" => rgb <= "000000";
					when "10011101100011101" => rgb <= "000000";
					when "10011101100011110" => rgb <= "000000";
					when "10011101100011111" => rgb <= "000000";
					when "10011101100100000" => rgb <= "000000";
					when "10011101100100001" => rgb <= "000000";
					when "10011101100100010" => rgb <= "000000";
					when "10011101100100011" => rgb <= "000000";
					when "10011101100100100" => rgb <= "000000";
					when "10011101100100101" => rgb <= "000000";
					when "10011101100100110" => rgb <= "000000";
					when "10011101100100111" => rgb <= "000000";
					when "10011101100101000" => rgb <= "000000";
					when "10011101100101001" => rgb <= "000000";
					when "10011101100101010" => rgb <= "000000";
					when "10011101100101011" => rgb <= "000000";
					when "10011101100101100" => rgb <= "000000";
					when "10011101100101101" => rgb <= "000000";
					when "10011101100101110" => rgb <= "000000";
					when "10011101100101111" => rgb <= "000000";
					when "10011101100110000" => rgb <= "000000";
					when "10011101100110001" => rgb <= "000000";
					when "10011101100110010" => rgb <= "000000";
					when "10011101100110011" => rgb <= "000000";
					when "10011101100110100" => rgb <= "000000";
					when "10011101100110101" => rgb <= "000000";
					when "10011101100110110" => rgb <= "000000";
					when "10011101100110111" => rgb <= "000000";
					when "10011101100111000" => rgb <= "000000";
					when "10011101100111001" => rgb <= "000000";
					when "10011101100111010" => rgb <= "000000";
					when "10011101100111011" => rgb <= "000000";
					when "10011101100111100" => rgb <= "000000";
					when "10011101100111101" => rgb <= "000000";
					when "10011101100111110" => rgb <= "000000";
					when "10011101100111111" => rgb <= "000000";
					when "10011110000000000" => rgb <= "000000";
					when "10011110000000001" => rgb <= "000000";
					when "10011110000000010" => rgb <= "000000";
					when "10011110000000011" => rgb <= "000000";
					when "10011110000000100" => rgb <= "000000";
					when "10011110000000101" => rgb <= "000000";
					when "10011110000000110" => rgb <= "000000";
					when "10011110000000111" => rgb <= "000000";
					when "10011110000001000" => rgb <= "000000";
					when "10011110000001001" => rgb <= "000000";
					when "10011110000001010" => rgb <= "000000";
					when "10011110000001011" => rgb <= "000000";
					when "10011110000001100" => rgb <= "000000";
					when "10011110000001101" => rgb <= "000000";
					when "10011110000001110" => rgb <= "000000";
					when "10011110000001111" => rgb <= "000000";
					when "10011110000010000" => rgb <= "000000";
					when "10011110000010001" => rgb <= "000000";
					when "10011110000010010" => rgb <= "000000";
					when "10011110000010011" => rgb <= "000000";
					when "10011110000010100" => rgb <= "000000";
					when "10011110000010101" => rgb <= "000000";
					when "10011110000010110" => rgb <= "000000";
					when "10011110000010111" => rgb <= "000000";
					when "10011110000011000" => rgb <= "000000";
					when "10011110000011001" => rgb <= "000000";
					when "10011110000011010" => rgb <= "000000";
					when "10011110000011011" => rgb <= "000000";
					when "10011110000011100" => rgb <= "000000";
					when "10011110000011101" => rgb <= "000000";
					when "10011110000011110" => rgb <= "000000";
					when "10011110000011111" => rgb <= "000000";
					when "10011110000100000" => rgb <= "000000";
					when "10011110000100001" => rgb <= "000000";
					when "10011110000100010" => rgb <= "000000";
					when "10011110000100011" => rgb <= "000000";
					when "10011110000100100" => rgb <= "000000";
					when "10011110000100101" => rgb <= "000000";
					when "10011110000100110" => rgb <= "000000";
					when "10011110000100111" => rgb <= "000000";
					when "10011110000101000" => rgb <= "000000";
					when "10011110000101001" => rgb <= "000000";
					when "10011110000101010" => rgb <= "000000";
					when "10011110000101011" => rgb <= "000000";
					when "10011110000101100" => rgb <= "000000";
					when "10011110000101101" => rgb <= "000000";
					when "10011110000101110" => rgb <= "000000";
					when "10011110000101111" => rgb <= "000000";
					when "10011110000110000" => rgb <= "000000";
					when "10011110000110001" => rgb <= "000000";
					when "10011110000110010" => rgb <= "000000";
					when "10011110000110011" => rgb <= "000000";
					when "10011110000110100" => rgb <= "000000";
					when "10011110000110101" => rgb <= "000000";
					when "10011110000110110" => rgb <= "000000";
					when "10011110000110111" => rgb <= "000000";
					when "10011110000111000" => rgb <= "000000";
					when "10011110000111001" => rgb <= "000000";
					when "10011110000111010" => rgb <= "000000";
					when "10011110000111011" => rgb <= "000000";
					when "10011110000111100" => rgb <= "000000";
					when "10011110000111101" => rgb <= "000000";
					when "10011110000111110" => rgb <= "000000";
					when "10011110000111111" => rgb <= "000000";
					when "10011110001000000" => rgb <= "000000";
					when "10011110001000001" => rgb <= "000000";
					when "10011110001000010" => rgb <= "000000";
					when "10011110001000011" => rgb <= "000000";
					when "10011110001000100" => rgb <= "000000";
					when "10011110001000101" => rgb <= "000000";
					when "10011110001000110" => rgb <= "000000";
					when "10011110001000111" => rgb <= "000000";
					when "10011110001001000" => rgb <= "000000";
					when "10011110001001001" => rgb <= "000000";
					when "10011110001001010" => rgb <= "000000";
					when "10011110001001011" => rgb <= "000000";
					when "10011110001001100" => rgb <= "000000";
					when "10011110001001101" => rgb <= "000000";
					when "10011110001001110" => rgb <= "000000";
					when "10011110001001111" => rgb <= "000000";
					when "10011110001010000" => rgb <= "000000";
					when "10011110001010001" => rgb <= "000000";
					when "10011110001010010" => rgb <= "000000";
					when "10011110001010011" => rgb <= "000000";
					when "10011110001010100" => rgb <= "000000";
					when "10011110001010101" => rgb <= "000000";
					when "10011110001010110" => rgb <= "000000";
					when "10011110001010111" => rgb <= "000000";
					when "10011110001011000" => rgb <= "000000";
					when "10011110001011001" => rgb <= "000000";
					when "10011110001011010" => rgb <= "000000";
					when "10011110001011011" => rgb <= "000000";
					when "10011110001011100" => rgb <= "000000";
					when "10011110001011101" => rgb <= "000000";
					when "10011110001011110" => rgb <= "000000";
					when "10011110001011111" => rgb <= "000000";
					when "10011110001100000" => rgb <= "000000";
					when "10011110001100001" => rgb <= "000000";
					when "10011110001100010" => rgb <= "000000";
					when "10011110001100011" => rgb <= "000000";
					when "10011110001100100" => rgb <= "000000";
					when "10011110001100101" => rgb <= "000000";
					when "10011110001100110" => rgb <= "000000";
					when "10011110001100111" => rgb <= "000000";
					when "10011110001101000" => rgb <= "000000";
					when "10011110001101001" => rgb <= "000000";
					when "10011110001101010" => rgb <= "000000";
					when "10011110001101011" => rgb <= "000000";
					when "10011110001101100" => rgb <= "000000";
					when "10011110001101101" => rgb <= "000000";
					when "10011110001101110" => rgb <= "000000";
					when "10011110001101111" => rgb <= "000000";
					when "10011110001110000" => rgb <= "000000";
					when "10011110001110001" => rgb <= "000000";
					when "10011110001110010" => rgb <= "000000";
					when "10011110001110011" => rgb <= "000000";
					when "10011110001110100" => rgb <= "000000";
					when "10011110001110101" => rgb <= "000000";
					when "10011110001110110" => rgb <= "000000";
					when "10011110001110111" => rgb <= "000000";
					when "10011110001111000" => rgb <= "000000";
					when "10011110001111001" => rgb <= "000000";
					when "10011110001111010" => rgb <= "000000";
					when "10011110001111011" => rgb <= "000000";
					when "10011110001111100" => rgb <= "000000";
					when "10011110001111101" => rgb <= "000000";
					when "10011110001111110" => rgb <= "000000";
					when "10011110001111111" => rgb <= "000000";
					when "10011110010000000" => rgb <= "000000";
					when "10011110010000001" => rgb <= "000000";
					when "10011110010000010" => rgb <= "000000";
					when "10011110010000011" => rgb <= "000000";
					when "10011110010000100" => rgb <= "000000";
					when "10011110010000101" => rgb <= "000000";
					when "10011110010000110" => rgb <= "000000";
					when "10011110010000111" => rgb <= "000000";
					when "10011110010001000" => rgb <= "000000";
					when "10011110010001001" => rgb <= "000000";
					when "10011110010001010" => rgb <= "000000";
					when "10011110010001011" => rgb <= "000000";
					when "10011110010001100" => rgb <= "000000";
					when "10011110010001101" => rgb <= "000000";
					when "10011110010001110" => rgb <= "000000";
					when "10011110010001111" => rgb <= "000000";
					when "10011110010010000" => rgb <= "000000";
					when "10011110010010001" => rgb <= "000000";
					when "10011110010010010" => rgb <= "000000";
					when "10011110010010011" => rgb <= "000000";
					when "10011110010010100" => rgb <= "000000";
					when "10011110010010101" => rgb <= "000000";
					when "10011110010010110" => rgb <= "000000";
					when "10011110010010111" => rgb <= "000000";
					when "10011110010011000" => rgb <= "000000";
					when "10011110010011001" => rgb <= "000000";
					when "10011110010011010" => rgb <= "000000";
					when "10011110010011011" => rgb <= "000000";
					when "10011110010011100" => rgb <= "000000";
					when "10011110010011101" => rgb <= "000000";
					when "10011110010011110" => rgb <= "000000";
					when "10011110010011111" => rgb <= "000000";
					when "10011110010100000" => rgb <= "000000";
					when "10011110010100001" => rgb <= "000000";
					when "10011110010100010" => rgb <= "000000";
					when "10011110010100011" => rgb <= "000000";
					when "10011110010100100" => rgb <= "000000";
					when "10011110010100101" => rgb <= "000000";
					when "10011110010100110" => rgb <= "000000";
					when "10011110010100111" => rgb <= "000000";
					when "10011110010101000" => rgb <= "000000";
					when "10011110010101001" => rgb <= "000000";
					when "10011110010101010" => rgb <= "000000";
					when "10011110010101011" => rgb <= "000000";
					when "10011110010101100" => rgb <= "000000";
					when "10011110010101101" => rgb <= "000000";
					when "10011110010101110" => rgb <= "000000";
					when "10011110010101111" => rgb <= "000000";
					when "10011110010110000" => rgb <= "000000";
					when "10011110010110001" => rgb <= "000000";
					when "10011110010110010" => rgb <= "000000";
					when "10011110010110011" => rgb <= "000000";
					when "10011110010110100" => rgb <= "000000";
					when "10011110010110101" => rgb <= "000000";
					when "10011110010110110" => rgb <= "000000";
					when "10011110010110111" => rgb <= "000000";
					when "10011110010111000" => rgb <= "000000";
					when "10011110010111001" => rgb <= "000000";
					when "10011110010111010" => rgb <= "000000";
					when "10011110010111011" => rgb <= "000000";
					when "10011110010111100" => rgb <= "000000";
					when "10011110010111101" => rgb <= "000000";
					when "10011110010111110" => rgb <= "000000";
					when "10011110010111111" => rgb <= "000000";
					when "10011110011000000" => rgb <= "000000";
					when "10011110011000001" => rgb <= "000000";
					when "10011110011000010" => rgb <= "000000";
					when "10011110011000011" => rgb <= "000000";
					when "10011110011000100" => rgb <= "000000";
					when "10011110011000101" => rgb <= "000000";
					when "10011110011000110" => rgb <= "000000";
					when "10011110011000111" => rgb <= "000000";
					when "10011110011001000" => rgb <= "000000";
					when "10011110011001001" => rgb <= "000000";
					when "10011110011001010" => rgb <= "000000";
					when "10011110011001011" => rgb <= "000000";
					when "10011110011001100" => rgb <= "000000";
					when "10011110011001101" => rgb <= "000000";
					when "10011110011001110" => rgb <= "000000";
					when "10011110011001111" => rgb <= "000000";
					when "10011110011010000" => rgb <= "000000";
					when "10011110011010001" => rgb <= "000000";
					when "10011110011010010" => rgb <= "000000";
					when "10011110011010011" => rgb <= "000000";
					when "10011110011010100" => rgb <= "000000";
					when "10011110011010101" => rgb <= "000000";
					when "10011110011010110" => rgb <= "000000";
					when "10011110011010111" => rgb <= "000000";
					when "10011110011011000" => rgb <= "000000";
					when "10011110011011001" => rgb <= "000000";
					when "10011110011011010" => rgb <= "000000";
					when "10011110011011011" => rgb <= "000000";
					when "10011110011011100" => rgb <= "000000";
					when "10011110011011101" => rgb <= "000000";
					when "10011110011011110" => rgb <= "000000";
					when "10011110011011111" => rgb <= "000000";
					when "10011110011100000" => rgb <= "000000";
					when "10011110011100001" => rgb <= "000000";
					when "10011110011100010" => rgb <= "000000";
					when "10011110011100011" => rgb <= "000000";
					when "10011110011100100" => rgb <= "000000";
					when "10011110011100101" => rgb <= "000000";
					when "10011110011100110" => rgb <= "000000";
					when "10011110011100111" => rgb <= "000000";
					when "10011110011101000" => rgb <= "000000";
					when "10011110011101001" => rgb <= "000000";
					when "10011110011101010" => rgb <= "000000";
					when "10011110011101011" => rgb <= "000000";
					when "10011110011101100" => rgb <= "000000";
					when "10011110011101101" => rgb <= "000000";
					when "10011110011101110" => rgb <= "000000";
					when "10011110011101111" => rgb <= "000000";
					when "10011110011110000" => rgb <= "000000";
					when "10011110011110001" => rgb <= "000000";
					when "10011110011110010" => rgb <= "000000";
					when "10011110011110011" => rgb <= "000000";
					when "10011110011110100" => rgb <= "000000";
					when "10011110011110101" => rgb <= "000000";
					when "10011110011110110" => rgb <= "000000";
					when "10011110011110111" => rgb <= "000000";
					when "10011110011111000" => rgb <= "000000";
					when "10011110011111001" => rgb <= "000000";
					when "10011110011111010" => rgb <= "000000";
					when "10011110011111011" => rgb <= "000000";
					when "10011110011111100" => rgb <= "000000";
					when "10011110011111101" => rgb <= "000000";
					when "10011110011111110" => rgb <= "000000";
					when "10011110011111111" => rgb <= "000000";
					when "10011110100000000" => rgb <= "000000";
					when "10011110100000001" => rgb <= "000000";
					when "10011110100000010" => rgb <= "000000";
					when "10011110100000011" => rgb <= "000000";
					when "10011110100000100" => rgb <= "000000";
					when "10011110100000101" => rgb <= "000000";
					when "10011110100000110" => rgb <= "000000";
					when "10011110100000111" => rgb <= "000000";
					when "10011110100001000" => rgb <= "000000";
					when "10011110100001001" => rgb <= "000000";
					when "10011110100001010" => rgb <= "000000";
					when "10011110100001011" => rgb <= "000000";
					when "10011110100001100" => rgb <= "000000";
					when "10011110100001101" => rgb <= "000000";
					when "10011110100001110" => rgb <= "000000";
					when "10011110100001111" => rgb <= "000000";
					when "10011110100010000" => rgb <= "000000";
					when "10011110100010001" => rgb <= "000000";
					when "10011110100010010" => rgb <= "000000";
					when "10011110100010011" => rgb <= "000000";
					when "10011110100010100" => rgb <= "000000";
					when "10011110100010101" => rgb <= "000000";
					when "10011110100010110" => rgb <= "000000";
					when "10011110100010111" => rgb <= "000000";
					when "10011110100011000" => rgb <= "000000";
					when "10011110100011001" => rgb <= "000000";
					when "10011110100011010" => rgb <= "000000";
					when "10011110100011011" => rgb <= "000000";
					when "10011110100011100" => rgb <= "000000";
					when "10011110100011101" => rgb <= "000000";
					when "10011110100011110" => rgb <= "000000";
					when "10011110100011111" => rgb <= "000000";
					when "10011110100100000" => rgb <= "000000";
					when "10011110100100001" => rgb <= "000000";
					when "10011110100100010" => rgb <= "000000";
					when "10011110100100011" => rgb <= "000000";
					when "10011110100100100" => rgb <= "000000";
					when "10011110100100101" => rgb <= "000000";
					when "10011110100100110" => rgb <= "000000";
					when "10011110100100111" => rgb <= "000000";
					when "10011110100101000" => rgb <= "000000";
					when "10011110100101001" => rgb <= "000000";
					when "10011110100101010" => rgb <= "000000";
					when "10011110100101011" => rgb <= "000000";
					when "10011110100101100" => rgb <= "000000";
					when "10011110100101101" => rgb <= "000000";
					when "10011110100101110" => rgb <= "000000";
					when "10011110100101111" => rgb <= "000000";
					when "10011110100110000" => rgb <= "000000";
					when "10011110100110001" => rgb <= "000000";
					when "10011110100110010" => rgb <= "000000";
					when "10011110100110011" => rgb <= "000000";
					when "10011110100110100" => rgb <= "000000";
					when "10011110100110101" => rgb <= "000000";
					when "10011110100110110" => rgb <= "000000";
					when "10011110100110111" => rgb <= "000000";
					when "10011110100111000" => rgb <= "000000";
					when "10011110100111001" => rgb <= "000000";
					when "10011110100111010" => rgb <= "000000";
					when "10011110100111011" => rgb <= "000000";
					when "10011110100111100" => rgb <= "000000";
					when "10011110100111101" => rgb <= "000000";
					when "10011110100111110" => rgb <= "000000";
					when "10011110100111111" => rgb <= "000000";
					when "10011111000000000" => rgb <= "000000";
					when "10011111000000001" => rgb <= "000000";
					when "10011111000000010" => rgb <= "000000";
					when "10011111000000011" => rgb <= "000000";
					when "10011111000000100" => rgb <= "000000";
					when "10011111000000101" => rgb <= "000000";
					when "10011111000000110" => rgb <= "000000";
					when "10011111000000111" => rgb <= "000000";
					when "10011111000001000" => rgb <= "000000";
					when "10011111000001001" => rgb <= "000000";
					when "10011111000001010" => rgb <= "000000";
					when "10011111000001011" => rgb <= "000000";
					when "10011111000001100" => rgb <= "000000";
					when "10011111000001101" => rgb <= "000000";
					when "10011111000001110" => rgb <= "000000";
					when "10011111000001111" => rgb <= "000000";
					when "10011111000010000" => rgb <= "000000";
					when "10011111000010001" => rgb <= "000000";
					when "10011111000010010" => rgb <= "000000";
					when "10011111000010011" => rgb <= "000000";
					when "10011111000010100" => rgb <= "000000";
					when "10011111000010101" => rgb <= "000000";
					when "10011111000010110" => rgb <= "000000";
					when "10011111000010111" => rgb <= "000000";
					when "10011111000011000" => rgb <= "000000";
					when "10011111000011001" => rgb <= "000000";
					when "10011111000011010" => rgb <= "000000";
					when "10011111000011011" => rgb <= "000000";
					when "10011111000011100" => rgb <= "000000";
					when "10011111000011101" => rgb <= "000000";
					when "10011111000011110" => rgb <= "000000";
					when "10011111000011111" => rgb <= "000000";
					when "10011111000100000" => rgb <= "000000";
					when "10011111000100001" => rgb <= "000000";
					when "10011111000100010" => rgb <= "000000";
					when "10011111000100011" => rgb <= "000000";
					when "10011111000100100" => rgb <= "000000";
					when "10011111000100101" => rgb <= "000000";
					when "10011111000100110" => rgb <= "000000";
					when "10011111000100111" => rgb <= "000000";
					when "10011111000101000" => rgb <= "000000";
					when "10011111000101001" => rgb <= "000000";
					when "10011111000101010" => rgb <= "000000";
					when "10011111000101011" => rgb <= "000000";
					when "10011111000101100" => rgb <= "000000";
					when "10011111000101101" => rgb <= "000000";
					when "10011111000101110" => rgb <= "000000";
					when "10011111000101111" => rgb <= "000000";
					when "10011111000110000" => rgb <= "000000";
					when "10011111000110001" => rgb <= "000000";
					when "10011111000110010" => rgb <= "000000";
					when "10011111000110011" => rgb <= "000000";
					when "10011111000110100" => rgb <= "000000";
					when "10011111000110101" => rgb <= "000000";
					when "10011111000110110" => rgb <= "000000";
					when "10011111000110111" => rgb <= "000000";
					when "10011111000111000" => rgb <= "000000";
					when "10011111000111001" => rgb <= "000000";
					when "10011111000111010" => rgb <= "000000";
					when "10011111000111011" => rgb <= "000000";
					when "10011111000111100" => rgb <= "000000";
					when "10011111000111101" => rgb <= "000000";
					when "10011111000111110" => rgb <= "000000";
					when "10011111000111111" => rgb <= "000000";
					when "10011111001000000" => rgb <= "000000";
					when "10011111001000001" => rgb <= "000000";
					when "10011111001000010" => rgb <= "000000";
					when "10011111001000011" => rgb <= "000000";
					when "10011111001000100" => rgb <= "000000";
					when "10011111001000101" => rgb <= "000000";
					when "10011111001000110" => rgb <= "000000";
					when "10011111001000111" => rgb <= "000000";
					when "10011111001001000" => rgb <= "000000";
					when "10011111001001001" => rgb <= "000000";
					when "10011111001001010" => rgb <= "000000";
					when "10011111001001011" => rgb <= "000000";
					when "10011111001001100" => rgb <= "000000";
					when "10011111001001101" => rgb <= "000000";
					when "10011111001001110" => rgb <= "000000";
					when "10011111001001111" => rgb <= "000000";
					when "10011111001010000" => rgb <= "000000";
					when "10011111001010001" => rgb <= "000000";
					when "10011111001010010" => rgb <= "000000";
					when "10011111001010011" => rgb <= "000000";
					when "10011111001010100" => rgb <= "000000";
					when "10011111001010101" => rgb <= "000000";
					when "10011111001010110" => rgb <= "000000";
					when "10011111001010111" => rgb <= "000000";
					when "10011111001011000" => rgb <= "000000";
					when "10011111001011001" => rgb <= "000000";
					when "10011111001011010" => rgb <= "000000";
					when "10011111001011011" => rgb <= "000000";
					when "10011111001011100" => rgb <= "000000";
					when "10011111001011101" => rgb <= "000000";
					when "10011111001011110" => rgb <= "000000";
					when "10011111001011111" => rgb <= "000000";
					when "10011111001100000" => rgb <= "000000";
					when "10011111001100001" => rgb <= "000000";
					when "10011111001100010" => rgb <= "000000";
					when "10011111001100011" => rgb <= "000000";
					when "10011111001100100" => rgb <= "000000";
					when "10011111001100101" => rgb <= "000000";
					when "10011111001100110" => rgb <= "000000";
					when "10011111001100111" => rgb <= "000000";
					when "10011111001101000" => rgb <= "000000";
					when "10011111001101001" => rgb <= "000000";
					when "10011111001101010" => rgb <= "000000";
					when "10011111001101011" => rgb <= "000000";
					when "10011111001101100" => rgb <= "000000";
					when "10011111001101101" => rgb <= "000000";
					when "10011111001101110" => rgb <= "000000";
					when "10011111001101111" => rgb <= "000000";
					when "10011111001110000" => rgb <= "000000";
					when "10011111001110001" => rgb <= "000000";
					when "10011111001110010" => rgb <= "000000";
					when "10011111001110011" => rgb <= "000000";
					when "10011111001110100" => rgb <= "000000";
					when "10011111001110101" => rgb <= "000000";
					when "10011111001110110" => rgb <= "000000";
					when "10011111001110111" => rgb <= "000000";
					when "10011111001111000" => rgb <= "000000";
					when "10011111001111001" => rgb <= "000000";
					when "10011111001111010" => rgb <= "000000";
					when "10011111001111011" => rgb <= "000000";
					when "10011111001111100" => rgb <= "000000";
					when "10011111001111101" => rgb <= "000000";
					when "10011111001111110" => rgb <= "000000";
					when "10011111001111111" => rgb <= "000000";
					when "10011111010000000" => rgb <= "000000";
					when "10011111010000001" => rgb <= "000000";
					when "10011111010000010" => rgb <= "000000";
					when "10011111010000011" => rgb <= "000000";
					when "10011111010000100" => rgb <= "000000";
					when "10011111010000101" => rgb <= "000000";
					when "10011111010000110" => rgb <= "000000";
					when "10011111010000111" => rgb <= "000000";
					when "10011111010001000" => rgb <= "000000";
					when "10011111010001001" => rgb <= "000000";
					when "10011111010001010" => rgb <= "000000";
					when "10011111010001011" => rgb <= "000000";
					when "10011111010001100" => rgb <= "000000";
					when "10011111010001101" => rgb <= "000000";
					when "10011111010001110" => rgb <= "000000";
					when "10011111010001111" => rgb <= "000000";
					when "10011111010010000" => rgb <= "000000";
					when "10011111010010001" => rgb <= "000000";
					when "10011111010010010" => rgb <= "000000";
					when "10011111010010011" => rgb <= "000000";
					when "10011111010010100" => rgb <= "000000";
					when "10011111010010101" => rgb <= "000000";
					when "10011111010010110" => rgb <= "000000";
					when "10011111010010111" => rgb <= "000000";
					when "10011111010011000" => rgb <= "000000";
					when "10011111010011001" => rgb <= "000000";
					when "10011111010011010" => rgb <= "000000";
					when "10011111010011011" => rgb <= "000000";
					when "10011111010011100" => rgb <= "000000";
					when "10011111010011101" => rgb <= "000000";
					when "10011111010011110" => rgb <= "000000";
					when "10011111010011111" => rgb <= "000000";
					when "10011111010100000" => rgb <= "000000";
					when "10011111010100001" => rgb <= "000000";
					when "10011111010100010" => rgb <= "000000";
					when "10011111010100011" => rgb <= "000000";
					when "10011111010100100" => rgb <= "000000";
					when "10011111010100101" => rgb <= "000000";
					when "10011111010100110" => rgb <= "000000";
					when "10011111010100111" => rgb <= "000000";
					when "10011111010101000" => rgb <= "000000";
					when "10011111010101001" => rgb <= "000000";
					when "10011111010101010" => rgb <= "000000";
					when "10011111010101011" => rgb <= "000000";
					when "10011111010101100" => rgb <= "000000";
					when "10011111010101101" => rgb <= "000000";
					when "10011111010101110" => rgb <= "000000";
					when "10011111010101111" => rgb <= "000000";
					when "10011111010110000" => rgb <= "000000";
					when "10011111010110001" => rgb <= "000000";
					when "10011111010110010" => rgb <= "000000";
					when "10011111010110011" => rgb <= "000000";
					when "10011111010110100" => rgb <= "000000";
					when "10011111010110101" => rgb <= "000000";
					when "10011111010110110" => rgb <= "000000";
					when "10011111010110111" => rgb <= "000000";
					when "10011111010111000" => rgb <= "000000";
					when "10011111010111001" => rgb <= "000000";
					when "10011111010111010" => rgb <= "000000";
					when "10011111010111011" => rgb <= "000000";
					when "10011111010111100" => rgb <= "000000";
					when "10011111010111101" => rgb <= "000000";
					when "10011111010111110" => rgb <= "000000";
					when "10011111010111111" => rgb <= "000000";
					when "10011111011000000" => rgb <= "000000";
					when "10011111011000001" => rgb <= "000000";
					when "10011111011000010" => rgb <= "000000";
					when "10011111011000011" => rgb <= "000000";
					when "10011111011000100" => rgb <= "000000";
					when "10011111011000101" => rgb <= "000000";
					when "10011111011000110" => rgb <= "000000";
					when "10011111011000111" => rgb <= "000000";
					when "10011111011001000" => rgb <= "000000";
					when "10011111011001001" => rgb <= "000000";
					when "10011111011001010" => rgb <= "000000";
					when "10011111011001011" => rgb <= "000000";
					when "10011111011001100" => rgb <= "000000";
					when "10011111011001101" => rgb <= "000000";
					when "10011111011001110" => rgb <= "000000";
					when "10011111011001111" => rgb <= "000000";
					when "10011111011010000" => rgb <= "000000";
					when "10011111011010001" => rgb <= "000000";
					when "10011111011010010" => rgb <= "000000";
					when "10011111011010011" => rgb <= "000000";
					when "10011111011010100" => rgb <= "000000";
					when "10011111011010101" => rgb <= "000000";
					when "10011111011010110" => rgb <= "000000";
					when "10011111011010111" => rgb <= "000000";
					when "10011111011011000" => rgb <= "000000";
					when "10011111011011001" => rgb <= "000000";
					when "10011111011011010" => rgb <= "000000";
					when "10011111011011011" => rgb <= "000000";
					when "10011111011011100" => rgb <= "000000";
					when "10011111011011101" => rgb <= "000000";
					when "10011111011011110" => rgb <= "000000";
					when "10011111011011111" => rgb <= "000000";
					when "10011111011100000" => rgb <= "000000";
					when "10011111011100001" => rgb <= "000000";
					when "10011111011100010" => rgb <= "000000";
					when "10011111011100011" => rgb <= "000000";
					when "10011111011100100" => rgb <= "000000";
					when "10011111011100101" => rgb <= "000000";
					when "10011111011100110" => rgb <= "000000";
					when "10011111011100111" => rgb <= "000000";
					when "10011111011101000" => rgb <= "000000";
					when "10011111011101001" => rgb <= "000000";
					when "10011111011101010" => rgb <= "000000";
					when "10011111011101011" => rgb <= "000000";
					when "10011111011101100" => rgb <= "000000";
					when "10011111011101101" => rgb <= "000000";
					when "10011111011101110" => rgb <= "000000";
					when "10011111011101111" => rgb <= "000000";
					when "10011111011110000" => rgb <= "000000";
					when "10011111011110001" => rgb <= "000000";
					when "10011111011110010" => rgb <= "000000";
					when "10011111011110011" => rgb <= "000000";
					when "10011111011110100" => rgb <= "000000";
					when "10011111011110101" => rgb <= "000000";
					when "10011111011110110" => rgb <= "000000";
					when "10011111011110111" => rgb <= "000000";
					when "10011111011111000" => rgb <= "000000";
					when "10011111011111001" => rgb <= "000000";
					when "10011111011111010" => rgb <= "000000";
					when "10011111011111011" => rgb <= "000000";
					when "10011111011111100" => rgb <= "000000";
					when "10011111011111101" => rgb <= "000000";
					when "10011111011111110" => rgb <= "000000";
					when "10011111011111111" => rgb <= "000000";
					when "10011111100000000" => rgb <= "000000";
					when "10011111100000001" => rgb <= "000000";
					when "10011111100000010" => rgb <= "000000";
					when "10011111100000011" => rgb <= "000000";
					when "10011111100000100" => rgb <= "000000";
					when "10011111100000101" => rgb <= "000000";
					when "10011111100000110" => rgb <= "000000";
					when "10011111100000111" => rgb <= "000000";
					when "10011111100001000" => rgb <= "000000";
					when "10011111100001001" => rgb <= "000000";
					when "10011111100001010" => rgb <= "000000";
					when "10011111100001011" => rgb <= "000000";
					when "10011111100001100" => rgb <= "000000";
					when "10011111100001101" => rgb <= "000000";
					when "10011111100001110" => rgb <= "000000";
					when "10011111100001111" => rgb <= "000000";
					when "10011111100010000" => rgb <= "000000";
					when "10011111100010001" => rgb <= "000000";
					when "10011111100010010" => rgb <= "000000";
					when "10011111100010011" => rgb <= "000000";
					when "10011111100010100" => rgb <= "000000";
					when "10011111100010101" => rgb <= "000000";
					when "10011111100010110" => rgb <= "000000";
					when "10011111100010111" => rgb <= "000000";
					when "10011111100011000" => rgb <= "000000";
					when "10011111100011001" => rgb <= "000000";
					when "10011111100011010" => rgb <= "000000";
					when "10011111100011011" => rgb <= "000000";
					when "10011111100011100" => rgb <= "000000";
					when "10011111100011101" => rgb <= "000000";
					when "10011111100011110" => rgb <= "000000";
					when "10011111100011111" => rgb <= "000000";
					when "10011111100100000" => rgb <= "000000";
					when "10011111100100001" => rgb <= "000000";
					when "10011111100100010" => rgb <= "000000";
					when "10011111100100011" => rgb <= "000000";
					when "10011111100100100" => rgb <= "000000";
					when "10011111100100101" => rgb <= "000000";
					when "10011111100100110" => rgb <= "000000";
					when "10011111100100111" => rgb <= "000000";
					when "10011111100101000" => rgb <= "000000";
					when "10011111100101001" => rgb <= "000000";
					when "10011111100101010" => rgb <= "000000";
					when "10011111100101011" => rgb <= "000000";
					when "10011111100101100" => rgb <= "000000";
					when "10011111100101101" => rgb <= "000000";
					when "10011111100101110" => rgb <= "000000";
					when "10011111100101111" => rgb <= "000000";
					when "10011111100110000" => rgb <= "000000";
					when "10011111100110001" => rgb <= "000000";
					when "10011111100110010" => rgb <= "000000";
					when "10011111100110011" => rgb <= "000000";
					when "10011111100110100" => rgb <= "000000";
					when "10011111100110101" => rgb <= "000000";
					when "10011111100110110" => rgb <= "000000";
					when "10011111100110111" => rgb <= "000000";
					when "10011111100111000" => rgb <= "000000";
					when "10011111100111001" => rgb <= "000000";
					when "10011111100111010" => rgb <= "000000";
					when "10011111100111011" => rgb <= "000000";
					when "10011111100111100" => rgb <= "000000";
					when "10011111100111101" => rgb <= "000000";
					when "10011111100111110" => rgb <= "000000";
					when "10011111100111111" => rgb <= "000000";
					when "10100000000000000" => rgb <= "000000";
					when "10100000000000001" => rgb <= "000000";
					when "10100000000000010" => rgb <= "000000";
					when "10100000000000011" => rgb <= "000000";
					when "10100000000000100" => rgb <= "000000";
					when "10100000000000101" => rgb <= "000000";
					when "10100000000000110" => rgb <= "000000";
					when "10100000000000111" => rgb <= "000000";
					when "10100000000001000" => rgb <= "000000";
					when "10100000000001001" => rgb <= "000000";
					when "10100000000001010" => rgb <= "000000";
					when "10100000000001011" => rgb <= "000000";
					when "10100000000001100" => rgb <= "000000";
					when "10100000000001101" => rgb <= "000000";
					when "10100000000001110" => rgb <= "000000";
					when "10100000000001111" => rgb <= "000000";
					when "10100000000010000" => rgb <= "000000";
					when "10100000000010001" => rgb <= "000000";
					when "10100000000010010" => rgb <= "000000";
					when "10100000000010011" => rgb <= "000000";
					when "10100000000010100" => rgb <= "000000";
					when "10100000000010101" => rgb <= "000000";
					when "10100000000010110" => rgb <= "000000";
					when "10100000000010111" => rgb <= "000000";
					when "10100000000011000" => rgb <= "000000";
					when "10100000000011001" => rgb <= "000000";
					when "10100000000011010" => rgb <= "000000";
					when "10100000000011011" => rgb <= "000000";
					when "10100000000011100" => rgb <= "000000";
					when "10100000000011101" => rgb <= "000000";
					when "10100000000011110" => rgb <= "000000";
					when "10100000000011111" => rgb <= "000000";
					when "10100000000100000" => rgb <= "000000";
					when "10100000000100001" => rgb <= "000000";
					when "10100000000100010" => rgb <= "000000";
					when "10100000000100011" => rgb <= "000000";
					when "10100000000100100" => rgb <= "000000";
					when "10100000000100101" => rgb <= "000000";
					when "10100000000100110" => rgb <= "000000";
					when "10100000000100111" => rgb <= "000000";
					when "10100000000101000" => rgb <= "000000";
					when "10100000000101001" => rgb <= "000000";
					when "10100000000101010" => rgb <= "000000";
					when "10100000000101011" => rgb <= "000000";
					when "10100000000101100" => rgb <= "000000";
					when "10100000000101101" => rgb <= "000000";
					when "10100000000101110" => rgb <= "000000";
					when "10100000000101111" => rgb <= "000000";
					when "10100000000110000" => rgb <= "000000";
					when "10100000000110001" => rgb <= "000000";
					when "10100000000110010" => rgb <= "000000";
					when "10100000000110011" => rgb <= "000000";
					when "10100000000110100" => rgb <= "000000";
					when "10100000000110101" => rgb <= "000000";
					when "10100000000110110" => rgb <= "000000";
					when "10100000000110111" => rgb <= "000000";
					when "10100000000111000" => rgb <= "000000";
					when "10100000000111001" => rgb <= "000000";
					when "10100000000111010" => rgb <= "000000";
					when "10100000000111011" => rgb <= "000000";
					when "10100000000111100" => rgb <= "000000";
					when "10100000000111101" => rgb <= "000000";
					when "10100000000111110" => rgb <= "000000";
					when "10100000000111111" => rgb <= "000000";
					when "10100000001000000" => rgb <= "000000";
					when "10100000001000001" => rgb <= "000000";
					when "10100000001000010" => rgb <= "000000";
					when "10100000001000011" => rgb <= "000000";
					when "10100000001000100" => rgb <= "000000";
					when "10100000001000101" => rgb <= "000000";
					when "10100000001000110" => rgb <= "000000";
					when "10100000001000111" => rgb <= "000000";
					when "10100000001001000" => rgb <= "000000";
					when "10100000001001001" => rgb <= "000000";
					when "10100000001001010" => rgb <= "000000";
					when "10100000001001011" => rgb <= "000000";
					when "10100000001001100" => rgb <= "000000";
					when "10100000001001101" => rgb <= "000000";
					when "10100000001001110" => rgb <= "000000";
					when "10100000001001111" => rgb <= "000000";
					when "10100000001010000" => rgb <= "000000";
					when "10100000001010001" => rgb <= "000000";
					when "10100000001010010" => rgb <= "000000";
					when "10100000001010011" => rgb <= "000000";
					when "10100000001010100" => rgb <= "000000";
					when "10100000001010101" => rgb <= "000000";
					when "10100000001010110" => rgb <= "000000";
					when "10100000001010111" => rgb <= "000000";
					when "10100000001011000" => rgb <= "000000";
					when "10100000001011001" => rgb <= "000000";
					when "10100000001011010" => rgb <= "000000";
					when "10100000001011011" => rgb <= "000000";
					when "10100000001011100" => rgb <= "000000";
					when "10100000001011101" => rgb <= "000000";
					when "10100000001011110" => rgb <= "000000";
					when "10100000001011111" => rgb <= "000000";
					when "10100000001100000" => rgb <= "000000";
					when "10100000001100001" => rgb <= "000000";
					when "10100000001100010" => rgb <= "000000";
					when "10100000001100011" => rgb <= "000000";
					when "10100000001100100" => rgb <= "000000";
					when "10100000001100101" => rgb <= "000000";
					when "10100000001100110" => rgb <= "000000";
					when "10100000001100111" => rgb <= "000000";
					when "10100000001101000" => rgb <= "000000";
					when "10100000001101001" => rgb <= "000000";
					when "10100000001101010" => rgb <= "000000";
					when "10100000001101011" => rgb <= "000000";
					when "10100000001101100" => rgb <= "000000";
					when "10100000001101101" => rgb <= "000000";
					when "10100000001101110" => rgb <= "000000";
					when "10100000001101111" => rgb <= "000000";
					when "10100000001110000" => rgb <= "000000";
					when "10100000001110001" => rgb <= "000000";
					when "10100000001110010" => rgb <= "000000";
					when "10100000001110011" => rgb <= "000000";
					when "10100000001110100" => rgb <= "000000";
					when "10100000001110101" => rgb <= "000000";
					when "10100000001110110" => rgb <= "000000";
					when "10100000001110111" => rgb <= "000000";
					when "10100000001111000" => rgb <= "000000";
					when "10100000001111001" => rgb <= "000000";
					when "10100000001111010" => rgb <= "000000";
					when "10100000001111011" => rgb <= "000000";
					when "10100000001111100" => rgb <= "000000";
					when "10100000001111101" => rgb <= "000000";
					when "10100000001111110" => rgb <= "000000";
					when "10100000001111111" => rgb <= "000000";
					when "10100000010000000" => rgb <= "000000";
					when "10100000010000001" => rgb <= "000000";
					when "10100000010000010" => rgb <= "000000";
					when "10100000010000011" => rgb <= "000000";
					when "10100000010000100" => rgb <= "000000";
					when "10100000010000101" => rgb <= "000000";
					when "10100000010000110" => rgb <= "000000";
					when "10100000010000111" => rgb <= "000000";
					when "10100000010001000" => rgb <= "000000";
					when "10100000010001001" => rgb <= "000000";
					when "10100000010001010" => rgb <= "000000";
					when "10100000010001011" => rgb <= "000000";
					when "10100000010001100" => rgb <= "000000";
					when "10100000010001101" => rgb <= "000000";
					when "10100000010001110" => rgb <= "000000";
					when "10100000010001111" => rgb <= "000000";
					when "10100000010010000" => rgb <= "000000";
					when "10100000010010001" => rgb <= "000000";
					when "10100000010010010" => rgb <= "000000";
					when "10100000010010011" => rgb <= "000000";
					when "10100000010010100" => rgb <= "000000";
					when "10100000010010101" => rgb <= "000000";
					when "10100000010010110" => rgb <= "000000";
					when "10100000010010111" => rgb <= "000000";
					when "10100000010011000" => rgb <= "000000";
					when "10100000010011001" => rgb <= "000000";
					when "10100000010011010" => rgb <= "000000";
					when "10100000010011011" => rgb <= "000000";
					when "10100000010011100" => rgb <= "000000";
					when "10100000010011101" => rgb <= "000000";
					when "10100000010011110" => rgb <= "000000";
					when "10100000010011111" => rgb <= "000000";
					when "10100000010100000" => rgb <= "000000";
					when "10100000010100001" => rgb <= "000000";
					when "10100000010100010" => rgb <= "000000";
					when "10100000010100011" => rgb <= "000000";
					when "10100000010100100" => rgb <= "000000";
					when "10100000010100101" => rgb <= "000000";
					when "10100000010100110" => rgb <= "000000";
					when "10100000010100111" => rgb <= "000000";
					when "10100000010101000" => rgb <= "000000";
					when "10100000010101001" => rgb <= "000000";
					when "10100000010101010" => rgb <= "000000";
					when "10100000010101011" => rgb <= "000000";
					when "10100000010101100" => rgb <= "000000";
					when "10100000010101101" => rgb <= "000000";
					when "10100000010101110" => rgb <= "000000";
					when "10100000010101111" => rgb <= "000000";
					when "10100000010110000" => rgb <= "000000";
					when "10100000010110001" => rgb <= "000000";
					when "10100000010110010" => rgb <= "000000";
					when "10100000010110011" => rgb <= "000000";
					when "10100000010110100" => rgb <= "000000";
					when "10100000010110101" => rgb <= "000000";
					when "10100000010110110" => rgb <= "000000";
					when "10100000010110111" => rgb <= "000000";
					when "10100000010111000" => rgb <= "000000";
					when "10100000010111001" => rgb <= "000000";
					when "10100000010111010" => rgb <= "000000";
					when "10100000010111011" => rgb <= "000000";
					when "10100000010111100" => rgb <= "000000";
					when "10100000010111101" => rgb <= "000000";
					when "10100000010111110" => rgb <= "000000";
					when "10100000010111111" => rgb <= "000000";
					when "10100000011000000" => rgb <= "000000";
					when "10100000011000001" => rgb <= "000000";
					when "10100000011000010" => rgb <= "000000";
					when "10100000011000011" => rgb <= "000000";
					when "10100000011000100" => rgb <= "000000";
					when "10100000011000101" => rgb <= "000000";
					when "10100000011000110" => rgb <= "000000";
					when "10100000011000111" => rgb <= "000000";
					when "10100000011001000" => rgb <= "000000";
					when "10100000011001001" => rgb <= "000000";
					when "10100000011001010" => rgb <= "000000";
					when "10100000011001011" => rgb <= "000000";
					when "10100000011001100" => rgb <= "000000";
					when "10100000011001101" => rgb <= "000000";
					when "10100000011001110" => rgb <= "000000";
					when "10100000011001111" => rgb <= "000000";
					when "10100000011010000" => rgb <= "000000";
					when "10100000011010001" => rgb <= "000000";
					when "10100000011010010" => rgb <= "000000";
					when "10100000011010011" => rgb <= "000000";
					when "10100000011010100" => rgb <= "000000";
					when "10100000011010101" => rgb <= "000000";
					when "10100000011010110" => rgb <= "000000";
					when "10100000011010111" => rgb <= "000000";
					when "10100000011011000" => rgb <= "000000";
					when "10100000011011001" => rgb <= "000000";
					when "10100000011011010" => rgb <= "000000";
					when "10100000011011011" => rgb <= "000000";
					when "10100000011011100" => rgb <= "000000";
					when "10100000011011101" => rgb <= "000000";
					when "10100000011011110" => rgb <= "000000";
					when "10100000011011111" => rgb <= "000000";
					when "10100000011100000" => rgb <= "000000";
					when "10100000011100001" => rgb <= "000000";
					when "10100000011100010" => rgb <= "000000";
					when "10100000011100011" => rgb <= "000000";
					when "10100000011100100" => rgb <= "000000";
					when "10100000011100101" => rgb <= "000000";
					when "10100000011100110" => rgb <= "000000";
					when "10100000011100111" => rgb <= "000000";
					when "10100000011101000" => rgb <= "000000";
					when "10100000011101001" => rgb <= "000000";
					when "10100000011101010" => rgb <= "000000";
					when "10100000011101011" => rgb <= "000000";
					when "10100000011101100" => rgb <= "000000";
					when "10100000011101101" => rgb <= "000000";
					when "10100000011101110" => rgb <= "000000";
					when "10100000011101111" => rgb <= "000000";
					when "10100000011110000" => rgb <= "000000";
					when "10100000011110001" => rgb <= "000000";
					when "10100000011110010" => rgb <= "000000";
					when "10100000011110011" => rgb <= "000000";
					when "10100000011110100" => rgb <= "000000";
					when "10100000011110101" => rgb <= "000000";
					when "10100000011110110" => rgb <= "000000";
					when "10100000011110111" => rgb <= "000000";
					when "10100000011111000" => rgb <= "000000";
					when "10100000011111001" => rgb <= "000000";
					when "10100000011111010" => rgb <= "000000";
					when "10100000011111011" => rgb <= "000000";
					when "10100000011111100" => rgb <= "000000";
					when "10100000011111101" => rgb <= "000000";
					when "10100000011111110" => rgb <= "000000";
					when "10100000011111111" => rgb <= "000000";
					when "10100000100000000" => rgb <= "000000";
					when "10100000100000001" => rgb <= "000000";
					when "10100000100000010" => rgb <= "000000";
					when "10100000100000011" => rgb <= "000000";
					when "10100000100000100" => rgb <= "000000";
					when "10100000100000101" => rgb <= "000000";
					when "10100000100000110" => rgb <= "000000";
					when "10100000100000111" => rgb <= "000000";
					when "10100000100001000" => rgb <= "000000";
					when "10100000100001001" => rgb <= "000000";
					when "10100000100001010" => rgb <= "000000";
					when "10100000100001011" => rgb <= "000000";
					when "10100000100001100" => rgb <= "000000";
					when "10100000100001101" => rgb <= "000000";
					when "10100000100001110" => rgb <= "000000";
					when "10100000100001111" => rgb <= "000000";
					when "10100000100010000" => rgb <= "000000";
					when "10100000100010001" => rgb <= "000000";
					when "10100000100010010" => rgb <= "000000";
					when "10100000100010011" => rgb <= "000000";
					when "10100000100010100" => rgb <= "000000";
					when "10100000100010101" => rgb <= "000000";
					when "10100000100010110" => rgb <= "000000";
					when "10100000100010111" => rgb <= "000000";
					when "10100000100011000" => rgb <= "000000";
					when "10100000100011001" => rgb <= "000000";
					when "10100000100011010" => rgb <= "000000";
					when "10100000100011011" => rgb <= "000000";
					when "10100000100011100" => rgb <= "000000";
					when "10100000100011101" => rgb <= "000000";
					when "10100000100011110" => rgb <= "000000";
					when "10100000100011111" => rgb <= "000000";
					when "10100000100100000" => rgb <= "000000";
					when "10100000100100001" => rgb <= "000000";
					when "10100000100100010" => rgb <= "000000";
					when "10100000100100011" => rgb <= "000000";
					when "10100000100100100" => rgb <= "000000";
					when "10100000100100101" => rgb <= "000000";
					when "10100000100100110" => rgb <= "000000";
					when "10100000100100111" => rgb <= "000000";
					when "10100000100101000" => rgb <= "000000";
					when "10100000100101001" => rgb <= "000000";
					when "10100000100101010" => rgb <= "000000";
					when "10100000100101011" => rgb <= "000000";
					when "10100000100101100" => rgb <= "000000";
					when "10100000100101101" => rgb <= "000000";
					when "10100000100101110" => rgb <= "000000";
					when "10100000100101111" => rgb <= "000000";
					when "10100000100110000" => rgb <= "000000";
					when "10100000100110001" => rgb <= "000000";
					when "10100000100110010" => rgb <= "000000";
					when "10100000100110011" => rgb <= "000000";
					when "10100000100110100" => rgb <= "000000";
					when "10100000100110101" => rgb <= "000000";
					when "10100000100110110" => rgb <= "000000";
					when "10100000100110111" => rgb <= "000000";
					when "10100000100111000" => rgb <= "000000";
					when "10100000100111001" => rgb <= "000000";
					when "10100000100111010" => rgb <= "000000";
					when "10100000100111011" => rgb <= "000000";
					when "10100000100111100" => rgb <= "000000";
					when "10100000100111101" => rgb <= "000000";
					when "10100000100111110" => rgb <= "000000";
					when "10100000100111111" => rgb <= "000000";
					when "10100001000000000" => rgb <= "000000";
					when "10100001000000001" => rgb <= "000000";
					when "10100001000000010" => rgb <= "000000";
					when "10100001000000011" => rgb <= "000000";
					when "10100001000000100" => rgb <= "000000";
					when "10100001000000101" => rgb <= "101010";
					when "10100001000000110" => rgb <= "101010";
					when "10100001000000111" => rgb <= "101010";
					when "10100001000001000" => rgb <= "101010";
					when "10100001000001001" => rgb <= "101010";
					when "10100001000001010" => rgb <= "101010";
					when "10100001000001011" => rgb <= "111111";
					when "10100001000001100" => rgb <= "010101";
					when "10100001000001101" => rgb <= "000000";
					when "10100001000001110" => rgb <= "000000";
					when "10100001000001111" => rgb <= "000000";
					when "10100001000010000" => rgb <= "000000";
					when "10100001000010001" => rgb <= "000000";
					when "10100001000010010" => rgb <= "000000";
					when "10100001000010011" => rgb <= "000000";
					when "10100001000010100" => rgb <= "000000";
					when "10100001000010101" => rgb <= "000000";
					when "10100001000010110" => rgb <= "000000";
					when "10100001000010111" => rgb <= "000000";
					when "10100001000011000" => rgb <= "000000";
					when "10100001000011001" => rgb <= "000000";
					when "10100001000011010" => rgb <= "000000";
					when "10100001000011011" => rgb <= "000000";
					when "10100001000011100" => rgb <= "000000";
					when "10100001000011101" => rgb <= "000000";
					when "10100001000011110" => rgb <= "000000";
					when "10100001000011111" => rgb <= "000000";
					when "10100001000100000" => rgb <= "000000";
					when "10100001000100001" => rgb <= "000000";
					when "10100001000100010" => rgb <= "000000";
					when "10100001000100011" => rgb <= "101010";
					when "10100001000100100" => rgb <= "111111";
					when "10100001000100101" => rgb <= "101010";
					when "10100001000100110" => rgb <= "101010";
					when "10100001000100111" => rgb <= "111111";
					when "10100001000101000" => rgb <= "101010";
					when "10100001000101001" => rgb <= "101010";
					when "10100001000101010" => rgb <= "101010";
					when "10100001000101011" => rgb <= "101010";
					when "10100001000101100" => rgb <= "101010";
					when "10100001000101101" => rgb <= "101010";
					when "10100001000101110" => rgb <= "101010";
					when "10100001000101111" => rgb <= "101010";
					when "10100001000110000" => rgb <= "101010";
					when "10100001000110001" => rgb <= "101010";
					when "10100001000110010" => rgb <= "000000";
					when "10100001000110011" => rgb <= "000000";
					when "10100001000110100" => rgb <= "000000";
					when "10100001000110101" => rgb <= "000000";
					when "10100001000110110" => rgb <= "000000";
					when "10100001000110111" => rgb <= "000000";
					when "10100001000111000" => rgb <= "000000";
					when "10100001000111001" => rgb <= "000000";
					when "10100001000111010" => rgb <= "000000";
					when "10100001000111011" => rgb <= "000000";
					when "10100001000111100" => rgb <= "000000";
					when "10100001000111101" => rgb <= "000000";
					when "10100001000111110" => rgb <= "000000";
					when "10100001000111111" => rgb <= "000000";
					when "10100001001000000" => rgb <= "000000";
					when "10100001001000001" => rgb <= "101010";
					when "10100001001000010" => rgb <= "111111";
					when "10100001001000011" => rgb <= "101010";
					when "10100001001000100" => rgb <= "101010";
					when "10100001001000101" => rgb <= "111111";
					when "10100001001000110" => rgb <= "101010";
					when "10100001001000111" => rgb <= "101010";
					when "10100001001001000" => rgb <= "101010";
					when "10100001001001001" => rgb <= "101010";
					when "10100001001001010" => rgb <= "101010";
					when "10100001001001011" => rgb <= "101010";
					when "10100001001001100" => rgb <= "101010";
					when "10100001001001101" => rgb <= "101010";
					when "10100001001001110" => rgb <= "101010";
					when "10100001001001111" => rgb <= "101010";
					when "10100001001010000" => rgb <= "101010";
					when "10100001001010001" => rgb <= "101010";
					when "10100001001010010" => rgb <= "101010";
					when "10100001001010011" => rgb <= "101010";
					when "10100001001010100" => rgb <= "111111";
					when "10100001001010101" => rgb <= "101010";
					when "10100001001010110" => rgb <= "101010";
					when "10100001001010111" => rgb <= "101010";
					when "10100001001011000" => rgb <= "000000";
					when "10100001001011001" => rgb <= "000000";
					when "10100001001011010" => rgb <= "000000";
					when "10100001001011011" => rgb <= "000000";
					when "10100001001011100" => rgb <= "000000";
					when "10100001001011101" => rgb <= "000000";
					when "10100001001011110" => rgb <= "000000";
					when "10100001001011111" => rgb <= "000000";
					when "10100001001100000" => rgb <= "000000";
					when "10100001001100001" => rgb <= "000000";
					when "10100001001100010" => rgb <= "000000";
					when "10100001001100011" => rgb <= "000000";
					when "10100001001100100" => rgb <= "000000";
					when "10100001001100101" => rgb <= "000000";
					when "10100001001100110" => rgb <= "010101";
					when "10100001001100111" => rgb <= "101010";
					when "10100001001101000" => rgb <= "101010";
					when "10100001001101001" => rgb <= "101010";
					when "10100001001101010" => rgb <= "101010";
					when "10100001001101011" => rgb <= "111111";
					when "10100001001101100" => rgb <= "111111";
					when "10100001001101101" => rgb <= "101010";
					when "10100001001101110" => rgb <= "000000";
					when "10100001001101111" => rgb <= "000000";
					when "10100001001110000" => rgb <= "000000";
					when "10100001001110001" => rgb <= "000000";
					when "10100001001110010" => rgb <= "000000";
					when "10100001001110011" => rgb <= "000000";
					when "10100001001110100" => rgb <= "000000";
					when "10100001001110101" => rgb <= "000000";
					when "10100001001110110" => rgb <= "000000";
					when "10100001001110111" => rgb <= "000000";
					when "10100001001111000" => rgb <= "000000";
					when "10100001001111001" => rgb <= "000000";
					when "10100001001111010" => rgb <= "000000";
					when "10100001001111011" => rgb <= "000000";
					when "10100001001111100" => rgb <= "000000";
					when "10100001001111101" => rgb <= "101010";
					when "10100001001111110" => rgb <= "111111";
					when "10100001001111111" => rgb <= "101010";
					when "10100001010000000" => rgb <= "101010";
					when "10100001010000001" => rgb <= "101010";
					when "10100001010000010" => rgb <= "101010";
					when "10100001010000011" => rgb <= "101010";
					when "10100001010000100" => rgb <= "101010";
					when "10100001010000101" => rgb <= "101010";
					when "10100001010000110" => rgb <= "101010";
					when "10100001010000111" => rgb <= "101010";
					when "10100001010001000" => rgb <= "101010";
					when "10100001010001001" => rgb <= "101010";
					when "10100001010001010" => rgb <= "101010";
					when "10100001010001011" => rgb <= "101010";
					when "10100001010001100" => rgb <= "000000";
					when "10100001010001101" => rgb <= "000000";
					when "10100001010001110" => rgb <= "000000";
					when "10100001010001111" => rgb <= "000000";
					when "10100001010010000" => rgb <= "000000";
					when "10100001010010001" => rgb <= "000000";
					when "10100001010010010" => rgb <= "000000";
					when "10100001010010011" => rgb <= "000000";
					when "10100001010010100" => rgb <= "000000";
					when "10100001010010101" => rgb <= "000000";
					when "10100001010010110" => rgb <= "000000";
					when "10100001010010111" => rgb <= "000000";
					when "10100001010011000" => rgb <= "000000";
					when "10100001010011001" => rgb <= "000000";
					when "10100001010011010" => rgb <= "000000";
					when "10100001010011011" => rgb <= "000000";
					when "10100001010011100" => rgb <= "000000";
					when "10100001010011101" => rgb <= "000000";
					when "10100001010011110" => rgb <= "000000";
					when "10100001010011111" => rgb <= "000000";
					when "10100001010100000" => rgb <= "000000";
					when "10100001010100001" => rgb <= "000000";
					when "10100001010100010" => rgb <= "010101";
					when "10100001010100011" => rgb <= "101010";
					when "10100001010100100" => rgb <= "101010";
					when "10100001010100101" => rgb <= "101010";
					when "10100001010100110" => rgb <= "111111";
					when "10100001010100111" => rgb <= "101010";
					when "10100001010101000" => rgb <= "101010";
					when "10100001010101001" => rgb <= "101010";
					when "10100001010101010" => rgb <= "000000";
					when "10100001010101011" => rgb <= "000000";
					when "10100001010101100" => rgb <= "000000";
					when "10100001010101101" => rgb <= "000000";
					when "10100001010101110" => rgb <= "000000";
					when "10100001010101111" => rgb <= "000000";
					when "10100001010110000" => rgb <= "000000";
					when "10100001010110001" => rgb <= "000000";
					when "10100001010110010" => rgb <= "000000";
					when "10100001010110011" => rgb <= "000000";
					when "10100001010110100" => rgb <= "000000";
					when "10100001010110101" => rgb <= "000000";
					when "10100001010110110" => rgb <= "000000";
					when "10100001010110111" => rgb <= "000000";
					when "10100001010111000" => rgb <= "000000";
					when "10100001010111001" => rgb <= "000000";
					when "10100001010111010" => rgb <= "000000";
					when "10100001010111011" => rgb <= "000000";
					when "10100001010111100" => rgb <= "000000";
					when "10100001010111101" => rgb <= "000000";
					when "10100001010111110" => rgb <= "000000";
					when "10100001010111111" => rgb <= "000000";
					when "10100001011000000" => rgb <= "010101";
					when "10100001011000001" => rgb <= "101010";
					when "10100001011000010" => rgb <= "111111";
					when "10100001011000011" => rgb <= "101010";
					when "10100001011000100" => rgb <= "101010";
					when "10100001011000101" => rgb <= "101010";
					when "10100001011000110" => rgb <= "101010";
					when "10100001011000111" => rgb <= "101010";
					when "10100001011001000" => rgb <= "101010";
					when "10100001011001001" => rgb <= "111111";
					when "10100001011001010" => rgb <= "101010";
					when "10100001011001011" => rgb <= "101010";
					when "10100001011001100" => rgb <= "111111";
					when "10100001011001101" => rgb <= "101010";
					when "10100001011001110" => rgb <= "101010";
					when "10100001011001111" => rgb <= "101010";
					when "10100001011010000" => rgb <= "000000";
					when "10100001011010001" => rgb <= "000000";
					when "10100001011010010" => rgb <= "000000";
					when "10100001011010011" => rgb <= "000000";
					when "10100001011010100" => rgb <= "000000";
					when "10100001011010101" => rgb <= "000000";
					when "10100001011010110" => rgb <= "000000";
					when "10100001011010111" => rgb <= "101010";
					when "10100001011011000" => rgb <= "101010";
					when "10100001011011001" => rgb <= "101010";
					when "10100001011011010" => rgb <= "101010";
					when "10100001011011011" => rgb <= "101010";
					when "10100001011011100" => rgb <= "101010";
					when "10100001011011101" => rgb <= "101010";
					when "10100001011011110" => rgb <= "101010";
					when "10100001011011111" => rgb <= "101010";
					when "10100001011100000" => rgb <= "111111";
					when "10100001011100001" => rgb <= "101010";
					when "10100001011100010" => rgb <= "111111";
					when "10100001011100011" => rgb <= "111111";
					when "10100001011100100" => rgb <= "101010";
					when "10100001011100101" => rgb <= "101010";
					when "10100001011100110" => rgb <= "000000";
					when "10100001011100111" => rgb <= "000000";
					when "10100001011101000" => rgb <= "000000";
					when "10100001011101001" => rgb <= "000000";
					when "10100001011101010" => rgb <= "000000";
					when "10100001011101011" => rgb <= "000000";
					when "10100001011101100" => rgb <= "000000";
					when "10100001011101101" => rgb <= "010101";
					when "10100001011101110" => rgb <= "101010";
					when "10100001011101111" => rgb <= "101010";
					when "10100001011110000" => rgb <= "111111";
					when "10100001011110001" => rgb <= "101010";
					when "10100001011110010" => rgb <= "101010";
					when "10100001011110011" => rgb <= "111111";
					when "10100001011110100" => rgb <= "101010";
					when "10100001011110101" => rgb <= "000000";
					when "10100001011110110" => rgb <= "000000";
					when "10100001011110111" => rgb <= "000000";
					when "10100001011111000" => rgb <= "000000";
					when "10100001011111001" => rgb <= "000000";
					when "10100001011111010" => rgb <= "000000";
					when "10100001011111011" => rgb <= "000000";
					when "10100001011111100" => rgb <= "000000";
					when "10100001011111101" => rgb <= "000000";
					when "10100001011111110" => rgb <= "000000";
					when "10100001011111111" => rgb <= "000000";
					when "10100001100000000" => rgb <= "000000";
					when "10100001100000001" => rgb <= "000000";
					when "10100001100000010" => rgb <= "000000";
					when "10100001100000011" => rgb <= "000000";
					when "10100001100000100" => rgb <= "000000";
					when "10100001100000101" => rgb <= "000000";
					when "10100001100000110" => rgb <= "000000";
					when "10100001100000111" => rgb <= "000000";
					when "10100001100001000" => rgb <= "000000";
					when "10100001100001001" => rgb <= "000000";
					when "10100001100001010" => rgb <= "000000";
					when "10100001100001011" => rgb <= "010101";
					when "10100001100001100" => rgb <= "101010";
					when "10100001100001101" => rgb <= "101010";
					when "10100001100001110" => rgb <= "101010";
					when "10100001100001111" => rgb <= "101010";
					when "10100001100010000" => rgb <= "101010";
					when "10100001100010001" => rgb <= "101010";
					when "10100001100010010" => rgb <= "101010";
					when "10100001100010011" => rgb <= "101010";
					when "10100001100010100" => rgb <= "101010";
					when "10100001100010101" => rgb <= "101010";
					when "10100001100010110" => rgb <= "101010";
					when "10100001100010111" => rgb <= "101010";
					when "10100001100011000" => rgb <= "101010";
					when "10100001100011001" => rgb <= "101010";
					when "10100001100011010" => rgb <= "010101";
					when "10100001100011011" => rgb <= "000000";
					when "10100001100011100" => rgb <= "000000";
					when "10100001100011101" => rgb <= "000000";
					when "10100001100011110" => rgb <= "000000";
					when "10100001100011111" => rgb <= "000000";
					when "10100001100100000" => rgb <= "000000";
					when "10100001100100001" => rgb <= "000000";
					when "10100001100100010" => rgb <= "101010";
					when "10100001100100011" => rgb <= "111111";
					when "10100001100100100" => rgb <= "101010";
					when "10100001100100101" => rgb <= "111111";
					when "10100001100100110" => rgb <= "101010";
					when "10100001100100111" => rgb <= "101010";
					when "10100001100101000" => rgb <= "101010";
					when "10100001100101001" => rgb <= "101010";
					when "10100001100101010" => rgb <= "101010";
					when "10100001100101011" => rgb <= "101010";
					when "10100001100101100" => rgb <= "101010";
					when "10100001100101101" => rgb <= "101010";
					when "10100001100101110" => rgb <= "101010";
					when "10100001100101111" => rgb <= "101010";
					when "10100001100110000" => rgb <= "111111";
					when "10100001100110001" => rgb <= "000000";
					when "10100001100110010" => rgb <= "000000";
					when "10100001100110011" => rgb <= "000000";
					when "10100001100110100" => rgb <= "000000";
					when "10100001100110101" => rgb <= "000000";
					when "10100001100110110" => rgb <= "000000";
					when "10100001100110111" => rgb <= "000000";
					when "10100001100111000" => rgb <= "000000";
					when "10100001100111001" => rgb <= "000000";
					when "10100001100111010" => rgb <= "000000";
					when "10100001100111011" => rgb <= "000000";
					when "10100001100111100" => rgb <= "000000";
					when "10100001100111101" => rgb <= "000000";
					when "10100001100111110" => rgb <= "000000";
					when "10100001100111111" => rgb <= "000000";
					when "10100010000000000" => rgb <= "000000";
					when "10100010000000001" => rgb <= "000000";
					when "10100010000000010" => rgb <= "000000";
					when "10100010000000011" => rgb <= "000000";
					when "10100010000000100" => rgb <= "000000";
					when "10100010000000101" => rgb <= "101010";
					when "10100010000000110" => rgb <= "111111";
					when "10100010000000111" => rgb <= "111111";
					when "10100010000001000" => rgb <= "111111";
					when "10100010000001001" => rgb <= "111111";
					when "10100010000001010" => rgb <= "101010";
					when "10100010000001011" => rgb <= "111111";
					when "10100010000001100" => rgb <= "010101";
					when "10100010000001101" => rgb <= "000000";
					when "10100010000001110" => rgb <= "000000";
					when "10100010000001111" => rgb <= "000000";
					when "10100010000010000" => rgb <= "000000";
					when "10100010000010001" => rgb <= "000000";
					when "10100010000010010" => rgb <= "000000";
					when "10100010000010011" => rgb <= "000000";
					when "10100010000010100" => rgb <= "000000";
					when "10100010000010101" => rgb <= "000000";
					when "10100010000010110" => rgb <= "000000";
					when "10100010000010111" => rgb <= "000000";
					when "10100010000011000" => rgb <= "000000";
					when "10100010000011001" => rgb <= "000000";
					when "10100010000011010" => rgb <= "000000";
					when "10100010000011011" => rgb <= "000000";
					when "10100010000011100" => rgb <= "000000";
					when "10100010000011101" => rgb <= "000000";
					when "10100010000011110" => rgb <= "000000";
					when "10100010000011111" => rgb <= "000000";
					when "10100010000100000" => rgb <= "000000";
					when "10100010000100001" => rgb <= "000000";
					when "10100010000100010" => rgb <= "000000";
					when "10100010000100011" => rgb <= "101010";
					when "10100010000100100" => rgb <= "111111";
					when "10100010000100101" => rgb <= "111111";
					when "10100010000100110" => rgb <= "101010";
					when "10100010000100111" => rgb <= "111111";
					when "10100010000101000" => rgb <= "111111";
					when "10100010000101001" => rgb <= "111111";
					when "10100010000101010" => rgb <= "111111";
					when "10100010000101011" => rgb <= "111111";
					when "10100010000101100" => rgb <= "111111";
					when "10100010000101101" => rgb <= "111111";
					when "10100010000101110" => rgb <= "111111";
					when "10100010000101111" => rgb <= "111111";
					when "10100010000110000" => rgb <= "101010";
					when "10100010000110001" => rgb <= "111111";
					when "10100010000110010" => rgb <= "000000";
					when "10100010000110011" => rgb <= "000000";
					when "10100010000110100" => rgb <= "000000";
					when "10100010000110101" => rgb <= "000000";
					when "10100010000110110" => rgb <= "000000";
					when "10100010000110111" => rgb <= "000000";
					when "10100010000111000" => rgb <= "000000";
					when "10100010000111001" => rgb <= "000000";
					when "10100010000111010" => rgb <= "000000";
					when "10100010000111011" => rgb <= "000000";
					when "10100010000111100" => rgb <= "000000";
					when "10100010000111101" => rgb <= "000000";
					when "10100010000111110" => rgb <= "000000";
					when "10100010000111111" => rgb <= "000000";
					when "10100010001000000" => rgb <= "000000";
					when "10100010001000001" => rgb <= "101010";
					when "10100010001000010" => rgb <= "101010";
					when "10100010001000011" => rgb <= "111111";
					when "10100010001000100" => rgb <= "101010";
					when "10100010001000101" => rgb <= "101010";
					when "10100010001000110" => rgb <= "111111";
					when "10100010001000111" => rgb <= "111111";
					when "10100010001001000" => rgb <= "111111";
					when "10100010001001001" => rgb <= "111111";
					when "10100010001001010" => rgb <= "111111";
					when "10100010001001011" => rgb <= "111111";
					when "10100010001001100" => rgb <= "111111";
					when "10100010001001101" => rgb <= "111111";
					when "10100010001001110" => rgb <= "111111";
					when "10100010001001111" => rgb <= "111111";
					when "10100010001010000" => rgb <= "111111";
					when "10100010001010001" => rgb <= "101010";
					when "10100010001010010" => rgb <= "111111";
					when "10100010001010011" => rgb <= "111111";
					when "10100010001010100" => rgb <= "101010";
					when "10100010001010101" => rgb <= "111111";
					when "10100010001010110" => rgb <= "101010";
					when "10100010001010111" => rgb <= "010101";
					when "10100010001011000" => rgb <= "000000";
					when "10100010001011001" => rgb <= "000000";
					when "10100010001011010" => rgb <= "000000";
					when "10100010001011011" => rgb <= "000000";
					when "10100010001011100" => rgb <= "000000";
					when "10100010001011101" => rgb <= "000000";
					when "10100010001011110" => rgb <= "000000";
					when "10100010001011111" => rgb <= "000000";
					when "10100010001100000" => rgb <= "000000";
					when "10100010001100001" => rgb <= "000000";
					when "10100010001100010" => rgb <= "000000";
					when "10100010001100011" => rgb <= "000000";
					when "10100010001100100" => rgb <= "000000";
					when "10100010001100101" => rgb <= "000000";
					when "10100010001100110" => rgb <= "010101";
					when "10100010001100111" => rgb <= "111111";
					when "10100010001101000" => rgb <= "101010";
					when "10100010001101001" => rgb <= "111111";
					when "10100010001101010" => rgb <= "101010";
					when "10100010001101011" => rgb <= "101010";
					when "10100010001101100" => rgb <= "101010";
					when "10100010001101101" => rgb <= "111111";
					when "10100010001101110" => rgb <= "000000";
					when "10100010001101111" => rgb <= "000000";
					when "10100010001110000" => rgb <= "000000";
					when "10100010001110001" => rgb <= "000000";
					when "10100010001110010" => rgb <= "000000";
					when "10100010001110011" => rgb <= "000000";
					when "10100010001110100" => rgb <= "000000";
					when "10100010001110101" => rgb <= "000000";
					when "10100010001110110" => rgb <= "000000";
					when "10100010001110111" => rgb <= "000000";
					when "10100010001111000" => rgb <= "000000";
					when "10100010001111001" => rgb <= "000000";
					when "10100010001111010" => rgb <= "000000";
					when "10100010001111011" => rgb <= "000000";
					when "10100010001111100" => rgb <= "000000";
					when "10100010001111101" => rgb <= "101010";
					when "10100010001111110" => rgb <= "111111";
					when "10100010001111111" => rgb <= "101010";
					when "10100010010000000" => rgb <= "111111";
					when "10100010010000001" => rgb <= "111111";
					when "10100010010000010" => rgb <= "111111";
					when "10100010010000011" => rgb <= "111111";
					when "10100010010000100" => rgb <= "111111";
					when "10100010010000101" => rgb <= "111111";
					when "10100010010000110" => rgb <= "111111";
					when "10100010010000111" => rgb <= "111111";
					when "10100010010001000" => rgb <= "111111";
					when "10100010010001001" => rgb <= "101010";
					when "10100010010001010" => rgb <= "111111";
					when "10100010010001011" => rgb <= "111111";
					when "10100010010001100" => rgb <= "000000";
					when "10100010010001101" => rgb <= "000000";
					when "10100010010001110" => rgb <= "000000";
					when "10100010010001111" => rgb <= "000000";
					when "10100010010010000" => rgb <= "000000";
					when "10100010010010001" => rgb <= "000000";
					when "10100010010010010" => rgb <= "000000";
					when "10100010010010011" => rgb <= "000000";
					when "10100010010010100" => rgb <= "000000";
					when "10100010010010101" => rgb <= "000000";
					when "10100010010010110" => rgb <= "000000";
					when "10100010010010111" => rgb <= "000000";
					when "10100010010011000" => rgb <= "000000";
					when "10100010010011001" => rgb <= "000000";
					when "10100010010011010" => rgb <= "000000";
					when "10100010010011011" => rgb <= "000000";
					when "10100010010011100" => rgb <= "000000";
					when "10100010010011101" => rgb <= "000000";
					when "10100010010011110" => rgb <= "000000";
					when "10100010010011111" => rgb <= "000000";
					when "10100010010100000" => rgb <= "000000";
					when "10100010010100001" => rgb <= "000000";
					when "10100010010100010" => rgb <= "010101";
					when "10100010010100011" => rgb <= "111111";
					when "10100010010100100" => rgb <= "101010";
					when "10100010010100101" => rgb <= "101010";
					when "10100010010100110" => rgb <= "111111";
					when "10100010010100111" => rgb <= "101010";
					when "10100010010101000" => rgb <= "101010";
					when "10100010010101001" => rgb <= "111111";
					when "10100010010101010" => rgb <= "000000";
					when "10100010010101011" => rgb <= "000000";
					when "10100010010101100" => rgb <= "000000";
					when "10100010010101101" => rgb <= "000000";
					when "10100010010101110" => rgb <= "000000";
					when "10100010010101111" => rgb <= "000000";
					when "10100010010110000" => rgb <= "000000";
					when "10100010010110001" => rgb <= "000000";
					when "10100010010110010" => rgb <= "000000";
					when "10100010010110011" => rgb <= "000000";
					when "10100010010110100" => rgb <= "000000";
					when "10100010010110101" => rgb <= "000000";
					when "10100010010110110" => rgb <= "000000";
					when "10100010010110111" => rgb <= "000000";
					when "10100010010111000" => rgb <= "000000";
					when "10100010010111001" => rgb <= "000000";
					when "10100010010111010" => rgb <= "000000";
					when "10100010010111011" => rgb <= "000000";
					when "10100010010111100" => rgb <= "000000";
					when "10100010010111101" => rgb <= "000000";
					when "10100010010111110" => rgb <= "000000";
					when "10100010010111111" => rgb <= "000000";
					when "10100010011000000" => rgb <= "010101";
					when "10100010011000001" => rgb <= "111111";
					when "10100010011000010" => rgb <= "101010";
					when "10100010011000011" => rgb <= "101010";
					when "10100010011000100" => rgb <= "111111";
					when "10100010011000101" => rgb <= "111111";
					when "10100010011000110" => rgb <= "101010";
					when "10100010011000111" => rgb <= "111111";
					when "10100010011001000" => rgb <= "101010";
					when "10100010011001001" => rgb <= "111111";
					when "10100010011001010" => rgb <= "111111";
					when "10100010011001011" => rgb <= "101010";
					when "10100010011001100" => rgb <= "111111";
					when "10100010011001101" => rgb <= "111111";
					when "10100010011001110" => rgb <= "101010";
					when "10100010011001111" => rgb <= "010101";
					when "10100010011010000" => rgb <= "000000";
					when "10100010011010001" => rgb <= "000000";
					when "10100010011010010" => rgb <= "000000";
					when "10100010011010011" => rgb <= "000000";
					when "10100010011010100" => rgb <= "000000";
					when "10100010011010101" => rgb <= "000000";
					when "10100010011010110" => rgb <= "000000";
					when "10100010011010111" => rgb <= "101010";
					when "10100010011011000" => rgb <= "111111";
					when "10100010011011001" => rgb <= "111111";
					when "10100010011011010" => rgb <= "101010";
					when "10100010011011011" => rgb <= "111111";
					when "10100010011011100" => rgb <= "111111";
					when "10100010011011101" => rgb <= "111111";
					when "10100010011011110" => rgb <= "111111";
					when "10100010011011111" => rgb <= "111111";
					when "10100010011100000" => rgb <= "111111";
					when "10100010011100001" => rgb <= "111111";
					when "10100010011100010" => rgb <= "101010";
					when "10100010011100011" => rgb <= "101010";
					when "10100010011100100" => rgb <= "101010";
					when "10100010011100101" => rgb <= "111111";
					when "10100010011100110" => rgb <= "000000";
					when "10100010011100111" => rgb <= "000000";
					when "10100010011101000" => rgb <= "000000";
					when "10100010011101001" => rgb <= "000000";
					when "10100010011101010" => rgb <= "000000";
					when "10100010011101011" => rgb <= "000000";
					when "10100010011101100" => rgb <= "000000";
					when "10100010011101101" => rgb <= "010101";
					when "10100010011101110" => rgb <= "111111";
					when "10100010011101111" => rgb <= "101010";
					when "10100010011110000" => rgb <= "111111";
					when "10100010011110001" => rgb <= "111111";
					when "10100010011110010" => rgb <= "111111";
					when "10100010011110011" => rgb <= "101010";
					when "10100010011110100" => rgb <= "101010";
					when "10100010011110101" => rgb <= "000000";
					when "10100010011110110" => rgb <= "000000";
					when "10100010011110111" => rgb <= "000000";
					when "10100010011111000" => rgb <= "000000";
					when "10100010011111001" => rgb <= "000000";
					when "10100010011111010" => rgb <= "000000";
					when "10100010011111011" => rgb <= "000000";
					when "10100010011111100" => rgb <= "000000";
					when "10100010011111101" => rgb <= "000000";
					when "10100010011111110" => rgb <= "000000";
					when "10100010011111111" => rgb <= "000000";
					when "10100010100000000" => rgb <= "000000";
					when "10100010100000001" => rgb <= "000000";
					when "10100010100000010" => rgb <= "000000";
					when "10100010100000011" => rgb <= "000000";
					when "10100010100000100" => rgb <= "000000";
					when "10100010100000101" => rgb <= "000000";
					when "10100010100000110" => rgb <= "000000";
					when "10100010100000111" => rgb <= "000000";
					when "10100010100001000" => rgb <= "000000";
					when "10100010100001001" => rgb <= "000000";
					when "10100010100001010" => rgb <= "000000";
					when "10100010100001011" => rgb <= "010101";
					when "10100010100001100" => rgb <= "111111";
					when "10100010100001101" => rgb <= "101010";
					when "10100010100001110" => rgb <= "111111";
					when "10100010100001111" => rgb <= "111111";
					when "10100010100010000" => rgb <= "111111";
					when "10100010100010001" => rgb <= "111111";
					when "10100010100010010" => rgb <= "111111";
					when "10100010100010011" => rgb <= "111111";
					when "10100010100010100" => rgb <= "111111";
					when "10100010100010101" => rgb <= "111111";
					when "10100010100010110" => rgb <= "111111";
					when "10100010100010111" => rgb <= "111111";
					when "10100010100011000" => rgb <= "101010";
					when "10100010100011001" => rgb <= "111111";
					when "10100010100011010" => rgb <= "101010";
					when "10100010100011011" => rgb <= "000000";
					when "10100010100011100" => rgb <= "000000";
					when "10100010100011101" => rgb <= "000000";
					when "10100010100011110" => rgb <= "000000";
					when "10100010100011111" => rgb <= "000000";
					when "10100010100100000" => rgb <= "000000";
					when "10100010100100001" => rgb <= "000000";
					when "10100010100100010" => rgb <= "101010";
					when "10100010100100011" => rgb <= "101010";
					when "10100010100100100" => rgb <= "101010";
					when "10100010100100101" => rgb <= "111111";
					when "10100010100100110" => rgb <= "111111";
					when "10100010100100111" => rgb <= "111111";
					when "10100010100101000" => rgb <= "111111";
					when "10100010100101001" => rgb <= "111111";
					when "10100010100101010" => rgb <= "111111";
					when "10100010100101011" => rgb <= "111111";
					when "10100010100101100" => rgb <= "111111";
					when "10100010100101101" => rgb <= "111111";
					when "10100010100101110" => rgb <= "111111";
					when "10100010100101111" => rgb <= "101010";
					when "10100010100110000" => rgb <= "101010";
					when "10100010100110001" => rgb <= "000000";
					when "10100010100110010" => rgb <= "000000";
					when "10100010100110011" => rgb <= "000000";
					when "10100010100110100" => rgb <= "000000";
					when "10100010100110101" => rgb <= "000000";
					when "10100010100110110" => rgb <= "000000";
					when "10100010100110111" => rgb <= "000000";
					when "10100010100111000" => rgb <= "000000";
					when "10100010100111001" => rgb <= "000000";
					when "10100010100111010" => rgb <= "000000";
					when "10100010100111011" => rgb <= "000000";
					when "10100010100111100" => rgb <= "000000";
					when "10100010100111101" => rgb <= "000000";
					when "10100010100111110" => rgb <= "000000";
					when "10100010100111111" => rgb <= "000000";
					when "10100011000000000" => rgb <= "000000";
					when "10100011000000001" => rgb <= "000000";
					when "10100011000000010" => rgb <= "000000";
					when "10100011000000011" => rgb <= "000000";
					when "10100011000000100" => rgb <= "000000";
					when "10100011000000101" => rgb <= "101010";
					when "10100011000000110" => rgb <= "101010";
					when "10100011000000111" => rgb <= "101010";
					when "10100011000001000" => rgb <= "101010";
					when "10100011000001001" => rgb <= "111111";
					when "10100011000001010" => rgb <= "101010";
					when "10100011000001011" => rgb <= "101010";
					when "10100011000001100" => rgb <= "010101";
					when "10100011000001101" => rgb <= "000000";
					when "10100011000001110" => rgb <= "000000";
					when "10100011000001111" => rgb <= "000000";
					when "10100011000010000" => rgb <= "000000";
					when "10100011000010001" => rgb <= "000000";
					when "10100011000010010" => rgb <= "000000";
					when "10100011000010011" => rgb <= "000000";
					when "10100011000010100" => rgb <= "000000";
					when "10100011000010101" => rgb <= "000000";
					when "10100011000010110" => rgb <= "000000";
					when "10100011000010111" => rgb <= "000000";
					when "10100011000011000" => rgb <= "000000";
					when "10100011000011001" => rgb <= "000000";
					when "10100011000011010" => rgb <= "000000";
					when "10100011000011011" => rgb <= "000000";
					when "10100011000011100" => rgb <= "000000";
					when "10100011000011101" => rgb <= "000000";
					when "10100011000011110" => rgb <= "000000";
					when "10100011000011111" => rgb <= "000000";
					when "10100011000100000" => rgb <= "000000";
					when "10100011000100001" => rgb <= "000000";
					when "10100011000100010" => rgb <= "000000";
					when "10100011000100011" => rgb <= "101010";
					when "10100011000100100" => rgb <= "111111";
					when "10100011000100101" => rgb <= "101010";
					when "10100011000100110" => rgb <= "111111";
					when "10100011000100111" => rgb <= "111111";
					when "10100011000101000" => rgb <= "111111";
					when "10100011000101001" => rgb <= "111111";
					when "10100011000101010" => rgb <= "111111";
					when "10100011000101011" => rgb <= "111111";
					when "10100011000101100" => rgb <= "111111";
					when "10100011000101101" => rgb <= "101010";
					when "10100011000101110" => rgb <= "101010";
					when "10100011000101111" => rgb <= "101010";
					when "10100011000110000" => rgb <= "111111";
					when "10100011000110001" => rgb <= "101010";
					when "10100011000110010" => rgb <= "000000";
					when "10100011000110011" => rgb <= "000000";
					when "10100011000110100" => rgb <= "000000";
					when "10100011000110101" => rgb <= "000000";
					when "10100011000110110" => rgb <= "000000";
					when "10100011000110111" => rgb <= "000000";
					when "10100011000111000" => rgb <= "000000";
					when "10100011000111001" => rgb <= "000000";
					when "10100011000111010" => rgb <= "000000";
					when "10100011000111011" => rgb <= "000000";
					when "10100011000111100" => rgb <= "000000";
					when "10100011000111101" => rgb <= "000000";
					when "10100011000111110" => rgb <= "000000";
					when "10100011000111111" => rgb <= "000000";
					when "10100011001000000" => rgb <= "000000";
					when "10100011001000001" => rgb <= "101010";
					when "10100011001000010" => rgb <= "101010";
					when "10100011001000011" => rgb <= "111111";
					when "10100011001000100" => rgb <= "101010";
					when "10100011001000101" => rgb <= "111111";
					when "10100011001000110" => rgb <= "111111";
					when "10100011001000111" => rgb <= "101010";
					when "10100011001001000" => rgb <= "111111";
					when "10100011001001001" => rgb <= "111111";
					when "10100011001001010" => rgb <= "111111";
					when "10100011001001011" => rgb <= "111111";
					when "10100011001001100" => rgb <= "111111";
					when "10100011001001101" => rgb <= "111111";
					when "10100011001001110" => rgb <= "111111";
					when "10100011001001111" => rgb <= "111111";
					when "10100011001010000" => rgb <= "111111";
					when "10100011001010001" => rgb <= "101010";
					when "10100011001010010" => rgb <= "111111";
					when "10100011001010011" => rgb <= "111111";
					when "10100011001010100" => rgb <= "101010";
					when "10100011001010101" => rgb <= "101010";
					when "10100011001010110" => rgb <= "111111";
					when "10100011001010111" => rgb <= "101010";
					when "10100011001011000" => rgb <= "000000";
					when "10100011001011001" => rgb <= "000000";
					when "10100011001011010" => rgb <= "000000";
					when "10100011001011011" => rgb <= "000000";
					when "10100011001011100" => rgb <= "000000";
					when "10100011001011101" => rgb <= "000000";
					when "10100011001011110" => rgb <= "000000";
					when "10100011001011111" => rgb <= "000000";
					when "10100011001100000" => rgb <= "000000";
					when "10100011001100001" => rgb <= "000000";
					when "10100011001100010" => rgb <= "000000";
					when "10100011001100011" => rgb <= "000000";
					when "10100011001100100" => rgb <= "000000";
					when "10100011001100101" => rgb <= "000000";
					when "10100011001100110" => rgb <= "010101";
					when "10100011001100111" => rgb <= "111111";
					when "10100011001101000" => rgb <= "101010";
					when "10100011001101001" => rgb <= "111111";
					when "10100011001101010" => rgb <= "111111";
					when "10100011001101011" => rgb <= "101010";
					when "10100011001101100" => rgb <= "111111";
					when "10100011001101101" => rgb <= "111111";
					when "10100011001101110" => rgb <= "000000";
					when "10100011001101111" => rgb <= "000000";
					when "10100011001110000" => rgb <= "000000";
					when "10100011001110001" => rgb <= "000000";
					when "10100011001110010" => rgb <= "000000";
					when "10100011001110011" => rgb <= "000000";
					when "10100011001110100" => rgb <= "000000";
					when "10100011001110101" => rgb <= "000000";
					when "10100011001110110" => rgb <= "000000";
					when "10100011001110111" => rgb <= "000000";
					when "10100011001111000" => rgb <= "000000";
					when "10100011001111001" => rgb <= "000000";
					when "10100011001111010" => rgb <= "000000";
					when "10100011001111011" => rgb <= "000000";
					when "10100011001111100" => rgb <= "000000";
					when "10100011001111101" => rgb <= "101010";
					when "10100011001111110" => rgb <= "101010";
					when "10100011001111111" => rgb <= "101010";
					when "10100011010000000" => rgb <= "111111";
					when "10100011010000001" => rgb <= "111111";
					when "10100011010000010" => rgb <= "111111";
					when "10100011010000011" => rgb <= "111111";
					when "10100011010000100" => rgb <= "111111";
					when "10100011010000101" => rgb <= "111111";
					when "10100011010000110" => rgb <= "111111";
					when "10100011010000111" => rgb <= "111111";
					when "10100011010001000" => rgb <= "111111";
					when "10100011010001001" => rgb <= "101010";
					when "10100011010001010" => rgb <= "101010";
					when "10100011010001011" => rgb <= "101010";
					when "10100011010001100" => rgb <= "000000";
					when "10100011010001101" => rgb <= "000000";
					when "10100011010001110" => rgb <= "000000";
					when "10100011010001111" => rgb <= "000000";
					when "10100011010010000" => rgb <= "000000";
					when "10100011010010001" => rgb <= "000000";
					when "10100011010010010" => rgb <= "000000";
					when "10100011010010011" => rgb <= "000000";
					when "10100011010010100" => rgb <= "000000";
					when "10100011010010101" => rgb <= "000000";
					when "10100011010010110" => rgb <= "000000";
					when "10100011010010111" => rgb <= "000000";
					when "10100011010011000" => rgb <= "000000";
					when "10100011010011001" => rgb <= "000000";
					when "10100011010011010" => rgb <= "000000";
					when "10100011010011011" => rgb <= "000000";
					when "10100011010011100" => rgb <= "000000";
					when "10100011010011101" => rgb <= "000000";
					when "10100011010011110" => rgb <= "000000";
					when "10100011010011111" => rgb <= "000000";
					when "10100011010100000" => rgb <= "000000";
					when "10100011010100001" => rgb <= "000000";
					when "10100011010100010" => rgb <= "010101";
					when "10100011010100011" => rgb <= "111111";
					when "10100011010100100" => rgb <= "101010";
					when "10100011010100101" => rgb <= "111111";
					when "10100011010100110" => rgb <= "101010";
					when "10100011010100111" => rgb <= "101010";
					when "10100011010101000" => rgb <= "111111";
					when "10100011010101001" => rgb <= "101010";
					when "10100011010101010" => rgb <= "000000";
					when "10100011010101011" => rgb <= "000000";
					when "10100011010101100" => rgb <= "000000";
					when "10100011010101101" => rgb <= "000000";
					when "10100011010101110" => rgb <= "000000";
					when "10100011010101111" => rgb <= "000000";
					when "10100011010110000" => rgb <= "000000";
					when "10100011010110001" => rgb <= "000000";
					when "10100011010110010" => rgb <= "000000";
					when "10100011010110011" => rgb <= "000000";
					when "10100011010110100" => rgb <= "000000";
					when "10100011010110101" => rgb <= "000000";
					when "10100011010110110" => rgb <= "000000";
					when "10100011010110111" => rgb <= "000000";
					when "10100011010111000" => rgb <= "000000";
					when "10100011010111001" => rgb <= "000000";
					when "10100011010111010" => rgb <= "000000";
					when "10100011010111011" => rgb <= "000000";
					when "10100011010111100" => rgb <= "000000";
					when "10100011010111101" => rgb <= "000000";
					when "10100011010111110" => rgb <= "000000";
					when "10100011010111111" => rgb <= "000000";
					when "10100011011000000" => rgb <= "010101";
					when "10100011011000001" => rgb <= "111111";
					when "10100011011000010" => rgb <= "101010";
					when "10100011011000011" => rgb <= "111111";
					when "10100011011000100" => rgb <= "111111";
					when "10100011011000101" => rgb <= "101010";
					when "10100011011000110" => rgb <= "111111";
					when "10100011011000111" => rgb <= "111111";
					when "10100011011001000" => rgb <= "111111";
					when "10100011011001001" => rgb <= "111111";
					when "10100011011001010" => rgb <= "111111";
					when "10100011011001011" => rgb <= "111111";
					when "10100011011001100" => rgb <= "101010";
					when "10100011011001101" => rgb <= "101010";
					when "10100011011001110" => rgb <= "101010";
					when "10100011011001111" => rgb <= "010101";
					when "10100011011010000" => rgb <= "000000";
					when "10100011011010001" => rgb <= "000000";
					when "10100011011010010" => rgb <= "000000";
					when "10100011011010011" => rgb <= "000000";
					when "10100011011010100" => rgb <= "000000";
					when "10100011011010101" => rgb <= "000000";
					when "10100011011010110" => rgb <= "000000";
					when "10100011011010111" => rgb <= "101010";
					when "10100011011011000" => rgb <= "111111";
					when "10100011011011001" => rgb <= "101010";
					when "10100011011011010" => rgb <= "101010";
					when "10100011011011011" => rgb <= "111111";
					when "10100011011011100" => rgb <= "111111";
					when "10100011011011101" => rgb <= "111111";
					when "10100011011011110" => rgb <= "101010";
					when "10100011011011111" => rgb <= "111111";
					when "10100011011100000" => rgb <= "101010";
					when "10100011011100001" => rgb <= "111111";
					when "10100011011100010" => rgb <= "101010";
					when "10100011011100011" => rgb <= "111111";
					when "10100011011100100" => rgb <= "111111";
					when "10100011011100101" => rgb <= "101010";
					when "10100011011100110" => rgb <= "000000";
					when "10100011011100111" => rgb <= "000000";
					when "10100011011101000" => rgb <= "000000";
					when "10100011011101001" => rgb <= "000000";
					when "10100011011101010" => rgb <= "000000";
					when "10100011011101011" => rgb <= "000000";
					when "10100011011101100" => rgb <= "000000";
					when "10100011011101101" => rgb <= "010101";
					when "10100011011101110" => rgb <= "101010";
					when "10100011011101111" => rgb <= "111111";
					when "10100011011110000" => rgb <= "101010";
					when "10100011011110001" => rgb <= "101010";
					when "10100011011110010" => rgb <= "101010";
					when "10100011011110011" => rgb <= "111111";
					when "10100011011110100" => rgb <= "101010";
					when "10100011011110101" => rgb <= "000000";
					when "10100011011110110" => rgb <= "000000";
					when "10100011011110111" => rgb <= "000000";
					when "10100011011111000" => rgb <= "000000";
					when "10100011011111001" => rgb <= "000000";
					when "10100011011111010" => rgb <= "000000";
					when "10100011011111011" => rgb <= "000000";
					when "10100011011111100" => rgb <= "000000";
					when "10100011011111101" => rgb <= "000000";
					when "10100011011111110" => rgb <= "000000";
					when "10100011011111111" => rgb <= "000000";
					when "10100011100000000" => rgb <= "000000";
					when "10100011100000001" => rgb <= "000000";
					when "10100011100000010" => rgb <= "000000";
					when "10100011100000011" => rgb <= "000000";
					when "10100011100000100" => rgb <= "000000";
					when "10100011100000101" => rgb <= "000000";
					when "10100011100000110" => rgb <= "000000";
					when "10100011100000111" => rgb <= "000000";
					when "10100011100001000" => rgb <= "000000";
					when "10100011100001001" => rgb <= "000000";
					when "10100011100001010" => rgb <= "000000";
					when "10100011100001011" => rgb <= "010101";
					when "10100011100001100" => rgb <= "101010";
					when "10100011100001101" => rgb <= "101010";
					when "10100011100001110" => rgb <= "111111";
					when "10100011100001111" => rgb <= "111111";
					when "10100011100010000" => rgb <= "111111";
					when "10100011100010001" => rgb <= "111111";
					when "10100011100010010" => rgb <= "111111";
					when "10100011100010011" => rgb <= "111111";
					when "10100011100010100" => rgb <= "111111";
					when "10100011100010101" => rgb <= "111111";
					when "10100011100010110" => rgb <= "111111";
					when "10100011100010111" => rgb <= "111111";
					when "10100011100011000" => rgb <= "101010";
					when "10100011100011001" => rgb <= "101010";
					when "10100011100011010" => rgb <= "010101";
					when "10100011100011011" => rgb <= "000000";
					when "10100011100011100" => rgb <= "000000";
					when "10100011100011101" => rgb <= "000000";
					when "10100011100011110" => rgb <= "000000";
					when "10100011100011111" => rgb <= "000000";
					when "10100011100100000" => rgb <= "000000";
					when "10100011100100001" => rgb <= "000000";
					when "10100011100100010" => rgb <= "101010";
					when "10100011100100011" => rgb <= "101010";
					when "10100011100100100" => rgb <= "111111";
					when "10100011100100101" => rgb <= "101010";
					when "10100011100100110" => rgb <= "101010";
					when "10100011100100111" => rgb <= "111111";
					when "10100011100101000" => rgb <= "111111";
					when "10100011100101001" => rgb <= "111111";
					when "10100011100101010" => rgb <= "111111";
					when "10100011100101011" => rgb <= "111111";
					when "10100011100101100" => rgb <= "111111";
					when "10100011100101101" => rgb <= "111111";
					when "10100011100101110" => rgb <= "101010";
					when "10100011100101111" => rgb <= "101010";
					when "10100011100110000" => rgb <= "111111";
					when "10100011100110001" => rgb <= "000000";
					when "10100011100110010" => rgb <= "000000";
					when "10100011100110011" => rgb <= "000000";
					when "10100011100110100" => rgb <= "000000";
					when "10100011100110101" => rgb <= "000000";
					when "10100011100110110" => rgb <= "000000";
					when "10100011100110111" => rgb <= "000000";
					when "10100011100111000" => rgb <= "000000";
					when "10100011100111001" => rgb <= "000000";
					when "10100011100111010" => rgb <= "000000";
					when "10100011100111011" => rgb <= "000000";
					when "10100011100111100" => rgb <= "000000";
					when "10100011100111101" => rgb <= "000000";
					when "10100011100111110" => rgb <= "000000";
					when "10100011100111111" => rgb <= "000000";
					when "10100100000000000" => rgb <= "000000";
					when "10100100000000001" => rgb <= "000000";
					when "10100100000000010" => rgb <= "000000";
					when "10100100000000011" => rgb <= "000000";
					when "10100100000000100" => rgb <= "000000";
					when "10100100000000101" => rgb <= "101010";
					when "10100100000000110" => rgb <= "111111";
					when "10100100000000111" => rgb <= "111111";
					when "10100100000001000" => rgb <= "111111";
					when "10100100000001001" => rgb <= "101010";
					when "10100100000001010" => rgb <= "111111";
					when "10100100000001011" => rgb <= "111111";
					when "10100100000001100" => rgb <= "010101";
					when "10100100000001101" => rgb <= "000000";
					when "10100100000001110" => rgb <= "000000";
					when "10100100000001111" => rgb <= "000000";
					when "10100100000010000" => rgb <= "000000";
					when "10100100000010001" => rgb <= "000000";
					when "10100100000010010" => rgb <= "000000";
					when "10100100000010011" => rgb <= "000000";
					when "10100100000010100" => rgb <= "000000";
					when "10100100000010101" => rgb <= "000000";
					when "10100100000010110" => rgb <= "000000";
					when "10100100000010111" => rgb <= "000000";
					when "10100100000011000" => rgb <= "000000";
					when "10100100000011001" => rgb <= "000000";
					when "10100100000011010" => rgb <= "000000";
					when "10100100000011011" => rgb <= "000000";
					when "10100100000011100" => rgb <= "000000";
					when "10100100000011101" => rgb <= "000000";
					when "10100100000011110" => rgb <= "000000";
					when "10100100000011111" => rgb <= "000000";
					when "10100100000100000" => rgb <= "000000";
					when "10100100000100001" => rgb <= "000000";
					when "10100100000100010" => rgb <= "000000";
					when "10100100000100011" => rgb <= "101010";
					when "10100100000100100" => rgb <= "111111";
					when "10100100000100101" => rgb <= "101010";
					when "10100100000100110" => rgb <= "111111";
					when "10100100000100111" => rgb <= "111111";
					when "10100100000101000" => rgb <= "111111";
					when "10100100000101001" => rgb <= "111111";
					when "10100100000101010" => rgb <= "111111";
					when "10100100000101011" => rgb <= "111111";
					when "10100100000101100" => rgb <= "111111";
					when "10100100000101101" => rgb <= "111111";
					when "10100100000101110" => rgb <= "111111";
					when "10100100000101111" => rgb <= "101010";
					when "10100100000110000" => rgb <= "111111";
					when "10100100000110001" => rgb <= "101010";
					when "10100100000110010" => rgb <= "000000";
					when "10100100000110011" => rgb <= "000000";
					when "10100100000110100" => rgb <= "000000";
					when "10100100000110101" => rgb <= "000000";
					when "10100100000110110" => rgb <= "000000";
					when "10100100000110111" => rgb <= "000000";
					when "10100100000111000" => rgb <= "000000";
					when "10100100000111001" => rgb <= "000000";
					when "10100100000111010" => rgb <= "000000";
					when "10100100000111011" => rgb <= "000000";
					when "10100100000111100" => rgb <= "000000";
					when "10100100000111101" => rgb <= "000000";
					when "10100100000111110" => rgb <= "000000";
					when "10100100000111111" => rgb <= "000000";
					when "10100100001000000" => rgb <= "000000";
					when "10100100001000001" => rgb <= "101010";
					when "10100100001000010" => rgb <= "111111";
					when "10100100001000011" => rgb <= "101010";
					when "10100100001000100" => rgb <= "101010";
					when "10100100001000101" => rgb <= "101010";
					when "10100100001000110" => rgb <= "101010";
					when "10100100001000111" => rgb <= "111111";
					when "10100100001001000" => rgb <= "111111";
					when "10100100001001001" => rgb <= "111111";
					when "10100100001001010" => rgb <= "111111";
					when "10100100001001011" => rgb <= "111111";
					when "10100100001001100" => rgb <= "111111";
					when "10100100001001101" => rgb <= "111111";
					when "10100100001001110" => rgb <= "111111";
					when "10100100001001111" => rgb <= "111111";
					when "10100100001010000" => rgb <= "111111";
					when "10100100001010001" => rgb <= "111111";
					when "10100100001010010" => rgb <= "101010";
					when "10100100001010011" => rgb <= "111111";
					when "10100100001010100" => rgb <= "111111";
					when "10100100001010101" => rgb <= "101010";
					when "10100100001010110" => rgb <= "101010";
					when "10100100001010111" => rgb <= "101010";
					when "10100100001011000" => rgb <= "000000";
					when "10100100001011001" => rgb <= "000000";
					when "10100100001011010" => rgb <= "000000";
					when "10100100001011011" => rgb <= "000000";
					when "10100100001011100" => rgb <= "000000";
					when "10100100001011101" => rgb <= "000000";
					when "10100100001011110" => rgb <= "000000";
					when "10100100001011111" => rgb <= "000000";
					when "10100100001100000" => rgb <= "000000";
					when "10100100001100001" => rgb <= "000000";
					when "10100100001100010" => rgb <= "000000";
					when "10100100001100011" => rgb <= "000000";
					when "10100100001100100" => rgb <= "000000";
					when "10100100001100101" => rgb <= "000000";
					when "10100100001100110" => rgb <= "010101";
					when "10100100001100111" => rgb <= "111111";
					when "10100100001101000" => rgb <= "111111";
					when "10100100001101001" => rgb <= "111111";
					when "10100100001101010" => rgb <= "101010";
					when "10100100001101011" => rgb <= "101010";
					when "10100100001101100" => rgb <= "111111";
					when "10100100001101101" => rgb <= "101010";
					when "10100100001101110" => rgb <= "000000";
					when "10100100001101111" => rgb <= "000000";
					when "10100100001110000" => rgb <= "000000";
					when "10100100001110001" => rgb <= "000000";
					when "10100100001110010" => rgb <= "000000";
					when "10100100001110011" => rgb <= "000000";
					when "10100100001110100" => rgb <= "000000";
					when "10100100001110101" => rgb <= "000000";
					when "10100100001110110" => rgb <= "000000";
					when "10100100001110111" => rgb <= "000000";
					when "10100100001111000" => rgb <= "000000";
					when "10100100001111001" => rgb <= "000000";
					when "10100100001111010" => rgb <= "000000";
					when "10100100001111011" => rgb <= "000000";
					when "10100100001111100" => rgb <= "000000";
					when "10100100001111101" => rgb <= "101010";
					when "10100100001111110" => rgb <= "111111";
					when "10100100001111111" => rgb <= "111111";
					when "10100100010000000" => rgb <= "111111";
					when "10100100010000001" => rgb <= "111111";
					when "10100100010000010" => rgb <= "111111";
					when "10100100010000011" => rgb <= "111111";
					when "10100100010000100" => rgb <= "111111";
					when "10100100010000101" => rgb <= "111111";
					when "10100100010000110" => rgb <= "111111";
					when "10100100010000111" => rgb <= "111111";
					when "10100100010001000" => rgb <= "111111";
					when "10100100010001001" => rgb <= "111111";
					when "10100100010001010" => rgb <= "111111";
					when "10100100010001011" => rgb <= "111111";
					when "10100100010001100" => rgb <= "000000";
					when "10100100010001101" => rgb <= "000000";
					when "10100100010001110" => rgb <= "000000";
					when "10100100010001111" => rgb <= "000000";
					when "10100100010010000" => rgb <= "000000";
					when "10100100010010001" => rgb <= "000000";
					when "10100100010010010" => rgb <= "000000";
					when "10100100010010011" => rgb <= "000000";
					when "10100100010010100" => rgb <= "000000";
					when "10100100010010101" => rgb <= "000000";
					when "10100100010010110" => rgb <= "000000";
					when "10100100010010111" => rgb <= "000000";
					when "10100100010011000" => rgb <= "000000";
					when "10100100010011001" => rgb <= "000000";
					when "10100100010011010" => rgb <= "000000";
					when "10100100010011011" => rgb <= "000000";
					when "10100100010011100" => rgb <= "000000";
					when "10100100010011101" => rgb <= "000000";
					when "10100100010011110" => rgb <= "000000";
					when "10100100010011111" => rgb <= "000000";
					when "10100100010100000" => rgb <= "000000";
					when "10100100010100001" => rgb <= "000000";
					when "10100100010100010" => rgb <= "010101";
					when "10100100010100011" => rgb <= "101010";
					when "10100100010100100" => rgb <= "101010";
					when "10100100010100101" => rgb <= "111111";
					when "10100100010100110" => rgb <= "101010";
					when "10100100010100111" => rgb <= "111111";
					when "10100100010101000" => rgb <= "101010";
					when "10100100010101001" => rgb <= "101010";
					when "10100100010101010" => rgb <= "000000";
					when "10100100010101011" => rgb <= "000000";
					when "10100100010101100" => rgb <= "000000";
					when "10100100010101101" => rgb <= "000000";
					when "10100100010101110" => rgb <= "000000";
					when "10100100010101111" => rgb <= "000000";
					when "10100100010110000" => rgb <= "000000";
					when "10100100010110001" => rgb <= "000000";
					when "10100100010110010" => rgb <= "000000";
					when "10100100010110011" => rgb <= "000000";
					when "10100100010110100" => rgb <= "000000";
					when "10100100010110101" => rgb <= "000000";
					when "10100100010110110" => rgb <= "000000";
					when "10100100010110111" => rgb <= "000000";
					when "10100100010111000" => rgb <= "000000";
					when "10100100010111001" => rgb <= "000000";
					when "10100100010111010" => rgb <= "000000";
					when "10100100010111011" => rgb <= "000000";
					when "10100100010111100" => rgb <= "000000";
					when "10100100010111101" => rgb <= "000000";
					when "10100100010111110" => rgb <= "000000";
					when "10100100010111111" => rgb <= "000000";
					when "10100100011000000" => rgb <= "010101";
					when "10100100011000001" => rgb <= "101010";
					when "10100100011000010" => rgb <= "101010";
					when "10100100011000011" => rgb <= "111111";
					when "10100100011000100" => rgb <= "101010";
					when "10100100011000101" => rgb <= "101010";
					when "10100100011000110" => rgb <= "111111";
					when "10100100011000111" => rgb <= "111111";
					when "10100100011001000" => rgb <= "111111";
					when "10100100011001001" => rgb <= "101010";
					when "10100100011001010" => rgb <= "101010";
					when "10100100011001011" => rgb <= "111111";
					when "10100100011001100" => rgb <= "111111";
					when "10100100011001101" => rgb <= "101010";
					when "10100100011001110" => rgb <= "101010";
					when "10100100011001111" => rgb <= "010101";
					when "10100100011010000" => rgb <= "000000";
					when "10100100011010001" => rgb <= "000000";
					when "10100100011010010" => rgb <= "000000";
					when "10100100011010011" => rgb <= "000000";
					when "10100100011010100" => rgb <= "000000";
					when "10100100011010101" => rgb <= "000000";
					when "10100100011010110" => rgb <= "000000";
					when "10100100011010111" => rgb <= "101010";
					when "10100100011011000" => rgb <= "111111";
					when "10100100011011001" => rgb <= "101010";
					when "10100100011011010" => rgb <= "101010";
					when "10100100011011011" => rgb <= "111111";
					when "10100100011011100" => rgb <= "111111";
					when "10100100011011101" => rgb <= "111111";
					when "10100100011011110" => rgb <= "111111";
					when "10100100011011111" => rgb <= "111111";
					when "10100100011100000" => rgb <= "111111";
					when "10100100011100001" => rgb <= "101010";
					when "10100100011100010" => rgb <= "111111";
					when "10100100011100011" => rgb <= "101010";
					when "10100100011100100" => rgb <= "111111";
					when "10100100011100101" => rgb <= "111111";
					when "10100100011100110" => rgb <= "000000";
					when "10100100011100111" => rgb <= "000000";
					when "10100100011101000" => rgb <= "000000";
					when "10100100011101001" => rgb <= "000000";
					when "10100100011101010" => rgb <= "000000";
					when "10100100011101011" => rgb <= "000000";
					when "10100100011101100" => rgb <= "000000";
					when "10100100011101101" => rgb <= "010101";
					when "10100100011101110" => rgb <= "111111";
					when "10100100011101111" => rgb <= "101010";
					when "10100100011110000" => rgb <= "111111";
					when "10100100011110001" => rgb <= "111111";
					when "10100100011110010" => rgb <= "101010";
					when "10100100011110011" => rgb <= "101010";
					when "10100100011110100" => rgb <= "101010";
					when "10100100011110101" => rgb <= "000000";
					when "10100100011110110" => rgb <= "000000";
					when "10100100011110111" => rgb <= "000000";
					when "10100100011111000" => rgb <= "000000";
					when "10100100011111001" => rgb <= "000000";
					when "10100100011111010" => rgb <= "000000";
					when "10100100011111011" => rgb <= "000000";
					when "10100100011111100" => rgb <= "000000";
					when "10100100011111101" => rgb <= "000000";
					when "10100100011111110" => rgb <= "000000";
					when "10100100011111111" => rgb <= "000000";
					when "10100100100000000" => rgb <= "000000";
					when "10100100100000001" => rgb <= "000000";
					when "10100100100000010" => rgb <= "000000";
					when "10100100100000011" => rgb <= "000000";
					when "10100100100000100" => rgb <= "000000";
					when "10100100100000101" => rgb <= "000000";
					when "10100100100000110" => rgb <= "000000";
					when "10100100100000111" => rgb <= "000000";
					when "10100100100001000" => rgb <= "000000";
					when "10100100100001001" => rgb <= "000000";
					when "10100100100001010" => rgb <= "000000";
					when "10100100100001011" => rgb <= "010101";
					when "10100100100001100" => rgb <= "111111";
					when "10100100100001101" => rgb <= "111111";
					when "10100100100001110" => rgb <= "111111";
					when "10100100100001111" => rgb <= "111111";
					when "10100100100010000" => rgb <= "111111";
					when "10100100100010001" => rgb <= "111111";
					when "10100100100010010" => rgb <= "111111";
					when "10100100100010011" => rgb <= "111111";
					when "10100100100010100" => rgb <= "111111";
					when "10100100100010101" => rgb <= "111111";
					when "10100100100010110" => rgb <= "111111";
					when "10100100100010111" => rgb <= "111111";
					when "10100100100011000" => rgb <= "101010";
					when "10100100100011001" => rgb <= "111111";
					when "10100100100011010" => rgb <= "010101";
					when "10100100100011011" => rgb <= "000000";
					when "10100100100011100" => rgb <= "000000";
					when "10100100100011101" => rgb <= "000000";
					when "10100100100011110" => rgb <= "000000";
					when "10100100100011111" => rgb <= "000000";
					when "10100100100100000" => rgb <= "000000";
					when "10100100100100001" => rgb <= "000000";
					when "10100100100100010" => rgb <= "101010";
					when "10100100100100011" => rgb <= "111111";
					when "10100100100100100" => rgb <= "101010";
					when "10100100100100101" => rgb <= "101010";
					when "10100100100100110" => rgb <= "111111";
					when "10100100100100111" => rgb <= "111111";
					when "10100100100101000" => rgb <= "111111";
					when "10100100100101001" => rgb <= "111111";
					when "10100100100101010" => rgb <= "111111";
					when "10100100100101011" => rgb <= "111111";
					when "10100100100101100" => rgb <= "111111";
					when "10100100100101101" => rgb <= "111111";
					when "10100100100101110" => rgb <= "101010";
					when "10100100100101111" => rgb <= "101010";
					when "10100100100110000" => rgb <= "101010";
					when "10100100100110001" => rgb <= "000000";
					when "10100100100110010" => rgb <= "000000";
					when "10100100100110011" => rgb <= "000000";
					when "10100100100110100" => rgb <= "000000";
					when "10100100100110101" => rgb <= "000000";
					when "10100100100110110" => rgb <= "000000";
					when "10100100100110111" => rgb <= "000000";
					when "10100100100111000" => rgb <= "000000";
					when "10100100100111001" => rgb <= "000000";
					when "10100100100111010" => rgb <= "000000";
					when "10100100100111011" => rgb <= "000000";
					when "10100100100111100" => rgb <= "000000";
					when "10100100100111101" => rgb <= "000000";
					when "10100100100111110" => rgb <= "000000";
					when "10100100100111111" => rgb <= "000000";
					when "10100101000000000" => rgb <= "000000";
					when "10100101000000001" => rgb <= "000000";
					when "10100101000000010" => rgb <= "000000";
					when "10100101000000011" => rgb <= "000000";
					when "10100101000000100" => rgb <= "000000";
					when "10100101000000101" => rgb <= "101010";
					when "10100101000000110" => rgb <= "101010";
					when "10100101000000111" => rgb <= "111111";
					when "10100101000001000" => rgb <= "111111";
					when "10100101000001001" => rgb <= "101010";
					when "10100101000001010" => rgb <= "101010";
					when "10100101000001011" => rgb <= "101010";
					when "10100101000001100" => rgb <= "010101";
					when "10100101000001101" => rgb <= "000000";
					when "10100101000001110" => rgb <= "000000";
					when "10100101000001111" => rgb <= "000000";
					when "10100101000010000" => rgb <= "000000";
					when "10100101000010001" => rgb <= "000000";
					when "10100101000010010" => rgb <= "000000";
					when "10100101000010011" => rgb <= "000000";
					when "10100101000010100" => rgb <= "000000";
					when "10100101000010101" => rgb <= "000000";
					when "10100101000010110" => rgb <= "000000";
					when "10100101000010111" => rgb <= "000000";
					when "10100101000011000" => rgb <= "000000";
					when "10100101000011001" => rgb <= "000000";
					when "10100101000011010" => rgb <= "000000";
					when "10100101000011011" => rgb <= "000000";
					when "10100101000011100" => rgb <= "000000";
					when "10100101000011101" => rgb <= "000000";
					when "10100101000011110" => rgb <= "000000";
					when "10100101000011111" => rgb <= "000000";
					when "10100101000100000" => rgb <= "000000";
					when "10100101000100001" => rgb <= "000000";
					when "10100101000100010" => rgb <= "000000";
					when "10100101000100011" => rgb <= "101010";
					when "10100101000100100" => rgb <= "101010";
					when "10100101000100101" => rgb <= "111111";
					when "10100101000100110" => rgb <= "111111";
					when "10100101000100111" => rgb <= "111111";
					when "10100101000101000" => rgb <= "111111";
					when "10100101000101001" => rgb <= "111111";
					when "10100101000101010" => rgb <= "111111";
					when "10100101000101011" => rgb <= "111111";
					when "10100101000101100" => rgb <= "111111";
					when "10100101000101101" => rgb <= "111111";
					when "10100101000101110" => rgb <= "111111";
					when "10100101000101111" => rgb <= "111111";
					when "10100101000110000" => rgb <= "111111";
					when "10100101000110001" => rgb <= "101010";
					when "10100101000110010" => rgb <= "000000";
					when "10100101000110011" => rgb <= "000000";
					when "10100101000110100" => rgb <= "000000";
					when "10100101000110101" => rgb <= "000000";
					when "10100101000110110" => rgb <= "000000";
					when "10100101000110111" => rgb <= "000000";
					when "10100101000111000" => rgb <= "000000";
					when "10100101000111001" => rgb <= "000000";
					when "10100101000111010" => rgb <= "000000";
					when "10100101000111011" => rgb <= "000000";
					when "10100101000111100" => rgb <= "000000";
					when "10100101000111101" => rgb <= "000000";
					when "10100101000111110" => rgb <= "000000";
					when "10100101000111111" => rgb <= "000000";
					when "10100101001000000" => rgb <= "000000";
					when "10100101001000001" => rgb <= "101010";
					when "10100101001000010" => rgb <= "101010";
					when "10100101001000011" => rgb <= "111111";
					when "10100101001000100" => rgb <= "111111";
					when "10100101001000101" => rgb <= "111111";
					when "10100101001000110" => rgb <= "101010";
					when "10100101001000111" => rgb <= "111111";
					when "10100101001001000" => rgb <= "101010";
					when "10100101001001001" => rgb <= "101010";
					when "10100101001001010" => rgb <= "101010";
					when "10100101001001011" => rgb <= "101010";
					when "10100101001001100" => rgb <= "101010";
					when "10100101001001101" => rgb <= "101010";
					when "10100101001001110" => rgb <= "101010";
					when "10100101001001111" => rgb <= "101010";
					when "10100101001010000" => rgb <= "101010";
					when "10100101001010001" => rgb <= "111111";
					when "10100101001010010" => rgb <= "101010";
					when "10100101001010011" => rgb <= "101010";
					when "10100101001010100" => rgb <= "111111";
					when "10100101001010101" => rgb <= "101010";
					when "10100101001010110" => rgb <= "101010";
					when "10100101001010111" => rgb <= "010101";
					when "10100101001011000" => rgb <= "000000";
					when "10100101001011001" => rgb <= "000000";
					when "10100101001011010" => rgb <= "000000";
					when "10100101001011011" => rgb <= "000000";
					when "10100101001011100" => rgb <= "000000";
					when "10100101001011101" => rgb <= "000000";
					when "10100101001011110" => rgb <= "000000";
					when "10100101001011111" => rgb <= "000000";
					when "10100101001100000" => rgb <= "000000";
					when "10100101001100001" => rgb <= "000000";
					when "10100101001100010" => rgb <= "000000";
					when "10100101001100011" => rgb <= "000000";
					when "10100101001100100" => rgb <= "000000";
					when "10100101001100101" => rgb <= "000000";
					when "10100101001100110" => rgb <= "010101";
					when "10100101001100111" => rgb <= "111111";
					when "10100101001101000" => rgb <= "111111";
					when "10100101001101001" => rgb <= "101010";
					when "10100101001101010" => rgb <= "111111";
					when "10100101001101011" => rgb <= "111111";
					when "10100101001101100" => rgb <= "101010";
					when "10100101001101101" => rgb <= "101010";
					when "10100101001101110" => rgb <= "000000";
					when "10100101001101111" => rgb <= "000000";
					when "10100101001110000" => rgb <= "000000";
					when "10100101001110001" => rgb <= "000000";
					when "10100101001110010" => rgb <= "000000";
					when "10100101001110011" => rgb <= "000000";
					when "10100101001110100" => rgb <= "000000";
					when "10100101001110101" => rgb <= "000000";
					when "10100101001110110" => rgb <= "000000";
					when "10100101001110111" => rgb <= "000000";
					when "10100101001111000" => rgb <= "000000";
					when "10100101001111001" => rgb <= "000000";
					when "10100101001111010" => rgb <= "000000";
					when "10100101001111011" => rgb <= "000000";
					when "10100101001111100" => rgb <= "000000";
					when "10100101001111101" => rgb <= "101010";
					when "10100101001111110" => rgb <= "101010";
					when "10100101001111111" => rgb <= "111111";
					when "10100101010000000" => rgb <= "111111";
					when "10100101010000001" => rgb <= "111111";
					when "10100101010000010" => rgb <= "111111";
					when "10100101010000011" => rgb <= "111111";
					when "10100101010000100" => rgb <= "111111";
					when "10100101010000101" => rgb <= "111111";
					when "10100101010000110" => rgb <= "111111";
					when "10100101010000111" => rgb <= "111111";
					when "10100101010001000" => rgb <= "101010";
					when "10100101010001001" => rgb <= "101010";
					when "10100101010001010" => rgb <= "101010";
					when "10100101010001011" => rgb <= "111111";
					when "10100101010001100" => rgb <= "000000";
					when "10100101010001101" => rgb <= "000000";
					when "10100101010001110" => rgb <= "000000";
					when "10100101010001111" => rgb <= "000000";
					when "10100101010010000" => rgb <= "000000";
					when "10100101010010001" => rgb <= "000000";
					when "10100101010010010" => rgb <= "000000";
					when "10100101010010011" => rgb <= "000000";
					when "10100101010010100" => rgb <= "000000";
					when "10100101010010101" => rgb <= "000000";
					when "10100101010010110" => rgb <= "000000";
					when "10100101010010111" => rgb <= "000000";
					when "10100101010011000" => rgb <= "000000";
					when "10100101010011001" => rgb <= "000000";
					when "10100101010011010" => rgb <= "000000";
					when "10100101010011011" => rgb <= "000000";
					when "10100101010011100" => rgb <= "000000";
					when "10100101010011101" => rgb <= "000000";
					when "10100101010011110" => rgb <= "000000";
					when "10100101010011111" => rgb <= "000000";
					when "10100101010100000" => rgb <= "000000";
					when "10100101010100001" => rgb <= "000000";
					when "10100101010100010" => rgb <= "010101";
					when "10100101010100011" => rgb <= "111111";
					when "10100101010100100" => rgb <= "101010";
					when "10100101010100101" => rgb <= "111111";
					when "10100101010100110" => rgb <= "111111";
					when "10100101010100111" => rgb <= "101010";
					when "10100101010101000" => rgb <= "111111";
					when "10100101010101001" => rgb <= "111111";
					when "10100101010101010" => rgb <= "000000";
					when "10100101010101011" => rgb <= "000000";
					when "10100101010101100" => rgb <= "000000";
					when "10100101010101101" => rgb <= "000000";
					when "10100101010101110" => rgb <= "000000";
					when "10100101010101111" => rgb <= "000000";
					when "10100101010110000" => rgb <= "000000";
					when "10100101010110001" => rgb <= "000000";
					when "10100101010110010" => rgb <= "000000";
					when "10100101010110011" => rgb <= "000000";
					when "10100101010110100" => rgb <= "000000";
					when "10100101010110101" => rgb <= "000000";
					when "10100101010110110" => rgb <= "000000";
					when "10100101010110111" => rgb <= "000000";
					when "10100101010111000" => rgb <= "000000";
					when "10100101010111001" => rgb <= "000000";
					when "10100101010111010" => rgb <= "000000";
					when "10100101010111011" => rgb <= "000000";
					when "10100101010111100" => rgb <= "000000";
					when "10100101010111101" => rgb <= "000000";
					when "10100101010111110" => rgb <= "000000";
					when "10100101010111111" => rgb <= "000000";
					when "10100101011000000" => rgb <= "010101";
					when "10100101011000001" => rgb <= "111111";
					when "10100101011000010" => rgb <= "111111";
					when "10100101011000011" => rgb <= "101010";
					when "10100101011000100" => rgb <= "111111";
					when "10100101011000101" => rgb <= "111111";
					when "10100101011000110" => rgb <= "111111";
					when "10100101011000111" => rgb <= "111111";
					when "10100101011001000" => rgb <= "101010";
					when "10100101011001001" => rgb <= "101010";
					when "10100101011001010" => rgb <= "101010";
					when "10100101011001011" => rgb <= "111111";
					when "10100101011001100" => rgb <= "101010";
					when "10100101011001101" => rgb <= "101010";
					when "10100101011001110" => rgb <= "111111";
					when "10100101011001111" => rgb <= "010101";
					when "10100101011010000" => rgb <= "000000";
					when "10100101011010001" => rgb <= "000000";
					when "10100101011010010" => rgb <= "000000";
					when "10100101011010011" => rgb <= "000000";
					when "10100101011010100" => rgb <= "000000";
					when "10100101011010101" => rgb <= "000000";
					when "10100101011010110" => rgb <= "000000";
					when "10100101011010111" => rgb <= "101010";
					when "10100101011011000" => rgb <= "111111";
					when "10100101011011001" => rgb <= "101010";
					when "10100101011011010" => rgb <= "101010";
					when "10100101011011011" => rgb <= "111111";
					when "10100101011011100" => rgb <= "111111";
					when "10100101011011101" => rgb <= "111111";
					when "10100101011011110" => rgb <= "111111";
					when "10100101011011111" => rgb <= "111111";
					when "10100101011100000" => rgb <= "111111";
					when "10100101011100001" => rgb <= "101010";
					when "10100101011100010" => rgb <= "111111";
					when "10100101011100011" => rgb <= "111111";
					when "10100101011100100" => rgb <= "101010";
					when "10100101011100101" => rgb <= "101010";
					when "10100101011100110" => rgb <= "000000";
					when "10100101011100111" => rgb <= "000000";
					when "10100101011101000" => rgb <= "000000";
					when "10100101011101001" => rgb <= "000000";
					when "10100101011101010" => rgb <= "000000";
					when "10100101011101011" => rgb <= "000000";
					when "10100101011101100" => rgb <= "000000";
					when "10100101011101101" => rgb <= "010101";
					when "10100101011101110" => rgb <= "111111";
					when "10100101011101111" => rgb <= "101010";
					when "10100101011110000" => rgb <= "111111";
					when "10100101011110001" => rgb <= "111111";
					when "10100101011110010" => rgb <= "111111";
					when "10100101011110011" => rgb <= "101010";
					when "10100101011110100" => rgb <= "101010";
					when "10100101011110101" => rgb <= "000000";
					when "10100101011110110" => rgb <= "000000";
					when "10100101011110111" => rgb <= "000000";
					when "10100101011111000" => rgb <= "000000";
					when "10100101011111001" => rgb <= "000000";
					when "10100101011111010" => rgb <= "000000";
					when "10100101011111011" => rgb <= "000000";
					when "10100101011111100" => rgb <= "000000";
					when "10100101011111101" => rgb <= "000000";
					when "10100101011111110" => rgb <= "000000";
					when "10100101011111111" => rgb <= "000000";
					when "10100101100000000" => rgb <= "000000";
					when "10100101100000001" => rgb <= "000000";
					when "10100101100000010" => rgb <= "000000";
					when "10100101100000011" => rgb <= "000000";
					when "10100101100000100" => rgb <= "000000";
					when "10100101100000101" => rgb <= "000000";
					when "10100101100000110" => rgb <= "000000";
					when "10100101100000111" => rgb <= "000000";
					when "10100101100001000" => rgb <= "000000";
					when "10100101100001001" => rgb <= "000000";
					when "10100101100001010" => rgb <= "000000";
					when "10100101100001011" => rgb <= "010101";
					when "10100101100001100" => rgb <= "101010";
					when "10100101100001101" => rgb <= "101010";
					when "10100101100001110" => rgb <= "101010";
					when "10100101100001111" => rgb <= "111111";
					when "10100101100010000" => rgb <= "111111";
					when "10100101100010001" => rgb <= "111111";
					when "10100101100010010" => rgb <= "111111";
					when "10100101100010011" => rgb <= "111111";
					when "10100101100010100" => rgb <= "111111";
					when "10100101100010101" => rgb <= "111111";
					when "10100101100010110" => rgb <= "111111";
					when "10100101100010111" => rgb <= "111111";
					when "10100101100011000" => rgb <= "101010";
					when "10100101100011001" => rgb <= "111111";
					when "10100101100011010" => rgb <= "010101";
					when "10100101100011011" => rgb <= "000000";
					when "10100101100011100" => rgb <= "000000";
					when "10100101100011101" => rgb <= "000000";
					when "10100101100011110" => rgb <= "000000";
					when "10100101100011111" => rgb <= "000000";
					when "10100101100100000" => rgb <= "000000";
					when "10100101100100001" => rgb <= "000000";
					when "10100101100100010" => rgb <= "101010";
					when "10100101100100011" => rgb <= "111111";
					when "10100101100100100" => rgb <= "101010";
					when "10100101100100101" => rgb <= "111111";
					when "10100101100100110" => rgb <= "111111";
					when "10100101100100111" => rgb <= "101010";
					when "10100101100101000" => rgb <= "111111";
					when "10100101100101001" => rgb <= "111111";
					when "10100101100101010" => rgb <= "111111";
					when "10100101100101011" => rgb <= "111111";
					when "10100101100101100" => rgb <= "111111";
					when "10100101100101101" => rgb <= "111111";
					when "10100101100101110" => rgb <= "101010";
					when "10100101100101111" => rgb <= "101010";
					when "10100101100110000" => rgb <= "111111";
					when "10100101100110001" => rgb <= "000000";
					when "10100101100110010" => rgb <= "000000";
					when "10100101100110011" => rgb <= "000000";
					when "10100101100110100" => rgb <= "000000";
					when "10100101100110101" => rgb <= "000000";
					when "10100101100110110" => rgb <= "000000";
					when "10100101100110111" => rgb <= "000000";
					when "10100101100111000" => rgb <= "000000";
					when "10100101100111001" => rgb <= "000000";
					when "10100101100111010" => rgb <= "000000";
					when "10100101100111011" => rgb <= "000000";
					when "10100101100111100" => rgb <= "000000";
					when "10100101100111101" => rgb <= "000000";
					when "10100101100111110" => rgb <= "000000";
					when "10100101100111111" => rgb <= "000000";
					when "10100110000000000" => rgb <= "000000";
					when "10100110000000001" => rgb <= "000000";
					when "10100110000000010" => rgb <= "000000";
					when "10100110000000011" => rgb <= "000000";
					when "10100110000000100" => rgb <= "000000";
					when "10100110000000101" => rgb <= "101010";
					when "10100110000000110" => rgb <= "111111";
					when "10100110000000111" => rgb <= "101010";
					when "10100110000001000" => rgb <= "101010";
					when "10100110000001001" => rgb <= "111111";
					when "10100110000001010" => rgb <= "111111";
					when "10100110000001011" => rgb <= "111111";
					when "10100110000001100" => rgb <= "010101";
					when "10100110000001101" => rgb <= "000000";
					when "10100110000001110" => rgb <= "000000";
					when "10100110000001111" => rgb <= "000000";
					when "10100110000010000" => rgb <= "000000";
					when "10100110000010001" => rgb <= "000000";
					when "10100110000010010" => rgb <= "000000";
					when "10100110000010011" => rgb <= "000000";
					when "10100110000010100" => rgb <= "000000";
					when "10100110000010101" => rgb <= "000000";
					when "10100110000010110" => rgb <= "000000";
					when "10100110000010111" => rgb <= "000000";
					when "10100110000011000" => rgb <= "000000";
					when "10100110000011001" => rgb <= "000000";
					when "10100110000011010" => rgb <= "000000";
					when "10100110000011011" => rgb <= "000000";
					when "10100110000011100" => rgb <= "000000";
					when "10100110000011101" => rgb <= "000000";
					when "10100110000011110" => rgb <= "000000";
					when "10100110000011111" => rgb <= "000000";
					when "10100110000100000" => rgb <= "000000";
					when "10100110000100001" => rgb <= "000000";
					when "10100110000100010" => rgb <= "000000";
					when "10100110000100011" => rgb <= "101010";
					when "10100110000100100" => rgb <= "111111";
					when "10100110000100101" => rgb <= "101010";
					when "10100110000100110" => rgb <= "101010";
					when "10100110000100111" => rgb <= "111111";
					when "10100110000101000" => rgb <= "111111";
					when "10100110000101001" => rgb <= "111111";
					when "10100110000101010" => rgb <= "111111";
					when "10100110000101011" => rgb <= "111111";
					when "10100110000101100" => rgb <= "111111";
					when "10100110000101101" => rgb <= "111111";
					when "10100110000101110" => rgb <= "101010";
					when "10100110000101111" => rgb <= "101010";
					when "10100110000110000" => rgb <= "111111";
					when "10100110000110001" => rgb <= "101010";
					when "10100110000110010" => rgb <= "000000";
					when "10100110000110011" => rgb <= "000000";
					when "10100110000110100" => rgb <= "000000";
					when "10100110000110101" => rgb <= "000000";
					when "10100110000110110" => rgb <= "000000";
					when "10100110000110111" => rgb <= "000000";
					when "10100110000111000" => rgb <= "000000";
					when "10100110000111001" => rgb <= "000000";
					when "10100110000111010" => rgb <= "000000";
					when "10100110000111011" => rgb <= "000000";
					when "10100110000111100" => rgb <= "000000";
					when "10100110000111101" => rgb <= "000000";
					when "10100110000111110" => rgb <= "000000";
					when "10100110000111111" => rgb <= "000000";
					when "10100110001000000" => rgb <= "000000";
					when "10100110001000001" => rgb <= "101010";
					when "10100110001000010" => rgb <= "101010";
					when "10100110001000011" => rgb <= "101010";
					when "10100110001000100" => rgb <= "101010";
					when "10100110001000101" => rgb <= "101010";
					when "10100110001000110" => rgb <= "101010";
					when "10100110001000111" => rgb <= "101010";
					when "10100110001001000" => rgb <= "101010";
					when "10100110001001001" => rgb <= "101010";
					when "10100110001001010" => rgb <= "101010";
					when "10100110001001011" => rgb <= "101010";
					when "10100110001001100" => rgb <= "101010";
					when "10100110001001101" => rgb <= "101010";
					when "10100110001001110" => rgb <= "101010";
					when "10100110001001111" => rgb <= "101010";
					when "10100110001010000" => rgb <= "101010";
					when "10100110001010001" => rgb <= "111111";
					when "10100110001010010" => rgb <= "101010";
					when "10100110001010011" => rgb <= "101010";
					when "10100110001010100" => rgb <= "101010";
					when "10100110001010101" => rgb <= "101010";
					when "10100110001010110" => rgb <= "111111";
					when "10100110001010111" => rgb <= "010101";
					when "10100110001011000" => rgb <= "000000";
					when "10100110001011001" => rgb <= "000000";
					when "10100110001011010" => rgb <= "000000";
					when "10100110001011011" => rgb <= "000000";
					when "10100110001011100" => rgb <= "000000";
					when "10100110001011101" => rgb <= "000000";
					when "10100110001011110" => rgb <= "000000";
					when "10100110001011111" => rgb <= "000000";
					when "10100110001100000" => rgb <= "000000";
					when "10100110001100001" => rgb <= "000000";
					when "10100110001100010" => rgb <= "000000";
					when "10100110001100011" => rgb <= "000000";
					when "10100110001100100" => rgb <= "000000";
					when "10100110001100101" => rgb <= "000000";
					when "10100110001100110" => rgb <= "010101";
					when "10100110001100111" => rgb <= "101010";
					when "10100110001101000" => rgb <= "101010";
					when "10100110001101001" => rgb <= "101010";
					when "10100110001101010" => rgb <= "111111";
					when "10100110001101011" => rgb <= "111111";
					when "10100110001101100" => rgb <= "111111";
					when "10100110001101101" => rgb <= "111111";
					when "10100110001101110" => rgb <= "000000";
					when "10100110001101111" => rgb <= "000000";
					when "10100110001110000" => rgb <= "000000";
					when "10100110001110001" => rgb <= "000000";
					when "10100110001110010" => rgb <= "000000";
					when "10100110001110011" => rgb <= "000000";
					when "10100110001110100" => rgb <= "000000";
					when "10100110001110101" => rgb <= "000000";
					when "10100110001110110" => rgb <= "000000";
					when "10100110001110111" => rgb <= "000000";
					when "10100110001111000" => rgb <= "000000";
					when "10100110001111001" => rgb <= "000000";
					when "10100110001111010" => rgb <= "000000";
					when "10100110001111011" => rgb <= "000000";
					when "10100110001111100" => rgb <= "000000";
					when "10100110001111101" => rgb <= "101010";
					when "10100110001111110" => rgb <= "111111";
					when "10100110001111111" => rgb <= "101010";
					when "10100110010000000" => rgb <= "111111";
					when "10100110010000001" => rgb <= "111111";
					when "10100110010000010" => rgb <= "111111";
					when "10100110010000011" => rgb <= "111111";
					when "10100110010000100" => rgb <= "111111";
					when "10100110010000101" => rgb <= "111111";
					when "10100110010000110" => rgb <= "111111";
					when "10100110010000111" => rgb <= "111111";
					when "10100110010001000" => rgb <= "101010";
					when "10100110010001001" => rgb <= "111111";
					when "10100110010001010" => rgb <= "111111";
					when "10100110010001011" => rgb <= "101010";
					when "10100110010001100" => rgb <= "000000";
					when "10100110010001101" => rgb <= "000000";
					when "10100110010001110" => rgb <= "000000";
					when "10100110010001111" => rgb <= "000000";
					when "10100110010010000" => rgb <= "000000";
					when "10100110010010001" => rgb <= "000000";
					when "10100110010010010" => rgb <= "000000";
					when "10100110010010011" => rgb <= "000000";
					when "10100110010010100" => rgb <= "000000";
					when "10100110010010101" => rgb <= "000000";
					when "10100110010010110" => rgb <= "000000";
					when "10100110010010111" => rgb <= "000000";
					when "10100110010011000" => rgb <= "000000";
					when "10100110010011001" => rgb <= "000000";
					when "10100110010011010" => rgb <= "000000";
					when "10100110010011011" => rgb <= "000000";
					when "10100110010011100" => rgb <= "000000";
					when "10100110010011101" => rgb <= "000000";
					when "10100110010011110" => rgb <= "000000";
					when "10100110010011111" => rgb <= "000000";
					when "10100110010100000" => rgb <= "000000";
					when "10100110010100001" => rgb <= "000000";
					when "10100110010100010" => rgb <= "010101";
					when "10100110010100011" => rgb <= "101010";
					when "10100110010100100" => rgb <= "101010";
					when "10100110010100101" => rgb <= "111111";
					when "10100110010100110" => rgb <= "111111";
					when "10100110010100111" => rgb <= "101010";
					when "10100110010101000" => rgb <= "101010";
					when "10100110010101001" => rgb <= "111111";
					when "10100110010101010" => rgb <= "000000";
					when "10100110010101011" => rgb <= "000000";
					when "10100110010101100" => rgb <= "000000";
					when "10100110010101101" => rgb <= "000000";
					when "10100110010101110" => rgb <= "000000";
					when "10100110010101111" => rgb <= "000000";
					when "10100110010110000" => rgb <= "000000";
					when "10100110010110001" => rgb <= "000000";
					when "10100110010110010" => rgb <= "000000";
					when "10100110010110011" => rgb <= "000000";
					when "10100110010110100" => rgb <= "000000";
					when "10100110010110101" => rgb <= "000000";
					when "10100110010110110" => rgb <= "000000";
					when "10100110010110111" => rgb <= "000000";
					when "10100110010111000" => rgb <= "000000";
					when "10100110010111001" => rgb <= "000000";
					when "10100110010111010" => rgb <= "000000";
					when "10100110010111011" => rgb <= "000000";
					when "10100110010111100" => rgb <= "000000";
					when "10100110010111101" => rgb <= "000000";
					when "10100110010111110" => rgb <= "000000";
					when "10100110010111111" => rgb <= "000000";
					when "10100110011000000" => rgb <= "010101";
					when "10100110011000001" => rgb <= "101010";
					when "10100110011000010" => rgb <= "101010";
					when "10100110011000011" => rgb <= "111111";
					when "10100110011000100" => rgb <= "111111";
					when "10100110011000101" => rgb <= "101010";
					when "10100110011000110" => rgb <= "101010";
					when "10100110011000111" => rgb <= "111111";
					when "10100110011001000" => rgb <= "101010";
					when "10100110011001001" => rgb <= "111111";
					when "10100110011001010" => rgb <= "111111";
					when "10100110011001011" => rgb <= "101010";
					when "10100110011001100" => rgb <= "101010";
					when "10100110011001101" => rgb <= "101010";
					when "10100110011001110" => rgb <= "111111";
					when "10100110011001111" => rgb <= "010101";
					when "10100110011010000" => rgb <= "000000";
					when "10100110011010001" => rgb <= "000000";
					when "10100110011010010" => rgb <= "000000";
					when "10100110011010011" => rgb <= "000000";
					when "10100110011010100" => rgb <= "000000";
					when "10100110011010101" => rgb <= "000000";
					when "10100110011010110" => rgb <= "000000";
					when "10100110011010111" => rgb <= "101010";
					when "10100110011011000" => rgb <= "111111";
					when "10100110011011001" => rgb <= "101010";
					when "10100110011011010" => rgb <= "101010";
					when "10100110011011011" => rgb <= "111111";
					when "10100110011011100" => rgb <= "111111";
					when "10100110011011101" => rgb <= "111111";
					when "10100110011011110" => rgb <= "111111";
					when "10100110011011111" => rgb <= "111111";
					when "10100110011100000" => rgb <= "111111";
					when "10100110011100001" => rgb <= "111111";
					when "10100110011100010" => rgb <= "101010";
					when "10100110011100011" => rgb <= "111111";
					when "10100110011100100" => rgb <= "111111";
					when "10100110011100101" => rgb <= "101010";
					when "10100110011100110" => rgb <= "000000";
					when "10100110011100111" => rgb <= "000000";
					when "10100110011101000" => rgb <= "000000";
					when "10100110011101001" => rgb <= "000000";
					when "10100110011101010" => rgb <= "000000";
					when "10100110011101011" => rgb <= "000000";
					when "10100110011101100" => rgb <= "000000";
					when "10100110011101101" => rgb <= "010101";
					when "10100110011101110" => rgb <= "101010";
					when "10100110011101111" => rgb <= "101010";
					when "10100110011110000" => rgb <= "111111";
					when "10100110011110001" => rgb <= "101010";
					when "10100110011110010" => rgb <= "101010";
					when "10100110011110011" => rgb <= "101010";
					when "10100110011110100" => rgb <= "101010";
					when "10100110011110101" => rgb <= "000000";
					when "10100110011110110" => rgb <= "000000";
					when "10100110011110111" => rgb <= "000000";
					when "10100110011111000" => rgb <= "000000";
					when "10100110011111001" => rgb <= "000000";
					when "10100110011111010" => rgb <= "000000";
					when "10100110011111011" => rgb <= "000000";
					when "10100110011111100" => rgb <= "000000";
					when "10100110011111101" => rgb <= "000000";
					when "10100110011111110" => rgb <= "000000";
					when "10100110011111111" => rgb <= "000000";
					when "10100110100000000" => rgb <= "000000";
					when "10100110100000001" => rgb <= "000000";
					when "10100110100000010" => rgb <= "000000";
					when "10100110100000011" => rgb <= "000000";
					when "10100110100000100" => rgb <= "000000";
					when "10100110100000101" => rgb <= "000000";
					when "10100110100000110" => rgb <= "000000";
					when "10100110100000111" => rgb <= "000000";
					when "10100110100001000" => rgb <= "000000";
					when "10100110100001001" => rgb <= "000000";
					when "10100110100001010" => rgb <= "000000";
					when "10100110100001011" => rgb <= "010101";
					when "10100110100001100" => rgb <= "101010";
					when "10100110100001101" => rgb <= "101010";
					when "10100110100001110" => rgb <= "111111";
					when "10100110100001111" => rgb <= "111111";
					when "10100110100010000" => rgb <= "111111";
					when "10100110100010001" => rgb <= "111111";
					when "10100110100010010" => rgb <= "111111";
					when "10100110100010011" => rgb <= "111111";
					when "10100110100010100" => rgb <= "111111";
					when "10100110100010101" => rgb <= "111111";
					when "10100110100010110" => rgb <= "111111";
					when "10100110100010111" => rgb <= "111111";
					when "10100110100011000" => rgb <= "101010";
					when "10100110100011001" => rgb <= "101010";
					when "10100110100011010" => rgb <= "010101";
					when "10100110100011011" => rgb <= "000000";
					when "10100110100011100" => rgb <= "000000";
					when "10100110100011101" => rgb <= "000000";
					when "10100110100011110" => rgb <= "000000";
					when "10100110100011111" => rgb <= "000000";
					when "10100110100100000" => rgb <= "000000";
					when "10100110100100001" => rgb <= "000000";
					when "10100110100100010" => rgb <= "101010";
					when "10100110100100011" => rgb <= "111111";
					when "10100110100100100" => rgb <= "101010";
					when "10100110100100101" => rgb <= "111111";
					when "10100110100100110" => rgb <= "101010";
					when "10100110100100111" => rgb <= "111111";
					when "10100110100101000" => rgb <= "111111";
					when "10100110100101001" => rgb <= "111111";
					when "10100110100101010" => rgb <= "111111";
					when "10100110100101011" => rgb <= "111111";
					when "10100110100101100" => rgb <= "111111";
					when "10100110100101101" => rgb <= "111111";
					when "10100110100101110" => rgb <= "101010";
					when "10100110100101111" => rgb <= "101010";
					when "10100110100110000" => rgb <= "111111";
					when "10100110100110001" => rgb <= "000000";
					when "10100110100110010" => rgb <= "000000";
					when "10100110100110011" => rgb <= "000000";
					when "10100110100110100" => rgb <= "000000";
					when "10100110100110101" => rgb <= "000000";
					when "10100110100110110" => rgb <= "000000";
					when "10100110100110111" => rgb <= "000000";
					when "10100110100111000" => rgb <= "000000";
					when "10100110100111001" => rgb <= "000000";
					when "10100110100111010" => rgb <= "000000";
					when "10100110100111011" => rgb <= "000000";
					when "10100110100111100" => rgb <= "000000";
					when "10100110100111101" => rgb <= "000000";
					when "10100110100111110" => rgb <= "000000";
					when "10100110100111111" => rgb <= "000000";
					when "10100111000000000" => rgb <= "000000";
					when "10100111000000001" => rgb <= "000000";
					when "10100111000000010" => rgb <= "000000";
					when "10100111000000011" => rgb <= "000000";
					when "10100111000000100" => rgb <= "000000";
					when "10100111000000101" => rgb <= "101010";
					when "10100111000000110" => rgb <= "101010";
					when "10100111000000111" => rgb <= "101010";
					when "10100111000001000" => rgb <= "101010";
					when "10100111000001001" => rgb <= "111111";
					when "10100111000001010" => rgb <= "101010";
					when "10100111000001011" => rgb <= "111111";
					when "10100111000001100" => rgb <= "010101";
					when "10100111000001101" => rgb <= "000000";
					when "10100111000001110" => rgb <= "000000";
					when "10100111000001111" => rgb <= "000000";
					when "10100111000010000" => rgb <= "000000";
					when "10100111000010001" => rgb <= "000000";
					when "10100111000010010" => rgb <= "000000";
					when "10100111000010011" => rgb <= "000000";
					when "10100111000010100" => rgb <= "000000";
					when "10100111000010101" => rgb <= "000000";
					when "10100111000010110" => rgb <= "000000";
					when "10100111000010111" => rgb <= "000000";
					when "10100111000011000" => rgb <= "000000";
					when "10100111000011001" => rgb <= "000000";
					when "10100111000011010" => rgb <= "000000";
					when "10100111000011011" => rgb <= "000000";
					when "10100111000011100" => rgb <= "000000";
					when "10100111000011101" => rgb <= "000000";
					when "10100111000011110" => rgb <= "000000";
					when "10100111000011111" => rgb <= "000000";
					when "10100111000100000" => rgb <= "000000";
					when "10100111000100001" => rgb <= "000000";
					when "10100111000100010" => rgb <= "000000";
					when "10100111000100011" => rgb <= "101010";
					when "10100111000100100" => rgb <= "111111";
					when "10100111000100101" => rgb <= "101010";
					when "10100111000100110" => rgb <= "111111";
					when "10100111000100111" => rgb <= "101010";
					when "10100111000101000" => rgb <= "111111";
					when "10100111000101001" => rgb <= "111111";
					when "10100111000101010" => rgb <= "111111";
					when "10100111000101011" => rgb <= "111111";
					when "10100111000101100" => rgb <= "111111";
					when "10100111000101101" => rgb <= "111111";
					when "10100111000101110" => rgb <= "111111";
					when "10100111000101111" => rgb <= "111111";
					when "10100111000110000" => rgb <= "111111";
					when "10100111000110001" => rgb <= "101010";
					when "10100111000110010" => rgb <= "000000";
					when "10100111000110011" => rgb <= "000000";
					when "10100111000110100" => rgb <= "000000";
					when "10100111000110101" => rgb <= "000000";
					when "10100111000110110" => rgb <= "000000";
					when "10100111000110111" => rgb <= "000000";
					when "10100111000111000" => rgb <= "000000";
					when "10100111000111001" => rgb <= "000000";
					when "10100111000111010" => rgb <= "000000";
					when "10100111000111011" => rgb <= "000000";
					when "10100111000111100" => rgb <= "000000";
					when "10100111000111101" => rgb <= "000000";
					when "10100111000111110" => rgb <= "000000";
					when "10100111000111111" => rgb <= "000000";
					when "10100111001000000" => rgb <= "000000";
					when "10100111001000001" => rgb <= "101010";
					when "10100111001000010" => rgb <= "101010";
					when "10100111001000011" => rgb <= "111111";
					when "10100111001000100" => rgb <= "111111";
					when "10100111001000101" => rgb <= "111111";
					when "10100111001000110" => rgb <= "101010";
					when "10100111001000111" => rgb <= "111111";
					when "10100111001001000" => rgb <= "111111";
					when "10100111001001001" => rgb <= "111111";
					when "10100111001001010" => rgb <= "111111";
					when "10100111001001011" => rgb <= "111111";
					when "10100111001001100" => rgb <= "111111";
					when "10100111001001101" => rgb <= "111111";
					when "10100111001001110" => rgb <= "111111";
					when "10100111001001111" => rgb <= "111111";
					when "10100111001010000" => rgb <= "111111";
					when "10100111001010001" => rgb <= "111111";
					when "10100111001010010" => rgb <= "101010";
					when "10100111001010011" => rgb <= "111111";
					when "10100111001010100" => rgb <= "111111";
					when "10100111001010101" => rgb <= "101010";
					when "10100111001010110" => rgb <= "111111";
					when "10100111001010111" => rgb <= "010101";
					when "10100111001011000" => rgb <= "000000";
					when "10100111001011001" => rgb <= "000000";
					when "10100111001011010" => rgb <= "000000";
					when "10100111001011011" => rgb <= "000000";
					when "10100111001011100" => rgb <= "000000";
					when "10100111001011101" => rgb <= "000000";
					when "10100111001011110" => rgb <= "000000";
					when "10100111001011111" => rgb <= "000000";
					when "10100111001100000" => rgb <= "000000";
					when "10100111001100001" => rgb <= "000000";
					when "10100111001100010" => rgb <= "000000";
					when "10100111001100011" => rgb <= "000000";
					when "10100111001100100" => rgb <= "000000";
					when "10100111001100101" => rgb <= "000000";
					when "10100111001100110" => rgb <= "010101";
					when "10100111001100111" => rgb <= "111111";
					when "10100111001101000" => rgb <= "101010";
					when "10100111001101001" => rgb <= "111111";
					when "10100111001101010" => rgb <= "111111";
					when "10100111001101011" => rgb <= "101010";
					when "10100111001101100" => rgb <= "111111";
					when "10100111001101101" => rgb <= "101010";
					when "10100111001101110" => rgb <= "000000";
					when "10100111001101111" => rgb <= "000000";
					when "10100111001110000" => rgb <= "000000";
					when "10100111001110001" => rgb <= "000000";
					when "10100111001110010" => rgb <= "000000";
					when "10100111001110011" => rgb <= "000000";
					when "10100111001110100" => rgb <= "000000";
					when "10100111001110101" => rgb <= "000000";
					when "10100111001110110" => rgb <= "000000";
					when "10100111001110111" => rgb <= "000000";
					when "10100111001111000" => rgb <= "000000";
					when "10100111001111001" => rgb <= "000000";
					when "10100111001111010" => rgb <= "000000";
					when "10100111001111011" => rgb <= "000000";
					when "10100111001111100" => rgb <= "000000";
					when "10100111001111101" => rgb <= "101010";
					when "10100111001111110" => rgb <= "111111";
					when "10100111001111111" => rgb <= "111111";
					when "10100111010000000" => rgb <= "111111";
					when "10100111010000001" => rgb <= "111111";
					when "10100111010000010" => rgb <= "111111";
					when "10100111010000011" => rgb <= "111111";
					when "10100111010000100" => rgb <= "111111";
					when "10100111010000101" => rgb <= "111111";
					when "10100111010000110" => rgb <= "111111";
					when "10100111010000111" => rgb <= "111111";
					when "10100111010001000" => rgb <= "111111";
					when "10100111010001001" => rgb <= "101010";
					when "10100111010001010" => rgb <= "101010";
					when "10100111010001011" => rgb <= "111111";
					when "10100111010001100" => rgb <= "000000";
					when "10100111010001101" => rgb <= "000000";
					when "10100111010001110" => rgb <= "000000";
					when "10100111010001111" => rgb <= "000000";
					when "10100111010010000" => rgb <= "000000";
					when "10100111010010001" => rgb <= "000000";
					when "10100111010010010" => rgb <= "000000";
					when "10100111010010011" => rgb <= "000000";
					when "10100111010010100" => rgb <= "000000";
					when "10100111010010101" => rgb <= "000000";
					when "10100111010010110" => rgb <= "000000";
					when "10100111010010111" => rgb <= "000000";
					when "10100111010011000" => rgb <= "000000";
					when "10100111010011001" => rgb <= "000000";
					when "10100111010011010" => rgb <= "000000";
					when "10100111010011011" => rgb <= "000000";
					when "10100111010011100" => rgb <= "000000";
					when "10100111010011101" => rgb <= "000000";
					when "10100111010011110" => rgb <= "000000";
					when "10100111010011111" => rgb <= "000000";
					when "10100111010100000" => rgb <= "000000";
					when "10100111010100001" => rgb <= "000000";
					when "10100111010100010" => rgb <= "010101";
					when "10100111010100011" => rgb <= "111111";
					when "10100111010100100" => rgb <= "101010";
					when "10100111010100101" => rgb <= "111111";
					when "10100111010100110" => rgb <= "101010";
					when "10100111010100111" => rgb <= "111111";
					when "10100111010101000" => rgb <= "101010";
					when "10100111010101001" => rgb <= "111111";
					when "10100111010101010" => rgb <= "000000";
					when "10100111010101011" => rgb <= "000000";
					when "10100111010101100" => rgb <= "000000";
					when "10100111010101101" => rgb <= "000000";
					when "10100111010101110" => rgb <= "000000";
					when "10100111010101111" => rgb <= "000000";
					when "10100111010110000" => rgb <= "000000";
					when "10100111010110001" => rgb <= "000000";
					when "10100111010110010" => rgb <= "000000";
					when "10100111010110011" => rgb <= "000000";
					when "10100111010110100" => rgb <= "000000";
					when "10100111010110101" => rgb <= "000000";
					when "10100111010110110" => rgb <= "000000";
					when "10100111010110111" => rgb <= "000000";
					when "10100111010111000" => rgb <= "000000";
					when "10100111010111001" => rgb <= "000000";
					when "10100111010111010" => rgb <= "000000";
					when "10100111010111011" => rgb <= "000000";
					when "10100111010111100" => rgb <= "000000";
					when "10100111010111101" => rgb <= "000000";
					when "10100111010111110" => rgb <= "000000";
					when "10100111010111111" => rgb <= "000000";
					when "10100111011000000" => rgb <= "010101";
					when "10100111011000001" => rgb <= "111111";
					when "10100111011000010" => rgb <= "101010";
					when "10100111011000011" => rgb <= "111111";
					when "10100111011000100" => rgb <= "101010";
					when "10100111011000101" => rgb <= "111111";
					when "10100111011000110" => rgb <= "111111";
					when "10100111011000111" => rgb <= "101010";
					when "10100111011001000" => rgb <= "101010";
					when "10100111011001001" => rgb <= "111111";
					when "10100111011001010" => rgb <= "101010";
					when "10100111011001011" => rgb <= "111111";
					when "10100111011001100" => rgb <= "111111";
					when "10100111011001101" => rgb <= "101010";
					when "10100111011001110" => rgb <= "111111";
					when "10100111011001111" => rgb <= "010101";
					when "10100111011010000" => rgb <= "000000";
					when "10100111011010001" => rgb <= "000000";
					when "10100111011010010" => rgb <= "000000";
					when "10100111011010011" => rgb <= "000000";
					when "10100111011010100" => rgb <= "000000";
					when "10100111011010101" => rgb <= "000000";
					when "10100111011010110" => rgb <= "000000";
					when "10100111011010111" => rgb <= "101010";
					when "10100111011011000" => rgb <= "111111";
					when "10100111011011001" => rgb <= "101010";
					when "10100111011011010" => rgb <= "101010";
					when "10100111011011011" => rgb <= "111111";
					when "10100111011011100" => rgb <= "111111";
					when "10100111011011101" => rgb <= "111111";
					when "10100111011011110" => rgb <= "111111";
					when "10100111011011111" => rgb <= "111111";
					when "10100111011100000" => rgb <= "111111";
					when "10100111011100001" => rgb <= "101010";
					when "10100111011100010" => rgb <= "111111";
					when "10100111011100011" => rgb <= "101010";
					when "10100111011100100" => rgb <= "111111";
					when "10100111011100101" => rgb <= "111111";
					when "10100111011100110" => rgb <= "000000";
					when "10100111011100111" => rgb <= "000000";
					when "10100111011101000" => rgb <= "000000";
					when "10100111011101001" => rgb <= "000000";
					when "10100111011101010" => rgb <= "000000";
					when "10100111011101011" => rgb <= "000000";
					when "10100111011101100" => rgb <= "000000";
					when "10100111011101101" => rgb <= "010101";
					when "10100111011101110" => rgb <= "101010";
					when "10100111011101111" => rgb <= "101010";
					when "10100111011110000" => rgb <= "101010";
					when "10100111011110001" => rgb <= "111111";
					when "10100111011110010" => rgb <= "111111";
					when "10100111011110011" => rgb <= "111111";
					when "10100111011110100" => rgb <= "101010";
					when "10100111011110101" => rgb <= "000000";
					when "10100111011110110" => rgb <= "000000";
					when "10100111011110111" => rgb <= "000000";
					when "10100111011111000" => rgb <= "000000";
					when "10100111011111001" => rgb <= "000000";
					when "10100111011111010" => rgb <= "000000";
					when "10100111011111011" => rgb <= "000000";
					when "10100111011111100" => rgb <= "000000";
					when "10100111011111101" => rgb <= "000000";
					when "10100111011111110" => rgb <= "000000";
					when "10100111011111111" => rgb <= "000000";
					when "10100111100000000" => rgb <= "000000";
					when "10100111100000001" => rgb <= "000000";
					when "10100111100000010" => rgb <= "000000";
					when "10100111100000011" => rgb <= "000000";
					when "10100111100000100" => rgb <= "000000";
					when "10100111100000101" => rgb <= "000000";
					when "10100111100000110" => rgb <= "000000";
					when "10100111100000111" => rgb <= "000000";
					when "10100111100001000" => rgb <= "000000";
					when "10100111100001001" => rgb <= "000000";
					when "10100111100001010" => rgb <= "000000";
					when "10100111100001011" => rgb <= "010101";
					when "10100111100001100" => rgb <= "111111";
					when "10100111100001101" => rgb <= "101010";
					when "10100111100001110" => rgb <= "101010";
					when "10100111100001111" => rgb <= "101010";
					when "10100111100010000" => rgb <= "111111";
					when "10100111100010001" => rgb <= "111111";
					when "10100111100010010" => rgb <= "111111";
					when "10100111100010011" => rgb <= "111111";
					when "10100111100010100" => rgb <= "111111";
					when "10100111100010101" => rgb <= "111111";
					when "10100111100010110" => rgb <= "111111";
					when "10100111100010111" => rgb <= "111111";
					when "10100111100011000" => rgb <= "101010";
					when "10100111100011001" => rgb <= "111111";
					when "10100111100011010" => rgb <= "010101";
					when "10100111100011011" => rgb <= "000000";
					when "10100111100011100" => rgb <= "000000";
					when "10100111100011101" => rgb <= "000000";
					when "10100111100011110" => rgb <= "000000";
					when "10100111100011111" => rgb <= "000000";
					when "10100111100100000" => rgb <= "000000";
					when "10100111100100001" => rgb <= "000000";
					when "10100111100100010" => rgb <= "101010";
					when "10100111100100011" => rgb <= "111111";
					when "10100111100100100" => rgb <= "101010";
					when "10100111100100101" => rgb <= "101010";
					when "10100111100100110" => rgb <= "111111";
					when "10100111100100111" => rgb <= "111111";
					when "10100111100101000" => rgb <= "111111";
					when "10100111100101001" => rgb <= "111111";
					when "10100111100101010" => rgb <= "111111";
					when "10100111100101011" => rgb <= "111111";
					when "10100111100101100" => rgb <= "111111";
					when "10100111100101101" => rgb <= "111111";
					when "10100111100101110" => rgb <= "101010";
					when "10100111100101111" => rgb <= "101010";
					when "10100111100110000" => rgb <= "111111";
					when "10100111100110001" => rgb <= "000000";
					when "10100111100110010" => rgb <= "000000";
					when "10100111100110011" => rgb <= "000000";
					when "10100111100110100" => rgb <= "000000";
					when "10100111100110101" => rgb <= "000000";
					when "10100111100110110" => rgb <= "000000";
					when "10100111100110111" => rgb <= "000000";
					when "10100111100111000" => rgb <= "000000";
					when "10100111100111001" => rgb <= "000000";
					when "10100111100111010" => rgb <= "000000";
					when "10100111100111011" => rgb <= "000000";
					when "10100111100111100" => rgb <= "000000";
					when "10100111100111101" => rgb <= "000000";
					when "10100111100111110" => rgb <= "000000";
					when "10100111100111111" => rgb <= "000000";
					when "10101000000000000" => rgb <= "000000";
					when "10101000000000001" => rgb <= "000000";
					when "10101000000000010" => rgb <= "000000";
					when "10101000000000011" => rgb <= "000000";
					when "10101000000000100" => rgb <= "000000";
					when "10101000000000101" => rgb <= "101010";
					when "10101000000000110" => rgb <= "111111";
					when "10101000000000111" => rgb <= "101010";
					when "10101000000001000" => rgb <= "111111";
					when "10101000000001001" => rgb <= "111111";
					when "10101000000001010" => rgb <= "101010";
					when "10101000000001011" => rgb <= "101010";
					when "10101000000001100" => rgb <= "010101";
					when "10101000000001101" => rgb <= "000000";
					when "10101000000001110" => rgb <= "000000";
					when "10101000000001111" => rgb <= "000000";
					when "10101000000010000" => rgb <= "000000";
					when "10101000000010001" => rgb <= "000000";
					when "10101000000010010" => rgb <= "000000";
					when "10101000000010011" => rgb <= "000000";
					when "10101000000010100" => rgb <= "000000";
					when "10101000000010101" => rgb <= "000000";
					when "10101000000010110" => rgb <= "000000";
					when "10101000000010111" => rgb <= "000000";
					when "10101000000011000" => rgb <= "000000";
					when "10101000000011001" => rgb <= "000000";
					when "10101000000011010" => rgb <= "000000";
					when "10101000000011011" => rgb <= "000000";
					when "10101000000011100" => rgb <= "000000";
					when "10101000000011101" => rgb <= "000000";
					when "10101000000011110" => rgb <= "000000";
					when "10101000000011111" => rgb <= "000000";
					when "10101000000100000" => rgb <= "000000";
					when "10101000000100001" => rgb <= "000000";
					when "10101000000100010" => rgb <= "000000";
					when "10101000000100011" => rgb <= "101010";
					when "10101000000100100" => rgb <= "111111";
					when "10101000000100101" => rgb <= "101010";
					when "10101000000100110" => rgb <= "101010";
					when "10101000000100111" => rgb <= "111111";
					when "10101000000101000" => rgb <= "111111";
					when "10101000000101001" => rgb <= "111111";
					when "10101000000101010" => rgb <= "101010";
					when "10101000000101011" => rgb <= "111111";
					when "10101000000101100" => rgb <= "111111";
					when "10101000000101101" => rgb <= "111111";
					when "10101000000101110" => rgb <= "111111";
					when "10101000000101111" => rgb <= "101010";
					when "10101000000110000" => rgb <= "111111";
					when "10101000000110001" => rgb <= "101010";
					when "10101000000110010" => rgb <= "000000";
					when "10101000000110011" => rgb <= "000000";
					when "10101000000110100" => rgb <= "000000";
					when "10101000000110101" => rgb <= "000000";
					when "10101000000110110" => rgb <= "000000";
					when "10101000000110111" => rgb <= "000000";
					when "10101000000111000" => rgb <= "000000";
					when "10101000000111001" => rgb <= "000000";
					when "10101000000111010" => rgb <= "010101";
					when "10101000000111011" => rgb <= "010101";
					when "10101000000111100" => rgb <= "010101";
					when "10101000000111101" => rgb <= "010101";
					when "10101000000111110" => rgb <= "010101";
					when "10101000000111111" => rgb <= "010101";
					when "10101000001000000" => rgb <= "010101";
					when "10101000001000001" => rgb <= "010101";
					when "10101000001000010" => rgb <= "010101";
					when "10101000001000011" => rgb <= "010101";
					when "10101000001000100" => rgb <= "010101";
					when "10101000001000101" => rgb <= "010101";
					when "10101000001000110" => rgb <= "010101";
					when "10101000001000111" => rgb <= "010101";
					when "10101000001001000" => rgb <= "010101";
					when "10101000001001001" => rgb <= "010101";
					when "10101000001001010" => rgb <= "010101";
					when "10101000001001011" => rgb <= "010101";
					when "10101000001001100" => rgb <= "010101";
					when "10101000001001101" => rgb <= "010101";
					when "10101000001001110" => rgb <= "010101";
					when "10101000001001111" => rgb <= "010101";
					when "10101000001010000" => rgb <= "101010";
					when "10101000001010001" => rgb <= "111111";
					when "10101000001010010" => rgb <= "101010";
					when "10101000001010011" => rgb <= "111111";
					when "10101000001010100" => rgb <= "111111";
					when "10101000001010101" => rgb <= "111111";
					when "10101000001010110" => rgb <= "101010";
					when "10101000001010111" => rgb <= "101010";
					when "10101000001011000" => rgb <= "010101";
					when "10101000001011001" => rgb <= "010101";
					when "10101000001011010" => rgb <= "010101";
					when "10101000001011011" => rgb <= "010101";
					when "10101000001011100" => rgb <= "010101";
					when "10101000001011101" => rgb <= "010101";
					when "10101000001011110" => rgb <= "010101";
					when "10101000001011111" => rgb <= "000000";
					when "10101000001100000" => rgb <= "000000";
					when "10101000001100001" => rgb <= "000000";
					when "10101000001100010" => rgb <= "000000";
					when "10101000001100011" => rgb <= "000000";
					when "10101000001100100" => rgb <= "000000";
					when "10101000001100101" => rgb <= "000000";
					when "10101000001100110" => rgb <= "010101";
					when "10101000001100111" => rgb <= "111111";
					when "10101000001101000" => rgb <= "101010";
					when "10101000001101001" => rgb <= "111111";
					when "10101000001101010" => rgb <= "111111";
					when "10101000001101011" => rgb <= "111111";
					when "10101000001101100" => rgb <= "111111";
					when "10101000001101101" => rgb <= "101010";
					when "10101000001101110" => rgb <= "000000";
					when "10101000001101111" => rgb <= "000000";
					when "10101000001110000" => rgb <= "000000";
					when "10101000001110001" => rgb <= "000000";
					when "10101000001110010" => rgb <= "000000";
					when "10101000001110011" => rgb <= "000000";
					when "10101000001110100" => rgb <= "000000";
					when "10101000001110101" => rgb <= "000000";
					when "10101000001110110" => rgb <= "000000";
					when "10101000001110111" => rgb <= "000000";
					when "10101000001111000" => rgb <= "000000";
					when "10101000001111001" => rgb <= "000000";
					when "10101000001111010" => rgb <= "000000";
					when "10101000001111011" => rgb <= "000000";
					when "10101000001111100" => rgb <= "000000";
					when "10101000001111101" => rgb <= "101010";
					when "10101000001111110" => rgb <= "111111";
					when "10101000001111111" => rgb <= "111111";
					when "10101000010000000" => rgb <= "111111";
					when "10101000010000001" => rgb <= "111111";
					when "10101000010000010" => rgb <= "111111";
					when "10101000010000011" => rgb <= "111111";
					when "10101000010000100" => rgb <= "111111";
					when "10101000010000101" => rgb <= "111111";
					when "10101000010000110" => rgb <= "111111";
					when "10101000010000111" => rgb <= "111111";
					when "10101000010001000" => rgb <= "111111";
					when "10101000010001001" => rgb <= "111111";
					when "10101000010001010" => rgb <= "111111";
					when "10101000010001011" => rgb <= "101010";
					when "10101000010001100" => rgb <= "000000";
					when "10101000010001101" => rgb <= "000000";
					when "10101000010001110" => rgb <= "000000";
					when "10101000010001111" => rgb <= "000000";
					when "10101000010010000" => rgb <= "000000";
					when "10101000010010001" => rgb <= "000000";
					when "10101000010010010" => rgb <= "000000";
					when "10101000010010011" => rgb <= "000000";
					when "10101000010010100" => rgb <= "000000";
					when "10101000010010101" => rgb <= "000000";
					when "10101000010010110" => rgb <= "000000";
					when "10101000010010111" => rgb <= "000000";
					when "10101000010011000" => rgb <= "000000";
					when "10101000010011001" => rgb <= "000000";
					when "10101000010011010" => rgb <= "000000";
					when "10101000010011011" => rgb <= "000000";
					when "10101000010011100" => rgb <= "000000";
					when "10101000010011101" => rgb <= "000000";
					when "10101000010011110" => rgb <= "000000";
					when "10101000010011111" => rgb <= "000000";
					when "10101000010100000" => rgb <= "000000";
					when "10101000010100001" => rgb <= "000000";
					when "10101000010100010" => rgb <= "010101";
					when "10101000010100011" => rgb <= "111111";
					when "10101000010100100" => rgb <= "101010";
					when "10101000010100101" => rgb <= "111111";
					when "10101000010100110" => rgb <= "111111";
					when "10101000010100111" => rgb <= "111111";
					when "10101000010101000" => rgb <= "111111";
					when "10101000010101001" => rgb <= "101010";
					when "10101000010101010" => rgb <= "000000";
					when "10101000010101011" => rgb <= "000000";
					when "10101000010101100" => rgb <= "000000";
					when "10101000010101101" => rgb <= "000000";
					when "10101000010101110" => rgb <= "000000";
					when "10101000010101111" => rgb <= "000000";
					when "10101000010110000" => rgb <= "000000";
					when "10101000010110001" => rgb <= "000000";
					when "10101000010110010" => rgb <= "000000";
					when "10101000010110011" => rgb <= "000000";
					when "10101000010110100" => rgb <= "000000";
					when "10101000010110101" => rgb <= "000000";
					when "10101000010110110" => rgb <= "000000";
					when "10101000010110111" => rgb <= "000000";
					when "10101000010111000" => rgb <= "000000";
					when "10101000010111001" => rgb <= "000000";
					when "10101000010111010" => rgb <= "000000";
					when "10101000010111011" => rgb <= "000000";
					when "10101000010111100" => rgb <= "000000";
					when "10101000010111101" => rgb <= "000000";
					when "10101000010111110" => rgb <= "000000";
					when "10101000010111111" => rgb <= "000000";
					when "10101000011000000" => rgb <= "010101";
					when "10101000011000001" => rgb <= "101010";
					when "10101000011000010" => rgb <= "101010";
					when "10101000011000011" => rgb <= "111111";
					when "10101000011000100" => rgb <= "111111";
					when "10101000011000101" => rgb <= "111111";
					when "10101000011000110" => rgb <= "111111";
					when "10101000011000111" => rgb <= "111111";
					when "10101000011001000" => rgb <= "111111";
					when "10101000011001001" => rgb <= "101010";
					when "10101000011001010" => rgb <= "111111";
					when "10101000011001011" => rgb <= "101010";
					when "10101000011001100" => rgb <= "111111";
					when "10101000011001101" => rgb <= "101010";
					when "10101000011001110" => rgb <= "111111";
					when "10101000011001111" => rgb <= "010101";
					when "10101000011010000" => rgb <= "000000";
					when "10101000011010001" => rgb <= "000000";
					when "10101000011010010" => rgb <= "000000";
					when "10101000011010011" => rgb <= "000000";
					when "10101000011010100" => rgb <= "000000";
					when "10101000011010101" => rgb <= "000000";
					when "10101000011010110" => rgb <= "000000";
					when "10101000011010111" => rgb <= "101010";
					when "10101000011011000" => rgb <= "101010";
					when "10101000011011001" => rgb <= "101010";
					when "10101000011011010" => rgb <= "101010";
					when "10101000011011011" => rgb <= "111111";
					when "10101000011011100" => rgb <= "111111";
					when "10101000011011101" => rgb <= "111111";
					when "10101000011011110" => rgb <= "111111";
					when "10101000011011111" => rgb <= "111111";
					when "10101000011100000" => rgb <= "101010";
					when "10101000011100001" => rgb <= "111111";
					when "10101000011100010" => rgb <= "111111";
					when "10101000011100011" => rgb <= "101010";
					when "10101000011100100" => rgb <= "101010";
					when "10101000011100101" => rgb <= "101010";
					when "10101000011100110" => rgb <= "000000";
					when "10101000011100111" => rgb <= "000000";
					when "10101000011101000" => rgb <= "000000";
					when "10101000011101001" => rgb <= "000000";
					when "10101000011101010" => rgb <= "000000";
					when "10101000011101011" => rgb <= "000000";
					when "10101000011101100" => rgb <= "000000";
					when "10101000011101101" => rgb <= "010101";
					when "10101000011101110" => rgb <= "101010";
					when "10101000011101111" => rgb <= "101010";
					when "10101000011110000" => rgb <= "111111";
					when "10101000011110001" => rgb <= "101010";
					when "10101000011110010" => rgb <= "111111";
					when "10101000011110011" => rgb <= "101010";
					when "10101000011110100" => rgb <= "101010";
					when "10101000011110101" => rgb <= "101010";
					when "10101000011110110" => rgb <= "010101";
					when "10101000011110111" => rgb <= "010101";
					when "10101000011111000" => rgb <= "010101";
					when "10101000011111001" => rgb <= "010101";
					when "10101000011111010" => rgb <= "010101";
					when "10101000011111011" => rgb <= "010101";
					when "10101000011111100" => rgb <= "010101";
					when "10101000011111101" => rgb <= "000000";
					when "10101000011111110" => rgb <= "000000";
					when "10101000011111111" => rgb <= "000000";
					when "10101000100000000" => rgb <= "000000";
					when "10101000100000001" => rgb <= "000000";
					when "10101000100000010" => rgb <= "000000";
					when "10101000100000011" => rgb <= "000000";
					when "10101000100000100" => rgb <= "000000";
					when "10101000100000101" => rgb <= "000000";
					when "10101000100000110" => rgb <= "000000";
					when "10101000100000111" => rgb <= "000000";
					when "10101000100001000" => rgb <= "000000";
					when "10101000100001001" => rgb <= "000000";
					when "10101000100001010" => rgb <= "000000";
					when "10101000100001011" => rgb <= "010101";
					when "10101000100001100" => rgb <= "111111";
					when "10101000100001101" => rgb <= "101010";
					when "10101000100001110" => rgb <= "111111";
					when "10101000100001111" => rgb <= "111111";
					when "10101000100010000" => rgb <= "111111";
					when "10101000100010001" => rgb <= "111111";
					when "10101000100010010" => rgb <= "111111";
					when "10101000100010011" => rgb <= "111111";
					when "10101000100010100" => rgb <= "111111";
					when "10101000100010101" => rgb <= "111111";
					when "10101000100010110" => rgb <= "111111";
					when "10101000100010111" => rgb <= "111111";
					when "10101000100011000" => rgb <= "101010";
					when "10101000100011001" => rgb <= "101010";
					when "10101000100011010" => rgb <= "010101";
					when "10101000100011011" => rgb <= "000000";
					when "10101000100011100" => rgb <= "000000";
					when "10101000100011101" => rgb <= "000000";
					when "10101000100011110" => rgb <= "000000";
					when "10101000100011111" => rgb <= "000000";
					when "10101000100100000" => rgb <= "000000";
					when "10101000100100001" => rgb <= "000000";
					when "10101000100100010" => rgb <= "101010";
					when "10101000100100011" => rgb <= "101010";
					when "10101000100100100" => rgb <= "101010";
					when "10101000100100101" => rgb <= "111111";
					when "10101000100100110" => rgb <= "111111";
					when "10101000100100111" => rgb <= "111111";
					when "10101000100101000" => rgb <= "101010";
					when "10101000100101001" => rgb <= "111111";
					when "10101000100101010" => rgb <= "111111";
					when "10101000100101011" => rgb <= "101010";
					when "10101000100101100" => rgb <= "111111";
					when "10101000100101101" => rgb <= "111111";
					when "10101000100101110" => rgb <= "101010";
					when "10101000100101111" => rgb <= "101010";
					when "10101000100110000" => rgb <= "101010";
					when "10101000100110001" => rgb <= "000000";
					when "10101000100110010" => rgb <= "000000";
					when "10101000100110011" => rgb <= "000000";
					when "10101000100110100" => rgb <= "000000";
					when "10101000100110101" => rgb <= "000000";
					when "10101000100110110" => rgb <= "000000";
					when "10101000100110111" => rgb <= "000000";
					when "10101000100111000" => rgb <= "000000";
					when "10101000100111001" => rgb <= "000000";
					when "10101000100111010" => rgb <= "000000";
					when "10101000100111011" => rgb <= "000000";
					when "10101000100111100" => rgb <= "000000";
					when "10101000100111101" => rgb <= "000000";
					when "10101000100111110" => rgb <= "000000";
					when "10101000100111111" => rgb <= "000000";
					when "10101001000000000" => rgb <= "000000";
					when "10101001000000001" => rgb <= "000000";
					when "10101001000000010" => rgb <= "000000";
					when "10101001000000011" => rgb <= "000000";
					when "10101001000000100" => rgb <= "000000";
					when "10101001000000101" => rgb <= "101010";
					when "10101001000000110" => rgb <= "111111";
					when "10101001000000111" => rgb <= "101010";
					when "10101001000001000" => rgb <= "111111";
					when "10101001000001001" => rgb <= "111111";
					when "10101001000001010" => rgb <= "101010";
					when "10101001000001011" => rgb <= "111111";
					when "10101001000001100" => rgb <= "101010";
					when "10101001000001101" => rgb <= "000000";
					when "10101001000001110" => rgb <= "000000";
					when "10101001000001111" => rgb <= "000000";
					when "10101001000010000" => rgb <= "000000";
					when "10101001000010001" => rgb <= "000000";
					when "10101001000010010" => rgb <= "000000";
					when "10101001000010011" => rgb <= "000000";
					when "10101001000010100" => rgb <= "000000";
					when "10101001000010101" => rgb <= "000000";
					when "10101001000010110" => rgb <= "000000";
					when "10101001000010111" => rgb <= "000000";
					when "10101001000011000" => rgb <= "000000";
					when "10101001000011001" => rgb <= "000000";
					when "10101001000011010" => rgb <= "000000";
					when "10101001000011011" => rgb <= "000000";
					when "10101001000011100" => rgb <= "000000";
					when "10101001000011101" => rgb <= "000000";
					when "10101001000011110" => rgb <= "000000";
					when "10101001000011111" => rgb <= "000000";
					when "10101001000100000" => rgb <= "000000";
					when "10101001000100001" => rgb <= "000000";
					when "10101001000100010" => rgb <= "000000";
					when "10101001000100011" => rgb <= "101010";
					when "10101001000100100" => rgb <= "111111";
					when "10101001000100101" => rgb <= "111111";
					when "10101001000100110" => rgb <= "111111";
					when "10101001000100111" => rgb <= "111111";
					when "10101001000101000" => rgb <= "111111";
					when "10101001000101001" => rgb <= "111111";
					when "10101001000101010" => rgb <= "101010";
					when "10101001000101011" => rgb <= "111111";
					when "10101001000101100" => rgb <= "111111";
					when "10101001000101101" => rgb <= "111111";
					when "10101001000101110" => rgb <= "111111";
					when "10101001000101111" => rgb <= "101010";
					when "10101001000110000" => rgb <= "111111";
					when "10101001000110001" => rgb <= "101010";
					when "10101001000110010" => rgb <= "000000";
					when "10101001000110011" => rgb <= "000000";
					when "10101001000110100" => rgb <= "000000";
					when "10101001000110101" => rgb <= "000000";
					when "10101001000110110" => rgb <= "000000";
					when "10101001000110111" => rgb <= "000000";
					when "10101001000111000" => rgb <= "000000";
					when "10101001000111001" => rgb <= "010101";
					when "10101001000111010" => rgb <= "101010";
					when "10101001000111011" => rgb <= "101010";
					when "10101001000111100" => rgb <= "111111";
					when "10101001000111101" => rgb <= "101010";
					when "10101001000111110" => rgb <= "111111";
					when "10101001000111111" => rgb <= "111111";
					when "10101001001000000" => rgb <= "101010";
					when "10101001001000001" => rgb <= "000000";
					when "10101001001000010" => rgb <= "000000";
					when "10101001001000011" => rgb <= "000000";
					when "10101001001000100" => rgb <= "000000";
					when "10101001001000101" => rgb <= "000000";
					when "10101001001000110" => rgb <= "000000";
					when "10101001001000111" => rgb <= "000000";
					when "10101001001001000" => rgb <= "000000";
					when "10101001001001001" => rgb <= "000000";
					when "10101001001001010" => rgb <= "000000";
					when "10101001001001011" => rgb <= "000000";
					when "10101001001001100" => rgb <= "000000";
					when "10101001001001101" => rgb <= "000000";
					when "10101001001001110" => rgb <= "000000";
					when "10101001001001111" => rgb <= "000000";
					when "10101001001010000" => rgb <= "101010";
					when "10101001001010001" => rgb <= "101010";
					when "10101001001010010" => rgb <= "101010";
					when "10101001001010011" => rgb <= "111111";
					when "10101001001010100" => rgb <= "101010";
					when "10101001001010101" => rgb <= "111111";
					when "10101001001010110" => rgb <= "101010";
					when "10101001001010111" => rgb <= "101010";
					when "10101001001011000" => rgb <= "111111";
					when "10101001001011001" => rgb <= "111111";
					when "10101001001011010" => rgb <= "111111";
					when "10101001001011011" => rgb <= "101010";
					when "10101001001011100" => rgb <= "111111";
					when "10101001001011101" => rgb <= "111111";
					when "10101001001011110" => rgb <= "101010";
					when "10101001001011111" => rgb <= "000000";
					when "10101001001100000" => rgb <= "000000";
					when "10101001001100001" => rgb <= "000000";
					when "10101001001100010" => rgb <= "000000";
					when "10101001001100011" => rgb <= "000000";
					when "10101001001100100" => rgb <= "000000";
					when "10101001001100101" => rgb <= "000000";
					when "10101001001100110" => rgb <= "010101";
					when "10101001001100111" => rgb <= "111111";
					when "10101001001101000" => rgb <= "101010";
					when "10101001001101001" => rgb <= "111111";
					when "10101001001101010" => rgb <= "101010";
					when "10101001001101011" => rgb <= "101010";
					when "10101001001101100" => rgb <= "111111";
					when "10101001001101101" => rgb <= "111111";
					when "10101001001101110" => rgb <= "000000";
					when "10101001001101111" => rgb <= "000000";
					when "10101001001110000" => rgb <= "000000";
					when "10101001001110001" => rgb <= "000000";
					when "10101001001110010" => rgb <= "000000";
					when "10101001001110011" => rgb <= "000000";
					when "10101001001110100" => rgb <= "000000";
					when "10101001001110101" => rgb <= "000000";
					when "10101001001110110" => rgb <= "000000";
					when "10101001001110111" => rgb <= "000000";
					when "10101001001111000" => rgb <= "000000";
					when "10101001001111001" => rgb <= "000000";
					when "10101001001111010" => rgb <= "000000";
					when "10101001001111011" => rgb <= "000000";
					when "10101001001111100" => rgb <= "000000";
					when "10101001001111101" => rgb <= "101010";
					when "10101001001111110" => rgb <= "111111";
					when "10101001001111111" => rgb <= "111111";
					when "10101001010000000" => rgb <= "111111";
					when "10101001010000001" => rgb <= "111111";
					when "10101001010000010" => rgb <= "111111";
					when "10101001010000011" => rgb <= "111111";
					when "10101001010000100" => rgb <= "111111";
					when "10101001010000101" => rgb <= "111111";
					when "10101001010000110" => rgb <= "111111";
					when "10101001010000111" => rgb <= "111111";
					when "10101001010001000" => rgb <= "111111";
					when "10101001010001001" => rgb <= "111111";
					when "10101001010001010" => rgb <= "111111";
					when "10101001010001011" => rgb <= "101010";
					when "10101001010001100" => rgb <= "000000";
					when "10101001010001101" => rgb <= "000000";
					when "10101001010001110" => rgb <= "000000";
					when "10101001010001111" => rgb <= "000000";
					when "10101001010010000" => rgb <= "000000";
					when "10101001010010001" => rgb <= "000000";
					when "10101001010010010" => rgb <= "000000";
					when "10101001010010011" => rgb <= "000000";
					when "10101001010010100" => rgb <= "000000";
					when "10101001010010101" => rgb <= "000000";
					when "10101001010010110" => rgb <= "000000";
					when "10101001010010111" => rgb <= "000000";
					when "10101001010011000" => rgb <= "000000";
					when "10101001010011001" => rgb <= "000000";
					when "10101001010011010" => rgb <= "000000";
					when "10101001010011011" => rgb <= "000000";
					when "10101001010011100" => rgb <= "000000";
					when "10101001010011101" => rgb <= "000000";
					when "10101001010011110" => rgb <= "000000";
					when "10101001010011111" => rgb <= "000000";
					when "10101001010100000" => rgb <= "000000";
					when "10101001010100001" => rgb <= "000000";
					when "10101001010100010" => rgb <= "010101";
					when "10101001010100011" => rgb <= "111111";
					when "10101001010100100" => rgb <= "101010";
					when "10101001010100101" => rgb <= "111111";
					when "10101001010100110" => rgb <= "111111";
					when "10101001010100111" => rgb <= "111111";
					when "10101001010101000" => rgb <= "111111";
					when "10101001010101001" => rgb <= "111111";
					when "10101001010101010" => rgb <= "000000";
					when "10101001010101011" => rgb <= "000000";
					when "10101001010101100" => rgb <= "000000";
					when "10101001010101101" => rgb <= "000000";
					when "10101001010101110" => rgb <= "000000";
					when "10101001010101111" => rgb <= "000000";
					when "10101001010110000" => rgb <= "000000";
					when "10101001010110001" => rgb <= "000000";
					when "10101001010110010" => rgb <= "000000";
					when "10101001010110011" => rgb <= "000000";
					when "10101001010110100" => rgb <= "000000";
					when "10101001010110101" => rgb <= "000000";
					when "10101001010110110" => rgb <= "000000";
					when "10101001010110111" => rgb <= "000000";
					when "10101001010111000" => rgb <= "000000";
					when "10101001010111001" => rgb <= "000000";
					when "10101001010111010" => rgb <= "000000";
					when "10101001010111011" => rgb <= "000000";
					when "10101001010111100" => rgb <= "000000";
					when "10101001010111101" => rgb <= "000000";
					when "10101001010111110" => rgb <= "000000";
					when "10101001010111111" => rgb <= "000000";
					when "10101001011000000" => rgb <= "010101";
					when "10101001011000001" => rgb <= "101010";
					when "10101001011000010" => rgb <= "101010";
					when "10101001011000011" => rgb <= "111111";
					when "10101001011000100" => rgb <= "111111";
					when "10101001011000101" => rgb <= "111111";
					when "10101001011000110" => rgb <= "111111";
					when "10101001011000111" => rgb <= "111111";
					when "10101001011001000" => rgb <= "111111";
					when "10101001011001001" => rgb <= "101010";
					when "10101001011001010" => rgb <= "111111";
					when "10101001011001011" => rgb <= "101010";
					when "10101001011001100" => rgb <= "111111";
					when "10101001011001101" => rgb <= "101010";
					when "10101001011001110" => rgb <= "111111";
					when "10101001011001111" => rgb <= "010101";
					when "10101001011010000" => rgb <= "000000";
					when "10101001011010001" => rgb <= "000000";
					when "10101001011010010" => rgb <= "000000";
					when "10101001011010011" => rgb <= "000000";
					when "10101001011010100" => rgb <= "000000";
					when "10101001011010101" => rgb <= "000000";
					when "10101001011010110" => rgb <= "000000";
					when "10101001011010111" => rgb <= "101010";
					when "10101001011011000" => rgb <= "101010";
					when "10101001011011001" => rgb <= "101010";
					when "10101001011011010" => rgb <= "101010";
					when "10101001011011011" => rgb <= "111111";
					when "10101001011011100" => rgb <= "111111";
					when "10101001011011101" => rgb <= "111111";
					when "10101001011011110" => rgb <= "111111";
					when "10101001011011111" => rgb <= "111111";
					when "10101001011100000" => rgb <= "111111";
					when "10101001011100001" => rgb <= "111111";
					when "10101001011100010" => rgb <= "111111";
					when "10101001011100011" => rgb <= "111111";
					when "10101001011100100" => rgb <= "111111";
					when "10101001011100101" => rgb <= "111111";
					when "10101001011100110" => rgb <= "000000";
					when "10101001011100111" => rgb <= "000000";
					when "10101001011101000" => rgb <= "000000";
					when "10101001011101001" => rgb <= "000000";
					when "10101001011101010" => rgb <= "000000";
					when "10101001011101011" => rgb <= "000000";
					when "10101001011101100" => rgb <= "000000";
					when "10101001011101101" => rgb <= "010101";
					when "10101001011101110" => rgb <= "111111";
					when "10101001011101111" => rgb <= "101010";
					when "10101001011110000" => rgb <= "101010";
					when "10101001011110001" => rgb <= "101010";
					when "10101001011110010" => rgb <= "111111";
					when "10101001011110011" => rgb <= "101010";
					when "10101001011110100" => rgb <= "111111";
					when "10101001011110101" => rgb <= "101010";
					when "10101001011110110" => rgb <= "111111";
					when "10101001011110111" => rgb <= "111111";
					when "10101001011111000" => rgb <= "111111";
					when "10101001011111001" => rgb <= "111111";
					when "10101001011111010" => rgb <= "111111";
					when "10101001011111011" => rgb <= "111111";
					when "10101001011111100" => rgb <= "010101";
					when "10101001011111101" => rgb <= "000000";
					when "10101001011111110" => rgb <= "000000";
					when "10101001011111111" => rgb <= "000000";
					when "10101001100000000" => rgb <= "000000";
					when "10101001100000001" => rgb <= "000000";
					when "10101001100000010" => rgb <= "000000";
					when "10101001100000011" => rgb <= "000000";
					when "10101001100000100" => rgb <= "000000";
					when "10101001100000101" => rgb <= "000000";
					when "10101001100000110" => rgb <= "000000";
					when "10101001100000111" => rgb <= "000000";
					when "10101001100001000" => rgb <= "000000";
					when "10101001100001001" => rgb <= "000000";
					when "10101001100001010" => rgb <= "000000";
					when "10101001100001011" => rgb <= "010101";
					when "10101001100001100" => rgb <= "111111";
					when "10101001100001101" => rgb <= "101010";
					when "10101001100001110" => rgb <= "111111";
					when "10101001100001111" => rgb <= "111111";
					when "10101001100010000" => rgb <= "111111";
					when "10101001100010001" => rgb <= "111111";
					when "10101001100010010" => rgb <= "111111";
					when "10101001100010011" => rgb <= "111111";
					when "10101001100010100" => rgb <= "111111";
					when "10101001100010101" => rgb <= "111111";
					when "10101001100010110" => rgb <= "111111";
					when "10101001100010111" => rgb <= "111111";
					when "10101001100011000" => rgb <= "111111";
					when "10101001100011001" => rgb <= "111111";
					when "10101001100011010" => rgb <= "101010";
					when "10101001100011011" => rgb <= "000000";
					when "10101001100011100" => rgb <= "000000";
					when "10101001100011101" => rgb <= "000000";
					when "10101001100011110" => rgb <= "000000";
					when "10101001100011111" => rgb <= "000000";
					when "10101001100100000" => rgb <= "000000";
					when "10101001100100001" => rgb <= "000000";
					when "10101001100100010" => rgb <= "101010";
					when "10101001100100011" => rgb <= "111111";
					when "10101001100100100" => rgb <= "101010";
					when "10101001100100101" => rgb <= "111111";
					when "10101001100100110" => rgb <= "111111";
					when "10101001100100111" => rgb <= "111111";
					when "10101001100101000" => rgb <= "101010";
					when "10101001100101001" => rgb <= "111111";
					when "10101001100101010" => rgb <= "111111";
					when "10101001100101011" => rgb <= "101010";
					when "10101001100101100" => rgb <= "111111";
					when "10101001100101101" => rgb <= "111111";
					when "10101001100101110" => rgb <= "101010";
					when "10101001100101111" => rgb <= "101010";
					when "10101001100110000" => rgb <= "111111";
					when "10101001100110001" => rgb <= "010101";
					when "10101001100110010" => rgb <= "000000";
					when "10101001100110011" => rgb <= "000000";
					when "10101001100110100" => rgb <= "000000";
					when "10101001100110101" => rgb <= "000000";
					when "10101001100110110" => rgb <= "000000";
					when "10101001100110111" => rgb <= "000000";
					when "10101001100111000" => rgb <= "000000";
					when "10101001100111001" => rgb <= "000000";
					when "10101001100111010" => rgb <= "000000";
					when "10101001100111011" => rgb <= "000000";
					when "10101001100111100" => rgb <= "000000";
					when "10101001100111101" => rgb <= "000000";
					when "10101001100111110" => rgb <= "000000";
					when "10101001100111111" => rgb <= "000000";
					when "10101010000000000" => rgb <= "000000";
					when "10101010000000001" => rgb <= "000000";
					when "10101010000000010" => rgb <= "000000";
					when "10101010000000011" => rgb <= "000000";
					when "10101010000000100" => rgb <= "000000";
					when "10101010000000101" => rgb <= "101010";
					when "10101010000000110" => rgb <= "111111";
					when "10101010000000111" => rgb <= "101010";
					when "10101010000001000" => rgb <= "111111";
					when "10101010000001001" => rgb <= "111111";
					when "10101010000001010" => rgb <= "101010";
					when "10101010000001011" => rgb <= "111111";
					when "10101010000001100" => rgb <= "101010";
					when "10101010000001101" => rgb <= "000000";
					when "10101010000001110" => rgb <= "000000";
					when "10101010000001111" => rgb <= "000000";
					when "10101010000010000" => rgb <= "000000";
					when "10101010000010001" => rgb <= "000000";
					when "10101010000010010" => rgb <= "000000";
					when "10101010000010011" => rgb <= "000000";
					when "10101010000010100" => rgb <= "000000";
					when "10101010000010101" => rgb <= "000000";
					when "10101010000010110" => rgb <= "000000";
					when "10101010000010111" => rgb <= "000000";
					when "10101010000011000" => rgb <= "000000";
					when "10101010000011001" => rgb <= "000000";
					when "10101010000011010" => rgb <= "000000";
					when "10101010000011011" => rgb <= "000000";
					when "10101010000011100" => rgb <= "000000";
					when "10101010000011101" => rgb <= "000000";
					when "10101010000011110" => rgb <= "000000";
					when "10101010000011111" => rgb <= "000000";
					when "10101010000100000" => rgb <= "000000";
					when "10101010000100001" => rgb <= "000000";
					when "10101010000100010" => rgb <= "000000";
					when "10101010000100011" => rgb <= "101010";
					when "10101010000100100" => rgb <= "111111";
					when "10101010000100101" => rgb <= "111111";
					when "10101010000100110" => rgb <= "111111";
					when "10101010000100111" => rgb <= "111111";
					when "10101010000101000" => rgb <= "111111";
					when "10101010000101001" => rgb <= "111111";
					when "10101010000101010" => rgb <= "101010";
					when "10101010000101011" => rgb <= "111111";
					when "10101010000101100" => rgb <= "111111";
					when "10101010000101101" => rgb <= "111111";
					when "10101010000101110" => rgb <= "111111";
					when "10101010000101111" => rgb <= "101010";
					when "10101010000110000" => rgb <= "101010";
					when "10101010000110001" => rgb <= "101010";
					when "10101010000110010" => rgb <= "000000";
					when "10101010000110011" => rgb <= "000000";
					when "10101010000110100" => rgb <= "000000";
					when "10101010000110101" => rgb <= "000000";
					when "10101010000110110" => rgb <= "000000";
					when "10101010000110111" => rgb <= "000000";
					when "10101010000111000" => rgb <= "000000";
					when "10101010000111001" => rgb <= "010101";
					when "10101010000111010" => rgb <= "101010";
					when "10101010000111011" => rgb <= "101010";
					when "10101010000111100" => rgb <= "101010";
					when "10101010000111101" => rgb <= "101010";
					when "10101010000111110" => rgb <= "101010";
					when "10101010000111111" => rgb <= "111111";
					when "10101010001000000" => rgb <= "101010";
					when "10101010001000001" => rgb <= "000000";
					when "10101010001000010" => rgb <= "000000";
					when "10101010001000011" => rgb <= "000000";
					when "10101010001000100" => rgb <= "000000";
					when "10101010001000101" => rgb <= "000000";
					when "10101010001000110" => rgb <= "000000";
					when "10101010001000111" => rgb <= "000000";
					when "10101010001001000" => rgb <= "000000";
					when "10101010001001001" => rgb <= "000000";
					when "10101010001001010" => rgb <= "000000";
					when "10101010001001011" => rgb <= "000000";
					when "10101010001001100" => rgb <= "000000";
					when "10101010001001101" => rgb <= "000000";
					when "10101010001001110" => rgb <= "000000";
					when "10101010001001111" => rgb <= "000000";
					when "10101010001010000" => rgb <= "101010";
					when "10101010001010001" => rgb <= "101010";
					when "10101010001010010" => rgb <= "111111";
					when "10101010001010011" => rgb <= "111111";
					when "10101010001010100" => rgb <= "101010";
					when "10101010001010101" => rgb <= "111111";
					when "10101010001010110" => rgb <= "111111";
					when "10101010001010111" => rgb <= "111111";
					when "10101010001011000" => rgb <= "101010";
					when "10101010001011001" => rgb <= "101010";
					when "10101010001011010" => rgb <= "101010";
					when "10101010001011011" => rgb <= "101010";
					when "10101010001011100" => rgb <= "101010";
					when "10101010001011101" => rgb <= "111111";
					when "10101010001011110" => rgb <= "101010";
					when "10101010001011111" => rgb <= "000000";
					when "10101010001100000" => rgb <= "000000";
					when "10101010001100001" => rgb <= "000000";
					when "10101010001100010" => rgb <= "000000";
					when "10101010001100011" => rgb <= "000000";
					when "10101010001100100" => rgb <= "000000";
					when "10101010001100101" => rgb <= "000000";
					when "10101010001100110" => rgb <= "010101";
					when "10101010001100111" => rgb <= "111111";
					when "10101010001101000" => rgb <= "101010";
					when "10101010001101001" => rgb <= "111111";
					when "10101010001101010" => rgb <= "101010";
					when "10101010001101011" => rgb <= "101010";
					when "10101010001101100" => rgb <= "101010";
					when "10101010001101101" => rgb <= "111111";
					when "10101010001101110" => rgb <= "000000";
					when "10101010001101111" => rgb <= "000000";
					when "10101010001110000" => rgb <= "000000";
					when "10101010001110001" => rgb <= "000000";
					when "10101010001110010" => rgb <= "000000";
					when "10101010001110011" => rgb <= "000000";
					when "10101010001110100" => rgb <= "000000";
					when "10101010001110101" => rgb <= "000000";
					when "10101010001110110" => rgb <= "000000";
					when "10101010001110111" => rgb <= "000000";
					when "10101010001111000" => rgb <= "000000";
					when "10101010001111001" => rgb <= "000000";
					when "10101010001111010" => rgb <= "000000";
					when "10101010001111011" => rgb <= "000000";
					when "10101010001111100" => rgb <= "000000";
					when "10101010001111101" => rgb <= "101010";
					when "10101010001111110" => rgb <= "111111";
					when "10101010001111111" => rgb <= "111111";
					when "10101010010000000" => rgb <= "111111";
					when "10101010010000001" => rgb <= "111111";
					when "10101010010000010" => rgb <= "111111";
					when "10101010010000011" => rgb <= "111111";
					when "10101010010000100" => rgb <= "111111";
					when "10101010010000101" => rgb <= "111111";
					when "10101010010000110" => rgb <= "111111";
					when "10101010010000111" => rgb <= "111111";
					when "10101010010001000" => rgb <= "111111";
					when "10101010010001001" => rgb <= "111111";
					when "10101010010001010" => rgb <= "111111";
					when "10101010010001011" => rgb <= "101010";
					when "10101010010001100" => rgb <= "000000";
					when "10101010010001101" => rgb <= "000000";
					when "10101010010001110" => rgb <= "000000";
					when "10101010010001111" => rgb <= "000000";
					when "10101010010010000" => rgb <= "000000";
					when "10101010010010001" => rgb <= "000000";
					when "10101010010010010" => rgb <= "000000";
					when "10101010010010011" => rgb <= "000000";
					when "10101010010010100" => rgb <= "000000";
					when "10101010010010101" => rgb <= "000000";
					when "10101010010010110" => rgb <= "000000";
					when "10101010010010111" => rgb <= "000000";
					when "10101010010011000" => rgb <= "000000";
					when "10101010010011001" => rgb <= "000000";
					when "10101010010011010" => rgb <= "000000";
					when "10101010010011011" => rgb <= "000000";
					when "10101010010011100" => rgb <= "000000";
					when "10101010010011101" => rgb <= "000000";
					when "10101010010011110" => rgb <= "000000";
					when "10101010010011111" => rgb <= "000000";
					when "10101010010100000" => rgb <= "000000";
					when "10101010010100001" => rgb <= "000000";
					when "10101010010100010" => rgb <= "010101";
					when "10101010010100011" => rgb <= "111111";
					when "10101010010100100" => rgb <= "101010";
					when "10101010010100101" => rgb <= "111111";
					when "10101010010100110" => rgb <= "111111";
					when "10101010010100111" => rgb <= "111111";
					when "10101010010101000" => rgb <= "101010";
					when "10101010010101001" => rgb <= "101010";
					when "10101010010101010" => rgb <= "000000";
					when "10101010010101011" => rgb <= "000000";
					when "10101010010101100" => rgb <= "000000";
					when "10101010010101101" => rgb <= "000000";
					when "10101010010101110" => rgb <= "000000";
					when "10101010010101111" => rgb <= "000000";
					when "10101010010110000" => rgb <= "000000";
					when "10101010010110001" => rgb <= "000000";
					when "10101010010110010" => rgb <= "000000";
					when "10101010010110011" => rgb <= "000000";
					when "10101010010110100" => rgb <= "000000";
					when "10101010010110101" => rgb <= "000000";
					when "10101010010110110" => rgb <= "000000";
					when "10101010010110111" => rgb <= "000000";
					when "10101010010111000" => rgb <= "000000";
					when "10101010010111001" => rgb <= "000000";
					when "10101010010111010" => rgb <= "000000";
					when "10101010010111011" => rgb <= "000000";
					when "10101010010111100" => rgb <= "000000";
					when "10101010010111101" => rgb <= "000000";
					when "10101010010111110" => rgb <= "000000";
					when "10101010010111111" => rgb <= "000000";
					when "10101010011000000" => rgb <= "010101";
					when "10101010011000001" => rgb <= "101010";
					when "10101010011000010" => rgb <= "101010";
					when "10101010011000011" => rgb <= "111111";
					when "10101010011000100" => rgb <= "111111";
					when "10101010011000101" => rgb <= "111111";
					when "10101010011000110" => rgb <= "111111";
					when "10101010011000111" => rgb <= "111111";
					when "10101010011001000" => rgb <= "111111";
					when "10101010011001001" => rgb <= "101010";
					when "10101010011001010" => rgb <= "111111";
					when "10101010011001011" => rgb <= "101010";
					when "10101010011001100" => rgb <= "111111";
					when "10101010011001101" => rgb <= "101010";
					when "10101010011001110" => rgb <= "111111";
					when "10101010011001111" => rgb <= "010101";
					when "10101010011010000" => rgb <= "000000";
					when "10101010011010001" => rgb <= "000000";
					when "10101010011010010" => rgb <= "000000";
					when "10101010011010011" => rgb <= "000000";
					when "10101010011010100" => rgb <= "000000";
					when "10101010011010101" => rgb <= "000000";
					when "10101010011010110" => rgb <= "000000";
					when "10101010011010111" => rgb <= "101010";
					when "10101010011011000" => rgb <= "101010";
					when "10101010011011001" => rgb <= "101010";
					when "10101010011011010" => rgb <= "101010";
					when "10101010011011011" => rgb <= "111111";
					when "10101010011011100" => rgb <= "111111";
					when "10101010011011101" => rgb <= "111111";
					when "10101010011011110" => rgb <= "111111";
					when "10101010011011111" => rgb <= "111111";
					when "10101010011100000" => rgb <= "111111";
					when "10101010011100001" => rgb <= "111111";
					when "10101010011100010" => rgb <= "101010";
					when "10101010011100011" => rgb <= "101010";
					when "10101010011100100" => rgb <= "111111";
					when "10101010011100101" => rgb <= "111111";
					when "10101010011100110" => rgb <= "000000";
					when "10101010011100111" => rgb <= "000000";
					when "10101010011101000" => rgb <= "000000";
					when "10101010011101001" => rgb <= "000000";
					when "10101010011101010" => rgb <= "000000";
					when "10101010011101011" => rgb <= "000000";
					when "10101010011101100" => rgb <= "000000";
					when "10101010011101101" => rgb <= "010101";
					when "10101010011101110" => rgb <= "111111";
					when "10101010011101111" => rgb <= "101010";
					when "10101010011110000" => rgb <= "111111";
					when "10101010011110001" => rgb <= "111111";
					when "10101010011110010" => rgb <= "111111";
					when "10101010011110011" => rgb <= "101010";
					when "10101010011110100" => rgb <= "101010";
					when "10101010011110101" => rgb <= "101010";
					when "10101010011110110" => rgb <= "101010";
					when "10101010011110111" => rgb <= "101010";
					when "10101010011111000" => rgb <= "101010";
					when "10101010011111001" => rgb <= "101010";
					when "10101010011111010" => rgb <= "101010";
					when "10101010011111011" => rgb <= "111111";
					when "10101010011111100" => rgb <= "010101";
					when "10101010011111101" => rgb <= "000000";
					when "10101010011111110" => rgb <= "000000";
					when "10101010011111111" => rgb <= "000000";
					when "10101010100000000" => rgb <= "000000";
					when "10101010100000001" => rgb <= "000000";
					when "10101010100000010" => rgb <= "000000";
					when "10101010100000011" => rgb <= "000000";
					when "10101010100000100" => rgb <= "000000";
					when "10101010100000101" => rgb <= "000000";
					when "10101010100000110" => rgb <= "000000";
					when "10101010100000111" => rgb <= "000000";
					when "10101010100001000" => rgb <= "000000";
					when "10101010100001001" => rgb <= "000000";
					when "10101010100001010" => rgb <= "000000";
					when "10101010100001011" => rgb <= "010101";
					when "10101010100001100" => rgb <= "111111";
					when "10101010100001101" => rgb <= "101010";
					when "10101010100001110" => rgb <= "111111";
					when "10101010100001111" => rgb <= "111111";
					when "10101010100010000" => rgb <= "111111";
					when "10101010100010001" => rgb <= "111111";
					when "10101010100010010" => rgb <= "111111";
					when "10101010100010011" => rgb <= "111111";
					when "10101010100010100" => rgb <= "111111";
					when "10101010100010101" => rgb <= "111111";
					when "10101010100010110" => rgb <= "111111";
					when "10101010100010111" => rgb <= "111111";
					when "10101010100011000" => rgb <= "101010";
					when "10101010100011001" => rgb <= "101010";
					when "10101010100011010" => rgb <= "101010";
					when "10101010100011011" => rgb <= "000000";
					when "10101010100011100" => rgb <= "000000";
					when "10101010100011101" => rgb <= "000000";
					when "10101010100011110" => rgb <= "000000";
					when "10101010100011111" => rgb <= "000000";
					when "10101010100100000" => rgb <= "000000";
					when "10101010100100001" => rgb <= "000000";
					when "10101010100100010" => rgb <= "101010";
					when "10101010100100011" => rgb <= "101010";
					when "10101010100100100" => rgb <= "101010";
					when "10101010100100101" => rgb <= "101010";
					when "10101010100100110" => rgb <= "111111";
					when "10101010100100111" => rgb <= "111111";
					when "10101010100101000" => rgb <= "101010";
					when "10101010100101001" => rgb <= "111111";
					when "10101010100101010" => rgb <= "111111";
					when "10101010100101011" => rgb <= "101010";
					when "10101010100101100" => rgb <= "111111";
					when "10101010100101101" => rgb <= "111111";
					when "10101010100101110" => rgb <= "101010";
					when "10101010100101111" => rgb <= "101010";
					when "10101010100110000" => rgb <= "111111";
					when "10101010100110001" => rgb <= "010101";
					when "10101010100110010" => rgb <= "000000";
					when "10101010100110011" => rgb <= "000000";
					when "10101010100110100" => rgb <= "000000";
					when "10101010100110101" => rgb <= "000000";
					when "10101010100110110" => rgb <= "000000";
					when "10101010100110111" => rgb <= "000000";
					when "10101010100111000" => rgb <= "000000";
					when "10101010100111001" => rgb <= "000000";
					when "10101010100111010" => rgb <= "000000";
					when "10101010100111011" => rgb <= "000000";
					when "10101010100111100" => rgb <= "000000";
					when "10101010100111101" => rgb <= "000000";
					when "10101010100111110" => rgb <= "000000";
					when "10101010100111111" => rgb <= "000000";
					when "10101011000000000" => rgb <= "000000";
					when "10101011000000001" => rgb <= "000000";
					when "10101011000000010" => rgb <= "000000";
					when "10101011000000011" => rgb <= "000000";
					when "10101011000000100" => rgb <= "000000";
					when "10101011000000101" => rgb <= "101010";
					when "10101011000000110" => rgb <= "111111";
					when "10101011000000111" => rgb <= "101010";
					when "10101011000001000" => rgb <= "111111";
					when "10101011000001001" => rgb <= "111111";
					when "10101011000001010" => rgb <= "101010";
					when "10101011000001011" => rgb <= "101010";
					when "10101011000001100" => rgb <= "101010";
					when "10101011000001101" => rgb <= "000000";
					when "10101011000001110" => rgb <= "000000";
					when "10101011000001111" => rgb <= "000000";
					when "10101011000010000" => rgb <= "000000";
					when "10101011000010001" => rgb <= "000000";
					when "10101011000010010" => rgb <= "000000";
					when "10101011000010011" => rgb <= "000000";
					when "10101011000010100" => rgb <= "000000";
					when "10101011000010101" => rgb <= "000000";
					when "10101011000010110" => rgb <= "000000";
					when "10101011000010111" => rgb <= "000000";
					when "10101011000011000" => rgb <= "000000";
					when "10101011000011001" => rgb <= "000000";
					when "10101011000011010" => rgb <= "000000";
					when "10101011000011011" => rgb <= "000000";
					when "10101011000011100" => rgb <= "000000";
					when "10101011000011101" => rgb <= "000000";
					when "10101011000011110" => rgb <= "000000";
					when "10101011000011111" => rgb <= "000000";
					when "10101011000100000" => rgb <= "000000";
					when "10101011000100001" => rgb <= "000000";
					when "10101011000100010" => rgb <= "000000";
					when "10101011000100011" => rgb <= "101010";
					when "10101011000100100" => rgb <= "101010";
					when "10101011000100101" => rgb <= "101010";
					when "10101011000100110" => rgb <= "111111";
					when "10101011000100111" => rgb <= "111111";
					when "10101011000101000" => rgb <= "111111";
					when "10101011000101001" => rgb <= "111111";
					when "10101011000101010" => rgb <= "101010";
					when "10101011000101011" => rgb <= "111111";
					when "10101011000101100" => rgb <= "111111";
					when "10101011000101101" => rgb <= "111111";
					when "10101011000101110" => rgb <= "111111";
					when "10101011000101111" => rgb <= "101010";
					when "10101011000110000" => rgb <= "111111";
					when "10101011000110001" => rgb <= "101010";
					when "10101011000110010" => rgb <= "000000";
					when "10101011000110011" => rgb <= "000000";
					when "10101011000110100" => rgb <= "000000";
					when "10101011000110101" => rgb <= "000000";
					when "10101011000110110" => rgb <= "000000";
					when "10101011000110111" => rgb <= "000000";
					when "10101011000111000" => rgb <= "000000";
					when "10101011000111001" => rgb <= "010101";
					when "10101011000111010" => rgb <= "111111";
					when "10101011000111011" => rgb <= "101010";
					when "10101011000111100" => rgb <= "111111";
					when "10101011000111101" => rgb <= "111111";
					when "10101011000111110" => rgb <= "111111";
					when "10101011000111111" => rgb <= "101010";
					when "10101011001000000" => rgb <= "101010";
					when "10101011001000001" => rgb <= "000000";
					when "10101011001000010" => rgb <= "000000";
					when "10101011001000011" => rgb <= "000000";
					when "10101011001000100" => rgb <= "000000";
					when "10101011001000101" => rgb <= "000000";
					when "10101011001000110" => rgb <= "000000";
					when "10101011001000111" => rgb <= "000000";
					when "10101011001001000" => rgb <= "000000";
					when "10101011001001001" => rgb <= "000000";
					when "10101011001001010" => rgb <= "000000";
					when "10101011001001011" => rgb <= "000000";
					when "10101011001001100" => rgb <= "000000";
					when "10101011001001101" => rgb <= "000000";
					when "10101011001001110" => rgb <= "000000";
					when "10101011001001111" => rgb <= "000000";
					when "10101011001010000" => rgb <= "101010";
					when "10101011001010001" => rgb <= "111111";
					when "10101011001010010" => rgb <= "101010";
					when "10101011001010011" => rgb <= "101010";
					when "10101011001010100" => rgb <= "111111";
					when "10101011001010101" => rgb <= "111111";
					when "10101011001010110" => rgb <= "101010";
					when "10101011001010111" => rgb <= "111111";
					when "10101011001011000" => rgb <= "111111";
					when "10101011001011001" => rgb <= "101010";
					when "10101011001011010" => rgb <= "111111";
					when "10101011001011011" => rgb <= "111111";
					when "10101011001011100" => rgb <= "101010";
					when "10101011001011101" => rgb <= "101010";
					when "10101011001011110" => rgb <= "101010";
					when "10101011001011111" => rgb <= "000000";
					when "10101011001100000" => rgb <= "000000";
					when "10101011001100001" => rgb <= "000000";
					when "10101011001100010" => rgb <= "000000";
					when "10101011001100011" => rgb <= "000000";
					when "10101011001100100" => rgb <= "000000";
					when "10101011001100101" => rgb <= "000000";
					when "10101011001100110" => rgb <= "010101";
					when "10101011001100111" => rgb <= "111111";
					when "10101011001101000" => rgb <= "101010";
					when "10101011001101001" => rgb <= "111111";
					when "10101011001101010" => rgb <= "101010";
					when "10101011001101011" => rgb <= "101010";
					when "10101011001101100" => rgb <= "101010";
					when "10101011001101101" => rgb <= "111111";
					when "10101011001101110" => rgb <= "000000";
					when "10101011001101111" => rgb <= "000000";
					when "10101011001110000" => rgb <= "000000";
					when "10101011001110001" => rgb <= "000000";
					when "10101011001110010" => rgb <= "000000";
					when "10101011001110011" => rgb <= "000000";
					when "10101011001110100" => rgb <= "000000";
					when "10101011001110101" => rgb <= "000000";
					when "10101011001110110" => rgb <= "000000";
					when "10101011001110111" => rgb <= "000000";
					when "10101011001111000" => rgb <= "000000";
					when "10101011001111001" => rgb <= "000000";
					when "10101011001111010" => rgb <= "000000";
					when "10101011001111011" => rgb <= "000000";
					when "10101011001111100" => rgb <= "000000";
					when "10101011001111101" => rgb <= "101010";
					when "10101011001111110" => rgb <= "111111";
					when "10101011001111111" => rgb <= "111111";
					when "10101011010000000" => rgb <= "111111";
					when "10101011010000001" => rgb <= "111111";
					when "10101011010000010" => rgb <= "111111";
					when "10101011010000011" => rgb <= "111111";
					when "10101011010000100" => rgb <= "111111";
					when "10101011010000101" => rgb <= "111111";
					when "10101011010000110" => rgb <= "111111";
					when "10101011010000111" => rgb <= "111111";
					when "10101011010001000" => rgb <= "111111";
					when "10101011010001001" => rgb <= "101010";
					when "10101011010001010" => rgb <= "111111";
					when "10101011010001011" => rgb <= "101010";
					when "10101011010001100" => rgb <= "000000";
					when "10101011010001101" => rgb <= "000000";
					when "10101011010001110" => rgb <= "000000";
					when "10101011010001111" => rgb <= "000000";
					when "10101011010010000" => rgb <= "000000";
					when "10101011010010001" => rgb <= "000000";
					when "10101011010010010" => rgb <= "000000";
					when "10101011010010011" => rgb <= "000000";
					when "10101011010010100" => rgb <= "000000";
					when "10101011010010101" => rgb <= "000000";
					when "10101011010010110" => rgb <= "000000";
					when "10101011010010111" => rgb <= "000000";
					when "10101011010011000" => rgb <= "000000";
					when "10101011010011001" => rgb <= "000000";
					when "10101011010011010" => rgb <= "000000";
					when "10101011010011011" => rgb <= "000000";
					when "10101011010011100" => rgb <= "000000";
					when "10101011010011101" => rgb <= "000000";
					when "10101011010011110" => rgb <= "000000";
					when "10101011010011111" => rgb <= "000000";
					when "10101011010100000" => rgb <= "000000";
					when "10101011010100001" => rgb <= "000000";
					when "10101011010100010" => rgb <= "010101";
					when "10101011010100011" => rgb <= "111111";
					when "10101011010100100" => rgb <= "101010";
					when "10101011010100101" => rgb <= "111111";
					when "10101011010100110" => rgb <= "111111";
					when "10101011010100111" => rgb <= "111111";
					when "10101011010101000" => rgb <= "111111";
					when "10101011010101001" => rgb <= "111111";
					when "10101011010101010" => rgb <= "000000";
					when "10101011010101011" => rgb <= "000000";
					when "10101011010101100" => rgb <= "000000";
					when "10101011010101101" => rgb <= "000000";
					when "10101011010101110" => rgb <= "000000";
					when "10101011010101111" => rgb <= "000000";
					when "10101011010110000" => rgb <= "000000";
					when "10101011010110001" => rgb <= "000000";
					when "10101011010110010" => rgb <= "000000";
					when "10101011010110011" => rgb <= "000000";
					when "10101011010110100" => rgb <= "000000";
					when "10101011010110101" => rgb <= "000000";
					when "10101011010110110" => rgb <= "000000";
					when "10101011010110111" => rgb <= "000000";
					when "10101011010111000" => rgb <= "000000";
					when "10101011010111001" => rgb <= "000000";
					when "10101011010111010" => rgb <= "000000";
					when "10101011010111011" => rgb <= "000000";
					when "10101011010111100" => rgb <= "000000";
					when "10101011010111101" => rgb <= "000000";
					when "10101011010111110" => rgb <= "000000";
					when "10101011010111111" => rgb <= "000000";
					when "10101011011000000" => rgb <= "010101";
					when "10101011011000001" => rgb <= "101010";
					when "10101011011000010" => rgb <= "101010";
					when "10101011011000011" => rgb <= "111111";
					when "10101011011000100" => rgb <= "111111";
					when "10101011011000101" => rgb <= "111111";
					when "10101011011000110" => rgb <= "111111";
					when "10101011011000111" => rgb <= "111111";
					when "10101011011001000" => rgb <= "111111";
					when "10101011011001001" => rgb <= "101010";
					when "10101011011001010" => rgb <= "111111";
					when "10101011011001011" => rgb <= "101010";
					when "10101011011001100" => rgb <= "111111";
					when "10101011011001101" => rgb <= "101010";
					when "10101011011001110" => rgb <= "111111";
					when "10101011011001111" => rgb <= "010101";
					when "10101011011010000" => rgb <= "000000";
					when "10101011011010001" => rgb <= "000000";
					when "10101011011010010" => rgb <= "000000";
					when "10101011011010011" => rgb <= "000000";
					when "10101011011010100" => rgb <= "000000";
					when "10101011011010101" => rgb <= "000000";
					when "10101011011010110" => rgb <= "000000";
					when "10101011011010111" => rgb <= "101010";
					when "10101011011011000" => rgb <= "101010";
					when "10101011011011001" => rgb <= "101010";
					when "10101011011011010" => rgb <= "101010";
					when "10101011011011011" => rgb <= "111111";
					when "10101011011011100" => rgb <= "111111";
					when "10101011011011101" => rgb <= "111111";
					when "10101011011011110" => rgb <= "111111";
					when "10101011011011111" => rgb <= "111111";
					when "10101011011100000" => rgb <= "111111";
					when "10101011011100001" => rgb <= "111111";
					when "10101011011100010" => rgb <= "101010";
					when "10101011011100011" => rgb <= "101010";
					when "10101011011100100" => rgb <= "101010";
					when "10101011011100101" => rgb <= "101010";
					when "10101011011100110" => rgb <= "000000";
					when "10101011011100111" => rgb <= "000000";
					when "10101011011101000" => rgb <= "000000";
					when "10101011011101001" => rgb <= "000000";
					when "10101011011101010" => rgb <= "000000";
					when "10101011011101011" => rgb <= "000000";
					when "10101011011101100" => rgb <= "000000";
					when "10101011011101101" => rgb <= "010101";
					when "10101011011101110" => rgb <= "111111";
					when "10101011011101111" => rgb <= "101010";
					when "10101011011110000" => rgb <= "101010";
					when "10101011011110001" => rgb <= "101010";
					when "10101011011110010" => rgb <= "111111";
					when "10101011011110011" => rgb <= "111111";
					when "10101011011110100" => rgb <= "111111";
					when "10101011011110101" => rgb <= "111111";
					when "10101011011110110" => rgb <= "111111";
					when "10101011011110111" => rgb <= "111111";
					when "10101011011111000" => rgb <= "101010";
					when "10101011011111001" => rgb <= "111111";
					when "10101011011111010" => rgb <= "101010";
					when "10101011011111011" => rgb <= "111111";
					when "10101011011111100" => rgb <= "010101";
					when "10101011011111101" => rgb <= "000000";
					when "10101011011111110" => rgb <= "000000";
					when "10101011011111111" => rgb <= "000000";
					when "10101011100000000" => rgb <= "000000";
					when "10101011100000001" => rgb <= "000000";
					when "10101011100000010" => rgb <= "000000";
					when "10101011100000011" => rgb <= "000000";
					when "10101011100000100" => rgb <= "000000";
					when "10101011100000101" => rgb <= "000000";
					when "10101011100000110" => rgb <= "000000";
					when "10101011100000111" => rgb <= "000000";
					when "10101011100001000" => rgb <= "000000";
					when "10101011100001001" => rgb <= "000000";
					when "10101011100001010" => rgb <= "000000";
					when "10101011100001011" => rgb <= "010101";
					when "10101011100001100" => rgb <= "111111";
					when "10101011100001101" => rgb <= "101010";
					when "10101011100001110" => rgb <= "111111";
					when "10101011100001111" => rgb <= "111111";
					when "10101011100010000" => rgb <= "111111";
					when "10101011100010001" => rgb <= "111111";
					when "10101011100010010" => rgb <= "111111";
					when "10101011100010011" => rgb <= "111111";
					when "10101011100010100" => rgb <= "111111";
					when "10101011100010101" => rgb <= "111111";
					when "10101011100010110" => rgb <= "111111";
					when "10101011100010111" => rgb <= "111111";
					when "10101011100011000" => rgb <= "101010";
					when "10101011100011001" => rgb <= "111111";
					when "10101011100011010" => rgb <= "101010";
					when "10101011100011011" => rgb <= "000000";
					when "10101011100011100" => rgb <= "000000";
					when "10101011100011101" => rgb <= "000000";
					when "10101011100011110" => rgb <= "000000";
					when "10101011100011111" => rgb <= "000000";
					when "10101011100100000" => rgb <= "000000";
					when "10101011100100001" => rgb <= "000000";
					when "10101011100100010" => rgb <= "101010";
					when "10101011100100011" => rgb <= "101010";
					when "10101011100100100" => rgb <= "101010";
					when "10101011100100101" => rgb <= "101010";
					when "10101011100100110" => rgb <= "111111";
					when "10101011100100111" => rgb <= "111111";
					when "10101011100101000" => rgb <= "101010";
					when "10101011100101001" => rgb <= "111111";
					when "10101011100101010" => rgb <= "111111";
					when "10101011100101011" => rgb <= "101010";
					when "10101011100101100" => rgb <= "111111";
					when "10101011100101101" => rgb <= "111111";
					when "10101011100101110" => rgb <= "101010";
					when "10101011100101111" => rgb <= "101010";
					when "10101011100110000" => rgb <= "111111";
					when "10101011100110001" => rgb <= "010101";
					when "10101011100110010" => rgb <= "000000";
					when "10101011100110011" => rgb <= "000000";
					when "10101011100110100" => rgb <= "000000";
					when "10101011100110101" => rgb <= "000000";
					when "10101011100110110" => rgb <= "000000";
					when "10101011100110111" => rgb <= "000000";
					when "10101011100111000" => rgb <= "000000";
					when "10101011100111001" => rgb <= "000000";
					when "10101011100111010" => rgb <= "000000";
					when "10101011100111011" => rgb <= "000000";
					when "10101011100111100" => rgb <= "000000";
					when "10101011100111101" => rgb <= "000000";
					when "10101011100111110" => rgb <= "000000";
					when "10101011100111111" => rgb <= "000000";
					when "10101100000000000" => rgb <= "000000";
					when "10101100000000001" => rgb <= "000000";
					when "10101100000000010" => rgb <= "000000";
					when "10101100000000011" => rgb <= "000000";
					when "10101100000000100" => rgb <= "000000";
					when "10101100000000101" => rgb <= "101010";
					when "10101100000000110" => rgb <= "111111";
					when "10101100000000111" => rgb <= "101010";
					when "10101100000001000" => rgb <= "111111";
					when "10101100000001001" => rgb <= "111111";
					when "10101100000001010" => rgb <= "101010";
					when "10101100000001011" => rgb <= "101010";
					when "10101100000001100" => rgb <= "101010";
					when "10101100000001101" => rgb <= "000000";
					when "10101100000001110" => rgb <= "000000";
					when "10101100000001111" => rgb <= "000000";
					when "10101100000010000" => rgb <= "000000";
					when "10101100000010001" => rgb <= "000000";
					when "10101100000010010" => rgb <= "000000";
					when "10101100000010011" => rgb <= "000000";
					when "10101100000010100" => rgb <= "000000";
					when "10101100000010101" => rgb <= "000000";
					when "10101100000010110" => rgb <= "000000";
					when "10101100000010111" => rgb <= "000000";
					when "10101100000011000" => rgb <= "000000";
					when "10101100000011001" => rgb <= "000000";
					when "10101100000011010" => rgb <= "000000";
					when "10101100000011011" => rgb <= "000000";
					when "10101100000011100" => rgb <= "000000";
					when "10101100000011101" => rgb <= "000000";
					when "10101100000011110" => rgb <= "000000";
					when "10101100000011111" => rgb <= "000000";
					when "10101100000100000" => rgb <= "000000";
					when "10101100000100001" => rgb <= "000000";
					when "10101100000100010" => rgb <= "000000";
					when "10101100000100011" => rgb <= "101010";
					when "10101100000100100" => rgb <= "111111";
					when "10101100000100101" => rgb <= "101010";
					when "10101100000100110" => rgb <= "101010";
					when "10101100000100111" => rgb <= "111111";
					when "10101100000101000" => rgb <= "111111";
					when "10101100000101001" => rgb <= "111111";
					when "10101100000101010" => rgb <= "101010";
					when "10101100000101011" => rgb <= "111111";
					when "10101100000101100" => rgb <= "111111";
					when "10101100000101101" => rgb <= "111111";
					when "10101100000101110" => rgb <= "111111";
					when "10101100000101111" => rgb <= "101010";
					when "10101100000110000" => rgb <= "111111";
					when "10101100000110001" => rgb <= "101010";
					when "10101100000110010" => rgb <= "000000";
					when "10101100000110011" => rgb <= "000000";
					when "10101100000110100" => rgb <= "000000";
					when "10101100000110101" => rgb <= "000000";
					when "10101100000110110" => rgb <= "000000";
					when "10101100000110111" => rgb <= "000000";
					when "10101100000111000" => rgb <= "000000";
					when "10101100000111001" => rgb <= "010101";
					when "10101100000111010" => rgb <= "101010";
					when "10101100000111011" => rgb <= "101010";
					when "10101100000111100" => rgb <= "111111";
					when "10101100000111101" => rgb <= "101010";
					when "10101100000111110" => rgb <= "111111";
					when "10101100000111111" => rgb <= "111111";
					when "10101100001000000" => rgb <= "101010";
					when "10101100001000001" => rgb <= "000000";
					when "10101100001000010" => rgb <= "000000";
					when "10101100001000011" => rgb <= "000000";
					when "10101100001000100" => rgb <= "000000";
					when "10101100001000101" => rgb <= "000000";
					when "10101100001000110" => rgb <= "000000";
					when "10101100001000111" => rgb <= "000000";
					when "10101100001001000" => rgb <= "000000";
					when "10101100001001001" => rgb <= "000000";
					when "10101100001001010" => rgb <= "000000";
					when "10101100001001011" => rgb <= "000000";
					when "10101100001001100" => rgb <= "000000";
					when "10101100001001101" => rgb <= "000000";
					when "10101100001001110" => rgb <= "000000";
					when "10101100001001111" => rgb <= "000000";
					when "10101100001010000" => rgb <= "101010";
					when "10101100001010001" => rgb <= "111111";
					when "10101100001010010" => rgb <= "101010";
					when "10101100001010011" => rgb <= "101010";
					when "10101100001010100" => rgb <= "111111";
					when "10101100001010101" => rgb <= "111111";
					when "10101100001010110" => rgb <= "101010";
					when "10101100001010111" => rgb <= "111111";
					when "10101100001011000" => rgb <= "111111";
					when "10101100001011001" => rgb <= "111111";
					when "10101100001011010" => rgb <= "101010";
					when "10101100001011011" => rgb <= "111111";
					when "10101100001011100" => rgb <= "111111";
					when "10101100001011101" => rgb <= "101010";
					when "10101100001011110" => rgb <= "101010";
					when "10101100001011111" => rgb <= "000000";
					when "10101100001100000" => rgb <= "000000";
					when "10101100001100001" => rgb <= "000000";
					when "10101100001100010" => rgb <= "000000";
					when "10101100001100011" => rgb <= "000000";
					when "10101100001100100" => rgb <= "000000";
					when "10101100001100101" => rgb <= "000000";
					when "10101100001100110" => rgb <= "010101";
					when "10101100001100111" => rgb <= "111111";
					when "10101100001101000" => rgb <= "101010";
					when "10101100001101001" => rgb <= "111111";
					when "10101100001101010" => rgb <= "111111";
					when "10101100001101011" => rgb <= "111111";
					when "10101100001101100" => rgb <= "111111";
					when "10101100001101101" => rgb <= "111111";
					when "10101100001101110" => rgb <= "000000";
					when "10101100001101111" => rgb <= "000000";
					when "10101100001110000" => rgb <= "000000";
					when "10101100001110001" => rgb <= "000000";
					when "10101100001110010" => rgb <= "000000";
					when "10101100001110011" => rgb <= "000000";
					when "10101100001110100" => rgb <= "000000";
					when "10101100001110101" => rgb <= "000000";
					when "10101100001110110" => rgb <= "000000";
					when "10101100001110111" => rgb <= "000000";
					when "10101100001111000" => rgb <= "000000";
					when "10101100001111001" => rgb <= "000000";
					when "10101100001111010" => rgb <= "000000";
					when "10101100001111011" => rgb <= "000000";
					when "10101100001111100" => rgb <= "000000";
					when "10101100001111101" => rgb <= "101010";
					when "10101100001111110" => rgb <= "111111";
					when "10101100001111111" => rgb <= "111111";
					when "10101100010000000" => rgb <= "111111";
					when "10101100010000001" => rgb <= "111111";
					when "10101100010000010" => rgb <= "111111";
					when "10101100010000011" => rgb <= "111111";
					when "10101100010000100" => rgb <= "111111";
					when "10101100010000101" => rgb <= "111111";
					when "10101100010000110" => rgb <= "111111";
					when "10101100010000111" => rgb <= "111111";
					when "10101100010001000" => rgb <= "111111";
					when "10101100010001001" => rgb <= "101010";
					when "10101100010001010" => rgb <= "111111";
					when "10101100010001011" => rgb <= "101010";
					when "10101100010001100" => rgb <= "000000";
					when "10101100010001101" => rgb <= "000000";
					when "10101100010001110" => rgb <= "000000";
					when "10101100010001111" => rgb <= "000000";
					when "10101100010010000" => rgb <= "000000";
					when "10101100010010001" => rgb <= "000000";
					when "10101100010010010" => rgb <= "000000";
					when "10101100010010011" => rgb <= "000000";
					when "10101100010010100" => rgb <= "000000";
					when "10101100010010101" => rgb <= "000000";
					when "10101100010010110" => rgb <= "000000";
					when "10101100010010111" => rgb <= "000000";
					when "10101100010011000" => rgb <= "000000";
					when "10101100010011001" => rgb <= "000000";
					when "10101100010011010" => rgb <= "000000";
					when "10101100010011011" => rgb <= "000000";
					when "10101100010011100" => rgb <= "000000";
					when "10101100010011101" => rgb <= "000000";
					when "10101100010011110" => rgb <= "000000";
					when "10101100010011111" => rgb <= "000000";
					when "10101100010100000" => rgb <= "000000";
					when "10101100010100001" => rgb <= "000000";
					when "10101100010100010" => rgb <= "010101";
					when "10101100010100011" => rgb <= "111111";
					when "10101100010100100" => rgb <= "101010";
					when "10101100010100101" => rgb <= "111111";
					when "10101100010100110" => rgb <= "111111";
					when "10101100010100111" => rgb <= "111111";
					when "10101100010101000" => rgb <= "111111";
					when "10101100010101001" => rgb <= "111111";
					when "10101100010101010" => rgb <= "000000";
					when "10101100010101011" => rgb <= "000000";
					when "10101100010101100" => rgb <= "000000";
					when "10101100010101101" => rgb <= "000000";
					when "10101100010101110" => rgb <= "000000";
					when "10101100010101111" => rgb <= "000000";
					when "10101100010110000" => rgb <= "000000";
					when "10101100010110001" => rgb <= "000000";
					when "10101100010110010" => rgb <= "000000";
					when "10101100010110011" => rgb <= "000000";
					when "10101100010110100" => rgb <= "000000";
					when "10101100010110101" => rgb <= "000000";
					when "10101100010110110" => rgb <= "000000";
					when "10101100010110111" => rgb <= "000000";
					when "10101100010111000" => rgb <= "000000";
					when "10101100010111001" => rgb <= "000000";
					when "10101100010111010" => rgb <= "000000";
					when "10101100010111011" => rgb <= "000000";
					when "10101100010111100" => rgb <= "000000";
					when "10101100010111101" => rgb <= "000000";
					when "10101100010111110" => rgb <= "000000";
					when "10101100010111111" => rgb <= "000000";
					when "10101100011000000" => rgb <= "010101";
					when "10101100011000001" => rgb <= "101010";
					when "10101100011000010" => rgb <= "101010";
					when "10101100011000011" => rgb <= "111111";
					when "10101100011000100" => rgb <= "111111";
					when "10101100011000101" => rgb <= "111111";
					when "10101100011000110" => rgb <= "111111";
					when "10101100011000111" => rgb <= "111111";
					when "10101100011001000" => rgb <= "111111";
					when "10101100011001001" => rgb <= "101010";
					when "10101100011001010" => rgb <= "111111";
					when "10101100011001011" => rgb <= "101010";
					when "10101100011001100" => rgb <= "111111";
					when "10101100011001101" => rgb <= "101010";
					when "10101100011001110" => rgb <= "111111";
					when "10101100011001111" => rgb <= "010101";
					when "10101100011010000" => rgb <= "000000";
					when "10101100011010001" => rgb <= "000000";
					when "10101100011010010" => rgb <= "000000";
					when "10101100011010011" => rgb <= "000000";
					when "10101100011010100" => rgb <= "000000";
					when "10101100011010101" => rgb <= "000000";
					when "10101100011010110" => rgb <= "000000";
					when "10101100011010111" => rgb <= "101010";
					when "10101100011011000" => rgb <= "101010";
					when "10101100011011001" => rgb <= "101010";
					when "10101100011011010" => rgb <= "101010";
					when "10101100011011011" => rgb <= "111111";
					when "10101100011011100" => rgb <= "111111";
					when "10101100011011101" => rgb <= "111111";
					when "10101100011011110" => rgb <= "111111";
					when "10101100011011111" => rgb <= "111111";
					when "10101100011100000" => rgb <= "111111";
					when "10101100011100001" => rgb <= "111111";
					when "10101100011100010" => rgb <= "111111";
					when "10101100011100011" => rgb <= "101010";
					when "10101100011100100" => rgb <= "111111";
					when "10101100011100101" => rgb <= "111111";
					when "10101100011100110" => rgb <= "000000";
					when "10101100011100111" => rgb <= "000000";
					when "10101100011101000" => rgb <= "000000";
					when "10101100011101001" => rgb <= "000000";
					when "10101100011101010" => rgb <= "000000";
					when "10101100011101011" => rgb <= "000000";
					when "10101100011101100" => rgb <= "000000";
					when "10101100011101101" => rgb <= "010101";
					when "10101100011101110" => rgb <= "111111";
					when "10101100011101111" => rgb <= "101010";
					when "10101100011110000" => rgb <= "111111";
					when "10101100011110001" => rgb <= "111111";
					when "10101100011110010" => rgb <= "101010";
					when "10101100011110011" => rgb <= "111111";
					when "10101100011110100" => rgb <= "101010";
					when "10101100011110101" => rgb <= "101010";
					when "10101100011110110" => rgb <= "101010";
					when "10101100011110111" => rgb <= "111111";
					when "10101100011111000" => rgb <= "111111";
					when "10101100011111001" => rgb <= "111111";
					when "10101100011111010" => rgb <= "101010";
					when "10101100011111011" => rgb <= "111111";
					when "10101100011111100" => rgb <= "010101";
					when "10101100011111101" => rgb <= "000000";
					when "10101100011111110" => rgb <= "000000";
					when "10101100011111111" => rgb <= "000000";
					when "10101100100000000" => rgb <= "000000";
					when "10101100100000001" => rgb <= "000000";
					when "10101100100000010" => rgb <= "000000";
					when "10101100100000011" => rgb <= "000000";
					when "10101100100000100" => rgb <= "000000";
					when "10101100100000101" => rgb <= "000000";
					when "10101100100000110" => rgb <= "000000";
					when "10101100100000111" => rgb <= "000000";
					when "10101100100001000" => rgb <= "000000";
					when "10101100100001001" => rgb <= "000000";
					when "10101100100001010" => rgb <= "000000";
					when "10101100100001011" => rgb <= "010101";
					when "10101100100001100" => rgb <= "111111";
					when "10101100100001101" => rgb <= "101010";
					when "10101100100001110" => rgb <= "111111";
					when "10101100100001111" => rgb <= "111111";
					when "10101100100010000" => rgb <= "111111";
					when "10101100100010001" => rgb <= "111111";
					when "10101100100010010" => rgb <= "111111";
					when "10101100100010011" => rgb <= "111111";
					when "10101100100010100" => rgb <= "111111";
					when "10101100100010101" => rgb <= "111111";
					when "10101100100010110" => rgb <= "111111";
					when "10101100100010111" => rgb <= "111111";
					when "10101100100011000" => rgb <= "101010";
					when "10101100100011001" => rgb <= "111111";
					when "10101100100011010" => rgb <= "101010";
					when "10101100100011011" => rgb <= "000000";
					when "10101100100011100" => rgb <= "000000";
					when "10101100100011101" => rgb <= "000000";
					when "10101100100011110" => rgb <= "000000";
					when "10101100100011111" => rgb <= "000000";
					when "10101100100100000" => rgb <= "000000";
					when "10101100100100001" => rgb <= "000000";
					when "10101100100100010" => rgb <= "101010";
					when "10101100100100011" => rgb <= "101010";
					when "10101100100100100" => rgb <= "101010";
					when "10101100100100101" => rgb <= "101010";
					when "10101100100100110" => rgb <= "111111";
					when "10101100100100111" => rgb <= "111111";
					when "10101100100101000" => rgb <= "101010";
					when "10101100100101001" => rgb <= "111111";
					when "10101100100101010" => rgb <= "111111";
					when "10101100100101011" => rgb <= "101010";
					when "10101100100101100" => rgb <= "111111";
					when "10101100100101101" => rgb <= "111111";
					when "10101100100101110" => rgb <= "101010";
					when "10101100100101111" => rgb <= "101010";
					when "10101100100110000" => rgb <= "111111";
					when "10101100100110001" => rgb <= "010101";
					when "10101100100110010" => rgb <= "000000";
					when "10101100100110011" => rgb <= "000000";
					when "10101100100110100" => rgb <= "000000";
					when "10101100100110101" => rgb <= "000000";
					when "10101100100110110" => rgb <= "000000";
					when "10101100100110111" => rgb <= "000000";
					when "10101100100111000" => rgb <= "000000";
					when "10101100100111001" => rgb <= "000000";
					when "10101100100111010" => rgb <= "000000";
					when "10101100100111011" => rgb <= "000000";
					when "10101100100111100" => rgb <= "000000";
					when "10101100100111101" => rgb <= "000000";
					when "10101100100111110" => rgb <= "000000";
					when "10101100100111111" => rgb <= "000000";
					when "10101101000000000" => rgb <= "000000";
					when "10101101000000001" => rgb <= "000000";
					when "10101101000000010" => rgb <= "000000";
					when "10101101000000011" => rgb <= "000000";
					when "10101101000000100" => rgb <= "000000";
					when "10101101000000101" => rgb <= "101010";
					when "10101101000000110" => rgb <= "111111";
					when "10101101000000111" => rgb <= "101010";
					when "10101101000001000" => rgb <= "111111";
					when "10101101000001001" => rgb <= "111111";
					when "10101101000001010" => rgb <= "101010";
					when "10101101000001011" => rgb <= "101010";
					when "10101101000001100" => rgb <= "101010";
					when "10101101000001101" => rgb <= "000000";
					when "10101101000001110" => rgb <= "000000";
					when "10101101000001111" => rgb <= "000000";
					when "10101101000010000" => rgb <= "000000";
					when "10101101000010001" => rgb <= "000000";
					when "10101101000010010" => rgb <= "000000";
					when "10101101000010011" => rgb <= "000000";
					when "10101101000010100" => rgb <= "000000";
					when "10101101000010101" => rgb <= "000000";
					when "10101101000010110" => rgb <= "000000";
					when "10101101000010111" => rgb <= "000000";
					when "10101101000011000" => rgb <= "000000";
					when "10101101000011001" => rgb <= "000000";
					when "10101101000011010" => rgb <= "000000";
					when "10101101000011011" => rgb <= "000000";
					when "10101101000011100" => rgb <= "000000";
					when "10101101000011101" => rgb <= "000000";
					when "10101101000011110" => rgb <= "000000";
					when "10101101000011111" => rgb <= "000000";
					when "10101101000100000" => rgb <= "000000";
					when "10101101000100001" => rgb <= "000000";
					when "10101101000100010" => rgb <= "000000";
					when "10101101000100011" => rgb <= "101010";
					when "10101101000100100" => rgb <= "111111";
					when "10101101000100101" => rgb <= "101010";
					when "10101101000100110" => rgb <= "101010";
					when "10101101000100111" => rgb <= "111111";
					when "10101101000101000" => rgb <= "111111";
					when "10101101000101001" => rgb <= "111111";
					when "10101101000101010" => rgb <= "101010";
					when "10101101000101011" => rgb <= "111111";
					when "10101101000101100" => rgb <= "111111";
					when "10101101000101101" => rgb <= "111111";
					when "10101101000101110" => rgb <= "111111";
					when "10101101000101111" => rgb <= "101010";
					when "10101101000110000" => rgb <= "111111";
					when "10101101000110001" => rgb <= "101010";
					when "10101101000110010" => rgb <= "000000";
					when "10101101000110011" => rgb <= "000000";
					when "10101101000110100" => rgb <= "000000";
					when "10101101000110101" => rgb <= "000000";
					when "10101101000110110" => rgb <= "000000";
					when "10101101000110111" => rgb <= "000000";
					when "10101101000111000" => rgb <= "000000";
					when "10101101000111001" => rgb <= "010101";
					when "10101101000111010" => rgb <= "101010";
					when "10101101000111011" => rgb <= "101010";
					when "10101101000111100" => rgb <= "101010";
					when "10101101000111101" => rgb <= "101010";
					when "10101101000111110" => rgb <= "111111";
					when "10101101000111111" => rgb <= "111111";
					when "10101101001000000" => rgb <= "101010";
					when "10101101001000001" => rgb <= "000000";
					when "10101101001000010" => rgb <= "000000";
					when "10101101001000011" => rgb <= "000000";
					when "10101101001000100" => rgb <= "000000";
					when "10101101001000101" => rgb <= "000000";
					when "10101101001000110" => rgb <= "000000";
					when "10101101001000111" => rgb <= "000000";
					when "10101101001001000" => rgb <= "000000";
					when "10101101001001001" => rgb <= "000000";
					when "10101101001001010" => rgb <= "000000";
					when "10101101001001011" => rgb <= "000000";
					when "10101101001001100" => rgb <= "000000";
					when "10101101001001101" => rgb <= "000000";
					when "10101101001001110" => rgb <= "000000";
					when "10101101001001111" => rgb <= "000000";
					when "10101101001010000" => rgb <= "101010";
					when "10101101001010001" => rgb <= "101010";
					when "10101101001010010" => rgb <= "101010";
					when "10101101001010011" => rgb <= "111111";
					when "10101101001010100" => rgb <= "111111";
					when "10101101001010101" => rgb <= "101010";
					when "10101101001010110" => rgb <= "101010";
					when "10101101001010111" => rgb <= "111111";
					when "10101101001011000" => rgb <= "101010";
					when "10101101001011001" => rgb <= "111111";
					when "10101101001011010" => rgb <= "101010";
					when "10101101001011011" => rgb <= "101010";
					when "10101101001011100" => rgb <= "111111";
					when "10101101001011101" => rgb <= "111111";
					when "10101101001011110" => rgb <= "101010";
					when "10101101001011111" => rgb <= "000000";
					when "10101101001100000" => rgb <= "000000";
					when "10101101001100001" => rgb <= "000000";
					when "10101101001100010" => rgb <= "000000";
					when "10101101001100011" => rgb <= "000000";
					when "10101101001100100" => rgb <= "000000";
					when "10101101001100101" => rgb <= "000000";
					when "10101101001100110" => rgb <= "010101";
					when "10101101001100111" => rgb <= "111111";
					when "10101101001101000" => rgb <= "101010";
					when "10101101001101001" => rgb <= "111111";
					when "10101101001101010" => rgb <= "101010";
					when "10101101001101011" => rgb <= "101010";
					when "10101101001101100" => rgb <= "101010";
					when "10101101001101101" => rgb <= "101010";
					when "10101101001101110" => rgb <= "000000";
					when "10101101001101111" => rgb <= "000000";
					when "10101101001110000" => rgb <= "000000";
					when "10101101001110001" => rgb <= "000000";
					when "10101101001110010" => rgb <= "000000";
					when "10101101001110011" => rgb <= "000000";
					when "10101101001110100" => rgb <= "000000";
					when "10101101001110101" => rgb <= "000000";
					when "10101101001110110" => rgb <= "000000";
					when "10101101001110111" => rgb <= "000000";
					when "10101101001111000" => rgb <= "000000";
					when "10101101001111001" => rgb <= "000000";
					when "10101101001111010" => rgb <= "000000";
					when "10101101001111011" => rgb <= "000000";
					when "10101101001111100" => rgb <= "000000";
					when "10101101001111101" => rgb <= "101010";
					when "10101101001111110" => rgb <= "111111";
					when "10101101001111111" => rgb <= "111111";
					when "10101101010000000" => rgb <= "111111";
					when "10101101010000001" => rgb <= "111111";
					when "10101101010000010" => rgb <= "111111";
					when "10101101010000011" => rgb <= "111111";
					when "10101101010000100" => rgb <= "111111";
					when "10101101010000101" => rgb <= "111111";
					when "10101101010000110" => rgb <= "111111";
					when "10101101010000111" => rgb <= "111111";
					when "10101101010001000" => rgb <= "111111";
					when "10101101010001001" => rgb <= "111111";
					when "10101101010001010" => rgb <= "111111";
					when "10101101010001011" => rgb <= "101010";
					when "10101101010001100" => rgb <= "000000";
					when "10101101010001101" => rgb <= "000000";
					when "10101101010001110" => rgb <= "000000";
					when "10101101010001111" => rgb <= "000000";
					when "10101101010010000" => rgb <= "000000";
					when "10101101010010001" => rgb <= "000000";
					when "10101101010010010" => rgb <= "000000";
					when "10101101010010011" => rgb <= "000000";
					when "10101101010010100" => rgb <= "000000";
					when "10101101010010101" => rgb <= "000000";
					when "10101101010010110" => rgb <= "000000";
					when "10101101010010111" => rgb <= "000000";
					when "10101101010011000" => rgb <= "000000";
					when "10101101010011001" => rgb <= "000000";
					when "10101101010011010" => rgb <= "000000";
					when "10101101010011011" => rgb <= "000000";
					when "10101101010011100" => rgb <= "000000";
					when "10101101010011101" => rgb <= "000000";
					when "10101101010011110" => rgb <= "000000";
					when "10101101010011111" => rgb <= "000000";
					when "10101101010100000" => rgb <= "000000";
					when "10101101010100001" => rgb <= "000000";
					when "10101101010100010" => rgb <= "010101";
					when "10101101010100011" => rgb <= "111111";
					when "10101101010100100" => rgb <= "101010";
					when "10101101010100101" => rgb <= "111111";
					when "10101101010100110" => rgb <= "111111";
					when "10101101010100111" => rgb <= "111111";
					when "10101101010101000" => rgb <= "101010";
					when "10101101010101001" => rgb <= "101010";
					when "10101101010101010" => rgb <= "000000";
					when "10101101010101011" => rgb <= "000000";
					when "10101101010101100" => rgb <= "000000";
					when "10101101010101101" => rgb <= "000000";
					when "10101101010101110" => rgb <= "000000";
					when "10101101010101111" => rgb <= "000000";
					when "10101101010110000" => rgb <= "000000";
					when "10101101010110001" => rgb <= "000000";
					when "10101101010110010" => rgb <= "000000";
					when "10101101010110011" => rgb <= "000000";
					when "10101101010110100" => rgb <= "000000";
					when "10101101010110101" => rgb <= "000000";
					when "10101101010110110" => rgb <= "000000";
					when "10101101010110111" => rgb <= "000000";
					when "10101101010111000" => rgb <= "000000";
					when "10101101010111001" => rgb <= "000000";
					when "10101101010111010" => rgb <= "000000";
					when "10101101010111011" => rgb <= "000000";
					when "10101101010111100" => rgb <= "000000";
					when "10101101010111101" => rgb <= "000000";
					when "10101101010111110" => rgb <= "000000";
					when "10101101010111111" => rgb <= "000000";
					when "10101101011000000" => rgb <= "010101";
					when "10101101011000001" => rgb <= "101010";
					when "10101101011000010" => rgb <= "101010";
					when "10101101011000011" => rgb <= "111111";
					when "10101101011000100" => rgb <= "111111";
					when "10101101011000101" => rgb <= "111111";
					when "10101101011000110" => rgb <= "111111";
					when "10101101011000111" => rgb <= "111111";
					when "10101101011001000" => rgb <= "111111";
					when "10101101011001001" => rgb <= "101010";
					when "10101101011001010" => rgb <= "111111";
					when "10101101011001011" => rgb <= "101010";
					when "10101101011001100" => rgb <= "111111";
					when "10101101011001101" => rgb <= "101010";
					when "10101101011001110" => rgb <= "111111";
					when "10101101011001111" => rgb <= "010101";
					when "10101101011010000" => rgb <= "000000";
					when "10101101011010001" => rgb <= "000000";
					when "10101101011010010" => rgb <= "000000";
					when "10101101011010011" => rgb <= "000000";
					when "10101101011010100" => rgb <= "000000";
					when "10101101011010101" => rgb <= "000000";
					when "10101101011010110" => rgb <= "000000";
					when "10101101011010111" => rgb <= "101010";
					when "10101101011011000" => rgb <= "101010";
					when "10101101011011001" => rgb <= "101010";
					when "10101101011011010" => rgb <= "101010";
					when "10101101011011011" => rgb <= "111111";
					when "10101101011011100" => rgb <= "111111";
					when "10101101011011101" => rgb <= "111111";
					when "10101101011011110" => rgb <= "111111";
					when "10101101011011111" => rgb <= "111111";
					when "10101101011100000" => rgb <= "111111";
					when "10101101011100001" => rgb <= "111111";
					when "10101101011100010" => rgb <= "111111";
					when "10101101011100011" => rgb <= "111111";
					when "10101101011100100" => rgb <= "111111";
					when "10101101011100101" => rgb <= "111111";
					when "10101101011100110" => rgb <= "000000";
					when "10101101011100111" => rgb <= "000000";
					when "10101101011101000" => rgb <= "000000";
					when "10101101011101001" => rgb <= "000000";
					when "10101101011101010" => rgb <= "000000";
					when "10101101011101011" => rgb <= "000000";
					when "10101101011101100" => rgb <= "000000";
					when "10101101011101101" => rgb <= "010101";
					when "10101101011101110" => rgb <= "111111";
					when "10101101011101111" => rgb <= "101010";
					when "10101101011110000" => rgb <= "101010";
					when "10101101011110001" => rgb <= "111111";
					when "10101101011110010" => rgb <= "111111";
					when "10101101011110011" => rgb <= "111111";
					when "10101101011110100" => rgb <= "101010";
					when "10101101011110101" => rgb <= "101010";
					when "10101101011110110" => rgb <= "101010";
					when "10101101011110111" => rgb <= "111111";
					when "10101101011111000" => rgb <= "101010";
					when "10101101011111001" => rgb <= "101010";
					when "10101101011111010" => rgb <= "101010";
					when "10101101011111011" => rgb <= "111111";
					when "10101101011111100" => rgb <= "010101";
					when "10101101011111101" => rgb <= "000000";
					when "10101101011111110" => rgb <= "000000";
					when "10101101011111111" => rgb <= "000000";
					when "10101101100000000" => rgb <= "000000";
					when "10101101100000001" => rgb <= "000000";
					when "10101101100000010" => rgb <= "000000";
					when "10101101100000011" => rgb <= "000000";
					when "10101101100000100" => rgb <= "000000";
					when "10101101100000101" => rgb <= "000000";
					when "10101101100000110" => rgb <= "000000";
					when "10101101100000111" => rgb <= "000000";
					when "10101101100001000" => rgb <= "000000";
					when "10101101100001001" => rgb <= "000000";
					when "10101101100001010" => rgb <= "000000";
					when "10101101100001011" => rgb <= "010101";
					when "10101101100001100" => rgb <= "111111";
					when "10101101100001101" => rgb <= "101010";
					when "10101101100001110" => rgb <= "111111";
					when "10101101100001111" => rgb <= "111111";
					when "10101101100010000" => rgb <= "111111";
					when "10101101100010001" => rgb <= "111111";
					when "10101101100010010" => rgb <= "111111";
					when "10101101100010011" => rgb <= "111111";
					when "10101101100010100" => rgb <= "111111";
					when "10101101100010101" => rgb <= "111111";
					when "10101101100010110" => rgb <= "111111";
					when "10101101100010111" => rgb <= "111111";
					when "10101101100011000" => rgb <= "101010";
					when "10101101100011001" => rgb <= "101010";
					when "10101101100011010" => rgb <= "101010";
					when "10101101100011011" => rgb <= "000000";
					when "10101101100011100" => rgb <= "000000";
					when "10101101100011101" => rgb <= "000000";
					when "10101101100011110" => rgb <= "000000";
					when "10101101100011111" => rgb <= "000000";
					when "10101101100100000" => rgb <= "000000";
					when "10101101100100001" => rgb <= "000000";
					when "10101101100100010" => rgb <= "101010";
					when "10101101100100011" => rgb <= "111111";
					when "10101101100100100" => rgb <= "101010";
					when "10101101100100101" => rgb <= "111111";
					when "10101101100100110" => rgb <= "111111";
					when "10101101100100111" => rgb <= "111111";
					when "10101101100101000" => rgb <= "101010";
					when "10101101100101001" => rgb <= "111111";
					when "10101101100101010" => rgb <= "111111";
					when "10101101100101011" => rgb <= "101010";
					when "10101101100101100" => rgb <= "111111";
					when "10101101100101101" => rgb <= "111111";
					when "10101101100101110" => rgb <= "101010";
					when "10101101100101111" => rgb <= "101010";
					when "10101101100110000" => rgb <= "111111";
					when "10101101100110001" => rgb <= "010101";
					when "10101101100110010" => rgb <= "000000";
					when "10101101100110011" => rgb <= "000000";
					when "10101101100110100" => rgb <= "000000";
					when "10101101100110101" => rgb <= "000000";
					when "10101101100110110" => rgb <= "000000";
					when "10101101100110111" => rgb <= "000000";
					when "10101101100111000" => rgb <= "000000";
					when "10101101100111001" => rgb <= "000000";
					when "10101101100111010" => rgb <= "000000";
					when "10101101100111011" => rgb <= "000000";
					when "10101101100111100" => rgb <= "000000";
					when "10101101100111101" => rgb <= "000000";
					when "10101101100111110" => rgb <= "000000";
					when "10101101100111111" => rgb <= "000000";
					when "10101110000000000" => rgb <= "000000";
					when "10101110000000001" => rgb <= "000000";
					when "10101110000000010" => rgb <= "000000";
					when "10101110000000011" => rgb <= "000000";
					when "10101110000000100" => rgb <= "000000";
					when "10101110000000101" => rgb <= "101010";
					when "10101110000000110" => rgb <= "111111";
					when "10101110000000111" => rgb <= "101010";
					when "10101110000001000" => rgb <= "111111";
					when "10101110000001001" => rgb <= "111111";
					when "10101110000001010" => rgb <= "101010";
					when "10101110000001011" => rgb <= "101010";
					when "10101110000001100" => rgb <= "101010";
					when "10101110000001101" => rgb <= "000000";
					when "10101110000001110" => rgb <= "000000";
					when "10101110000001111" => rgb <= "000000";
					when "10101110000010000" => rgb <= "000000";
					when "10101110000010001" => rgb <= "000000";
					when "10101110000010010" => rgb <= "000000";
					when "10101110000010011" => rgb <= "000000";
					when "10101110000010100" => rgb <= "000000";
					when "10101110000010101" => rgb <= "000000";
					when "10101110000010110" => rgb <= "000000";
					when "10101110000010111" => rgb <= "000000";
					when "10101110000011000" => rgb <= "000000";
					when "10101110000011001" => rgb <= "000000";
					when "10101110000011010" => rgb <= "000000";
					when "10101110000011011" => rgb <= "000000";
					when "10101110000011100" => rgb <= "000000";
					when "10101110000011101" => rgb <= "000000";
					when "10101110000011110" => rgb <= "000000";
					when "10101110000011111" => rgb <= "000000";
					when "10101110000100000" => rgb <= "000000";
					when "10101110000100001" => rgb <= "000000";
					when "10101110000100010" => rgb <= "000000";
					when "10101110000100011" => rgb <= "101010";
					when "10101110000100100" => rgb <= "101010";
					when "10101110000100101" => rgb <= "101010";
					when "10101110000100110" => rgb <= "111111";
					when "10101110000100111" => rgb <= "111111";
					when "10101110000101000" => rgb <= "111111";
					when "10101110000101001" => rgb <= "111111";
					when "10101110000101010" => rgb <= "101010";
					when "10101110000101011" => rgb <= "111111";
					when "10101110000101100" => rgb <= "111111";
					when "10101110000101101" => rgb <= "111111";
					when "10101110000101110" => rgb <= "111111";
					when "10101110000101111" => rgb <= "101010";
					when "10101110000110000" => rgb <= "111111";
					when "10101110000110001" => rgb <= "101010";
					when "10101110000110010" => rgb <= "000000";
					when "10101110000110011" => rgb <= "000000";
					when "10101110000110100" => rgb <= "000000";
					when "10101110000110101" => rgb <= "000000";
					when "10101110000110110" => rgb <= "000000";
					when "10101110000110111" => rgb <= "000000";
					when "10101110000111000" => rgb <= "000000";
					when "10101110000111001" => rgb <= "010101";
					when "10101110000111010" => rgb <= "101010";
					when "10101110000111011" => rgb <= "111111";
					when "10101110000111100" => rgb <= "111111";
					when "10101110000111101" => rgb <= "111111";
					when "10101110000111110" => rgb <= "111111";
					when "10101110000111111" => rgb <= "101010";
					when "10101110001000000" => rgb <= "101010";
					when "10101110001000001" => rgb <= "000000";
					when "10101110001000010" => rgb <= "000000";
					when "10101110001000011" => rgb <= "000000";
					when "10101110001000100" => rgb <= "000000";
					when "10101110001000101" => rgb <= "000000";
					when "10101110001000110" => rgb <= "000000";
					when "10101110001000111" => rgb <= "000000";
					when "10101110001001000" => rgb <= "000000";
					when "10101110001001001" => rgb <= "000000";
					when "10101110001001010" => rgb <= "000000";
					when "10101110001001011" => rgb <= "000000";
					when "10101110001001100" => rgb <= "000000";
					when "10101110001001101" => rgb <= "000000";
					when "10101110001001110" => rgb <= "000000";
					when "10101110001001111" => rgb <= "000000";
					when "10101110001010000" => rgb <= "101010";
					when "10101110001010001" => rgb <= "101010";
					when "10101110001010010" => rgb <= "101010";
					when "10101110001010011" => rgb <= "111111";
					when "10101110001010100" => rgb <= "101010";
					when "10101110001010101" => rgb <= "101010";
					when "10101110001010110" => rgb <= "111111";
					when "10101110001010111" => rgb <= "101010";
					when "10101110001011000" => rgb <= "111111";
					when "10101110001011001" => rgb <= "111111";
					when "10101110001011010" => rgb <= "111111";
					when "10101110001011011" => rgb <= "101010";
					when "10101110001011100" => rgb <= "101010";
					when "10101110001011101" => rgb <= "111111";
					when "10101110001011110" => rgb <= "101010";
					when "10101110001011111" => rgb <= "000000";
					when "10101110001100000" => rgb <= "000000";
					when "10101110001100001" => rgb <= "000000";
					when "10101110001100010" => rgb <= "000000";
					when "10101110001100011" => rgb <= "000000";
					when "10101110001100100" => rgb <= "000000";
					when "10101110001100101" => rgb <= "000000";
					when "10101110001100110" => rgb <= "010101";
					when "10101110001100111" => rgb <= "111111";
					when "10101110001101000" => rgb <= "101010";
					when "10101110001101001" => rgb <= "111111";
					when "10101110001101010" => rgb <= "101010";
					when "10101110001101011" => rgb <= "101010";
					when "10101110001101100" => rgb <= "101010";
					when "10101110001101101" => rgb <= "101010";
					when "10101110001101110" => rgb <= "000000";
					when "10101110001101111" => rgb <= "000000";
					when "10101110001110000" => rgb <= "000000";
					when "10101110001110001" => rgb <= "000000";
					when "10101110001110010" => rgb <= "000000";
					when "10101110001110011" => rgb <= "000000";
					when "10101110001110100" => rgb <= "000000";
					when "10101110001110101" => rgb <= "000000";
					when "10101110001110110" => rgb <= "000000";
					when "10101110001110111" => rgb <= "000000";
					when "10101110001111000" => rgb <= "000000";
					when "10101110001111001" => rgb <= "000000";
					when "10101110001111010" => rgb <= "000000";
					when "10101110001111011" => rgb <= "000000";
					when "10101110001111100" => rgb <= "000000";
					when "10101110001111101" => rgb <= "101010";
					when "10101110001111110" => rgb <= "111111";
					when "10101110001111111" => rgb <= "111111";
					when "10101110010000000" => rgb <= "111111";
					when "10101110010000001" => rgb <= "111111";
					when "10101110010000010" => rgb <= "111111";
					when "10101110010000011" => rgb <= "111111";
					when "10101110010000100" => rgb <= "111111";
					when "10101110010000101" => rgb <= "111111";
					when "10101110010000110" => rgb <= "111111";
					when "10101110010000111" => rgb <= "111111";
					when "10101110010001000" => rgb <= "111111";
					when "10101110010001001" => rgb <= "111111";
					when "10101110010001010" => rgb <= "111111";
					when "10101110010001011" => rgb <= "101010";
					when "10101110010001100" => rgb <= "000000";
					when "10101110010001101" => rgb <= "000000";
					when "10101110010001110" => rgb <= "000000";
					when "10101110010001111" => rgb <= "000000";
					when "10101110010010000" => rgb <= "000000";
					when "10101110010010001" => rgb <= "000000";
					when "10101110010010010" => rgb <= "000000";
					when "10101110010010011" => rgb <= "000000";
					when "10101110010010100" => rgb <= "000000";
					when "10101110010010101" => rgb <= "000000";
					when "10101110010010110" => rgb <= "000000";
					when "10101110010010111" => rgb <= "000000";
					when "10101110010011000" => rgb <= "000000";
					when "10101110010011001" => rgb <= "000000";
					when "10101110010011010" => rgb <= "000000";
					when "10101110010011011" => rgb <= "000000";
					when "10101110010011100" => rgb <= "000000";
					when "10101110010011101" => rgb <= "000000";
					when "10101110010011110" => rgb <= "000000";
					when "10101110010011111" => rgb <= "000000";
					when "10101110010100000" => rgb <= "000000";
					when "10101110010100001" => rgb <= "000000";
					when "10101110010100010" => rgb <= "010101";
					when "10101110010100011" => rgb <= "111111";
					when "10101110010100100" => rgb <= "101010";
					when "10101110010100101" => rgb <= "111111";
					when "10101110010100110" => rgb <= "111111";
					when "10101110010100111" => rgb <= "111111";
					when "10101110010101000" => rgb <= "111111";
					when "10101110010101001" => rgb <= "111111";
					when "10101110010101010" => rgb <= "000000";
					when "10101110010101011" => rgb <= "000000";
					when "10101110010101100" => rgb <= "000000";
					when "10101110010101101" => rgb <= "000000";
					when "10101110010101110" => rgb <= "000000";
					when "10101110010101111" => rgb <= "000000";
					when "10101110010110000" => rgb <= "000000";
					when "10101110010110001" => rgb <= "000000";
					when "10101110010110010" => rgb <= "000000";
					when "10101110010110011" => rgb <= "000000";
					when "10101110010110100" => rgb <= "000000";
					when "10101110010110101" => rgb <= "000000";
					when "10101110010110110" => rgb <= "000000";
					when "10101110010110111" => rgb <= "000000";
					when "10101110010111000" => rgb <= "000000";
					when "10101110010111001" => rgb <= "000000";
					when "10101110010111010" => rgb <= "000000";
					when "10101110010111011" => rgb <= "000000";
					when "10101110010111100" => rgb <= "000000";
					when "10101110010111101" => rgb <= "000000";
					when "10101110010111110" => rgb <= "000000";
					when "10101110010111111" => rgb <= "000000";
					when "10101110011000000" => rgb <= "010101";
					when "10101110011000001" => rgb <= "101010";
					when "10101110011000010" => rgb <= "101010";
					when "10101110011000011" => rgb <= "111111";
					when "10101110011000100" => rgb <= "111111";
					when "10101110011000101" => rgb <= "111111";
					when "10101110011000110" => rgb <= "111111";
					when "10101110011000111" => rgb <= "111111";
					when "10101110011001000" => rgb <= "111111";
					when "10101110011001001" => rgb <= "101010";
					when "10101110011001010" => rgb <= "111111";
					when "10101110011001011" => rgb <= "101010";
					when "10101110011001100" => rgb <= "111111";
					when "10101110011001101" => rgb <= "101010";
					when "10101110011001110" => rgb <= "111111";
					when "10101110011001111" => rgb <= "010101";
					when "10101110011010000" => rgb <= "000000";
					when "10101110011010001" => rgb <= "000000";
					when "10101110011010010" => rgb <= "000000";
					when "10101110011010011" => rgb <= "000000";
					when "10101110011010100" => rgb <= "000000";
					when "10101110011010101" => rgb <= "000000";
					when "10101110011010110" => rgb <= "000000";
					when "10101110011010111" => rgb <= "101010";
					when "10101110011011000" => rgb <= "101010";
					when "10101110011011001" => rgb <= "101010";
					when "10101110011011010" => rgb <= "101010";
					when "10101110011011011" => rgb <= "111111";
					when "10101110011011100" => rgb <= "111111";
					when "10101110011011101" => rgb <= "111111";
					when "10101110011011110" => rgb <= "111111";
					when "10101110011011111" => rgb <= "111111";
					when "10101110011100000" => rgb <= "111111";
					when "10101110011100001" => rgb <= "111111";
					when "10101110011100010" => rgb <= "101010";
					when "10101110011100011" => rgb <= "101010";
					when "10101110011100100" => rgb <= "111111";
					when "10101110011100101" => rgb <= "111111";
					when "10101110011100110" => rgb <= "000000";
					when "10101110011100111" => rgb <= "000000";
					when "10101110011101000" => rgb <= "000000";
					when "10101110011101001" => rgb <= "000000";
					when "10101110011101010" => rgb <= "000000";
					when "10101110011101011" => rgb <= "000000";
					when "10101110011101100" => rgb <= "000000";
					when "10101110011101101" => rgb <= "010101";
					when "10101110011101110" => rgb <= "111111";
					when "10101110011101111" => rgb <= "111111";
					when "10101110011110000" => rgb <= "101010";
					when "10101110011110001" => rgb <= "111111";
					when "10101110011110010" => rgb <= "101010";
					when "10101110011110011" => rgb <= "101010";
					when "10101110011110100" => rgb <= "111111";
					when "10101110011110101" => rgb <= "101010";
					when "10101110011110110" => rgb <= "101010";
					when "10101110011110111" => rgb <= "111111";
					when "10101110011111000" => rgb <= "111111";
					when "10101110011111001" => rgb <= "111111";
					when "10101110011111010" => rgb <= "111111";
					when "10101110011111011" => rgb <= "111111";
					when "10101110011111100" => rgb <= "010101";
					when "10101110011111101" => rgb <= "000000";
					when "10101110011111110" => rgb <= "000000";
					when "10101110011111111" => rgb <= "000000";
					when "10101110100000000" => rgb <= "000000";
					when "10101110100000001" => rgb <= "000000";
					when "10101110100000010" => rgb <= "000000";
					when "10101110100000011" => rgb <= "000000";
					when "10101110100000100" => rgb <= "000000";
					when "10101110100000101" => rgb <= "000000";
					when "10101110100000110" => rgb <= "000000";
					when "10101110100000111" => rgb <= "000000";
					when "10101110100001000" => rgb <= "000000";
					when "10101110100001001" => rgb <= "000000";
					when "10101110100001010" => rgb <= "000000";
					when "10101110100001011" => rgb <= "010101";
					when "10101110100001100" => rgb <= "111111";
					when "10101110100001101" => rgb <= "101010";
					when "10101110100001110" => rgb <= "111111";
					when "10101110100001111" => rgb <= "111111";
					when "10101110100010000" => rgb <= "111111";
					when "10101110100010001" => rgb <= "111111";
					when "10101110100010010" => rgb <= "111111";
					when "10101110100010011" => rgb <= "111111";
					when "10101110100010100" => rgb <= "111111";
					when "10101110100010101" => rgb <= "111111";
					when "10101110100010110" => rgb <= "111111";
					when "10101110100010111" => rgb <= "111111";
					when "10101110100011000" => rgb <= "111111";
					when "10101110100011001" => rgb <= "111111";
					when "10101110100011010" => rgb <= "101010";
					when "10101110100011011" => rgb <= "000000";
					when "10101110100011100" => rgb <= "000000";
					when "10101110100011101" => rgb <= "000000";
					when "10101110100011110" => rgb <= "000000";
					when "10101110100011111" => rgb <= "000000";
					when "10101110100100000" => rgb <= "000000";
					when "10101110100100001" => rgb <= "000000";
					when "10101110100100010" => rgb <= "101010";
					when "10101110100100011" => rgb <= "101010";
					when "10101110100100100" => rgb <= "101010";
					when "10101110100100101" => rgb <= "111111";
					when "10101110100100110" => rgb <= "111111";
					when "10101110100100111" => rgb <= "111111";
					when "10101110100101000" => rgb <= "101010";
					when "10101110100101001" => rgb <= "111111";
					when "10101110100101010" => rgb <= "111111";
					when "10101110100101011" => rgb <= "101010";
					when "10101110100101100" => rgb <= "111111";
					when "10101110100101101" => rgb <= "111111";
					when "10101110100101110" => rgb <= "101010";
					when "10101110100101111" => rgb <= "101010";
					when "10101110100110000" => rgb <= "111111";
					when "10101110100110001" => rgb <= "010101";
					when "10101110100110010" => rgb <= "000000";
					when "10101110100110011" => rgb <= "000000";
					when "10101110100110100" => rgb <= "000000";
					when "10101110100110101" => rgb <= "000000";
					when "10101110100110110" => rgb <= "000000";
					when "10101110100110111" => rgb <= "000000";
					when "10101110100111000" => rgb <= "000000";
					when "10101110100111001" => rgb <= "000000";
					when "10101110100111010" => rgb <= "000000";
					when "10101110100111011" => rgb <= "000000";
					when "10101110100111100" => rgb <= "000000";
					when "10101110100111101" => rgb <= "000000";
					when "10101110100111110" => rgb <= "000000";
					when "10101110100111111" => rgb <= "000000";
					when "10101111000000000" => rgb <= "000000";
					when "10101111000000001" => rgb <= "000000";
					when "10101111000000010" => rgb <= "000000";
					when "10101111000000011" => rgb <= "000000";
					when "10101111000000100" => rgb <= "000000";
					when "10101111000000101" => rgb <= "101010";
					when "10101111000000110" => rgb <= "111111";
					when "10101111000000111" => rgb <= "101010";
					when "10101111000001000" => rgb <= "111111";
					when "10101111000001001" => rgb <= "111111";
					when "10101111000001010" => rgb <= "101010";
					when "10101111000001011" => rgb <= "101010";
					when "10101111000001100" => rgb <= "101010";
					when "10101111000001101" => rgb <= "000000";
					when "10101111000001110" => rgb <= "000000";
					when "10101111000001111" => rgb <= "000000";
					when "10101111000010000" => rgb <= "000000";
					when "10101111000010001" => rgb <= "000000";
					when "10101111000010010" => rgb <= "000000";
					when "10101111000010011" => rgb <= "000000";
					when "10101111000010100" => rgb <= "000000";
					when "10101111000010101" => rgb <= "000000";
					when "10101111000010110" => rgb <= "000000";
					when "10101111000010111" => rgb <= "000000";
					when "10101111000011000" => rgb <= "000000";
					when "10101111000011001" => rgb <= "000000";
					when "10101111000011010" => rgb <= "000000";
					when "10101111000011011" => rgb <= "000000";
					when "10101111000011100" => rgb <= "000000";
					when "10101111000011101" => rgb <= "000000";
					when "10101111000011110" => rgb <= "000000";
					when "10101111000011111" => rgb <= "000000";
					when "10101111000100000" => rgb <= "000000";
					when "10101111000100001" => rgb <= "000000";
					when "10101111000100010" => rgb <= "000000";
					when "10101111000100011" => rgb <= "101010";
					when "10101111000100100" => rgb <= "101010";
					when "10101111000100101" => rgb <= "101010";
					when "10101111000100110" => rgb <= "111111";
					when "10101111000100111" => rgb <= "111111";
					when "10101111000101000" => rgb <= "111111";
					when "10101111000101001" => rgb <= "111111";
					when "10101111000101010" => rgb <= "101010";
					when "10101111000101011" => rgb <= "111111";
					when "10101111000101100" => rgb <= "111111";
					when "10101111000101101" => rgb <= "111111";
					when "10101111000101110" => rgb <= "111111";
					when "10101111000101111" => rgb <= "101010";
					when "10101111000110000" => rgb <= "101010";
					when "10101111000110001" => rgb <= "101010";
					when "10101111000110010" => rgb <= "000000";
					when "10101111000110011" => rgb <= "000000";
					when "10101111000110100" => rgb <= "000000";
					when "10101111000110101" => rgb <= "000000";
					when "10101111000110110" => rgb <= "000000";
					when "10101111000110111" => rgb <= "000000";
					when "10101111000111000" => rgb <= "000000";
					when "10101111000111001" => rgb <= "010101";
					when "10101111000111010" => rgb <= "111111";
					when "10101111000111011" => rgb <= "101010";
					when "10101111000111100" => rgb <= "101010";
					when "10101111000111101" => rgb <= "101010";
					when "10101111000111110" => rgb <= "111111";
					when "10101111000111111" => rgb <= "111111";
					when "10101111001000000" => rgb <= "101010";
					when "10101111001000001" => rgb <= "000000";
					when "10101111001000010" => rgb <= "000000";
					when "10101111001000011" => rgb <= "000000";
					when "10101111001000100" => rgb <= "000000";
					when "10101111001000101" => rgb <= "000000";
					when "10101111001000110" => rgb <= "000000";
					when "10101111001000111" => rgb <= "000000";
					when "10101111001001000" => rgb <= "000000";
					when "10101111001001001" => rgb <= "000000";
					when "10101111001001010" => rgb <= "000000";
					when "10101111001001011" => rgb <= "000000";
					when "10101111001001100" => rgb <= "000000";
					when "10101111001001101" => rgb <= "000000";
					when "10101111001001110" => rgb <= "000000";
					when "10101111001001111" => rgb <= "000000";
					when "10101111001010000" => rgb <= "101010";
					when "10101111001010001" => rgb <= "101010";
					when "10101111001010010" => rgb <= "101010";
					when "10101111001010011" => rgb <= "111111";
					when "10101111001010100" => rgb <= "101010";
					when "10101111001010101" => rgb <= "111111";
					when "10101111001010110" => rgb <= "111111";
					when "10101111001010111" => rgb <= "101010";
					when "10101111001011000" => rgb <= "111111";
					when "10101111001011001" => rgb <= "101010";
					when "10101111001011010" => rgb <= "101010";
					when "10101111001011011" => rgb <= "111111";
					when "10101111001011100" => rgb <= "101010";
					when "10101111001011101" => rgb <= "111111";
					when "10101111001011110" => rgb <= "101010";
					when "10101111001011111" => rgb <= "000000";
					when "10101111001100000" => rgb <= "000000";
					when "10101111001100001" => rgb <= "000000";
					when "10101111001100010" => rgb <= "000000";
					when "10101111001100011" => rgb <= "000000";
					when "10101111001100100" => rgb <= "000000";
					when "10101111001100101" => rgb <= "000000";
					when "10101111001100110" => rgb <= "010101";
					when "10101111001100111" => rgb <= "111111";
					when "10101111001101000" => rgb <= "101010";
					when "10101111001101001" => rgb <= "111111";
					when "10101111001101010" => rgb <= "111111";
					when "10101111001101011" => rgb <= "101010";
					when "10101111001101100" => rgb <= "101010";
					when "10101111001101101" => rgb <= "101010";
					when "10101111001101110" => rgb <= "000000";
					when "10101111001101111" => rgb <= "000000";
					when "10101111001110000" => rgb <= "000000";
					when "10101111001110001" => rgb <= "000000";
					when "10101111001110010" => rgb <= "000000";
					when "10101111001110011" => rgb <= "000000";
					when "10101111001110100" => rgb <= "000000";
					when "10101111001110101" => rgb <= "000000";
					when "10101111001110110" => rgb <= "000000";
					when "10101111001110111" => rgb <= "000000";
					when "10101111001111000" => rgb <= "000000";
					when "10101111001111001" => rgb <= "000000";
					when "10101111001111010" => rgb <= "000000";
					when "10101111001111011" => rgb <= "000000";
					when "10101111001111100" => rgb <= "000000";
					when "10101111001111101" => rgb <= "101010";
					when "10101111001111110" => rgb <= "111111";
					when "10101111001111111" => rgb <= "111111";
					when "10101111010000000" => rgb <= "111111";
					when "10101111010000001" => rgb <= "111111";
					when "10101111010000010" => rgb <= "111111";
					when "10101111010000011" => rgb <= "111111";
					when "10101111010000100" => rgb <= "111111";
					when "10101111010000101" => rgb <= "111111";
					when "10101111010000110" => rgb <= "111111";
					when "10101111010000111" => rgb <= "111111";
					when "10101111010001000" => rgb <= "111111";
					when "10101111010001001" => rgb <= "101010";
					when "10101111010001010" => rgb <= "111111";
					when "10101111010001011" => rgb <= "101010";
					when "10101111010001100" => rgb <= "000000";
					when "10101111010001101" => rgb <= "000000";
					when "10101111010001110" => rgb <= "000000";
					when "10101111010001111" => rgb <= "000000";
					when "10101111010010000" => rgb <= "000000";
					when "10101111010010001" => rgb <= "000000";
					when "10101111010010010" => rgb <= "000000";
					when "10101111010010011" => rgb <= "000000";
					when "10101111010010100" => rgb <= "000000";
					when "10101111010010101" => rgb <= "000000";
					when "10101111010010110" => rgb <= "000000";
					when "10101111010010111" => rgb <= "000000";
					when "10101111010011000" => rgb <= "000000";
					when "10101111010011001" => rgb <= "000000";
					when "10101111010011010" => rgb <= "000000";
					when "10101111010011011" => rgb <= "000000";
					when "10101111010011100" => rgb <= "000000";
					when "10101111010011101" => rgb <= "000000";
					when "10101111010011110" => rgb <= "000000";
					when "10101111010011111" => rgb <= "000000";
					when "10101111010100000" => rgb <= "000000";
					when "10101111010100001" => rgb <= "000000";
					when "10101111010100010" => rgb <= "010101";
					when "10101111010100011" => rgb <= "111111";
					when "10101111010100100" => rgb <= "101010";
					when "10101111010100101" => rgb <= "111111";
					when "10101111010100110" => rgb <= "111111";
					when "10101111010100111" => rgb <= "111111";
					when "10101111010101000" => rgb <= "101010";
					when "10101111010101001" => rgb <= "101010";
					when "10101111010101010" => rgb <= "000000";
					when "10101111010101011" => rgb <= "000000";
					when "10101111010101100" => rgb <= "000000";
					when "10101111010101101" => rgb <= "000000";
					when "10101111010101110" => rgb <= "000000";
					when "10101111010101111" => rgb <= "000000";
					when "10101111010110000" => rgb <= "000000";
					when "10101111010110001" => rgb <= "000000";
					when "10101111010110010" => rgb <= "000000";
					when "10101111010110011" => rgb <= "000000";
					when "10101111010110100" => rgb <= "000000";
					when "10101111010110101" => rgb <= "000000";
					when "10101111010110110" => rgb <= "000000";
					when "10101111010110111" => rgb <= "000000";
					when "10101111010111000" => rgb <= "000000";
					when "10101111010111001" => rgb <= "000000";
					when "10101111010111010" => rgb <= "000000";
					when "10101111010111011" => rgb <= "000000";
					when "10101111010111100" => rgb <= "000000";
					when "10101111010111101" => rgb <= "000000";
					when "10101111010111110" => rgb <= "000000";
					when "10101111010111111" => rgb <= "000000";
					when "10101111011000000" => rgb <= "010101";
					when "10101111011000001" => rgb <= "101010";
					when "10101111011000010" => rgb <= "101010";
					when "10101111011000011" => rgb <= "111111";
					when "10101111011000100" => rgb <= "111111";
					when "10101111011000101" => rgb <= "111111";
					when "10101111011000110" => rgb <= "111111";
					when "10101111011000111" => rgb <= "111111";
					when "10101111011001000" => rgb <= "111111";
					when "10101111011001001" => rgb <= "101010";
					when "10101111011001010" => rgb <= "111111";
					when "10101111011001011" => rgb <= "101010";
					when "10101111011001100" => rgb <= "111111";
					when "10101111011001101" => rgb <= "101010";
					when "10101111011001110" => rgb <= "111111";
					when "10101111011001111" => rgb <= "010101";
					when "10101111011010000" => rgb <= "000000";
					when "10101111011010001" => rgb <= "000000";
					when "10101111011010010" => rgb <= "000000";
					when "10101111011010011" => rgb <= "000000";
					when "10101111011010100" => rgb <= "000000";
					when "10101111011010101" => rgb <= "000000";
					when "10101111011010110" => rgb <= "000000";
					when "10101111011010111" => rgb <= "101010";
					when "10101111011011000" => rgb <= "101010";
					when "10101111011011001" => rgb <= "101010";
					when "10101111011011010" => rgb <= "101010";
					when "10101111011011011" => rgb <= "111111";
					when "10101111011011100" => rgb <= "111111";
					when "10101111011011101" => rgb <= "111111";
					when "10101111011011110" => rgb <= "111111";
					when "10101111011011111" => rgb <= "111111";
					when "10101111011100000" => rgb <= "111111";
					when "10101111011100001" => rgb <= "111111";
					when "10101111011100010" => rgb <= "111111";
					when "10101111011100011" => rgb <= "101010";
					when "10101111011100100" => rgb <= "111111";
					when "10101111011100101" => rgb <= "111111";
					when "10101111011100110" => rgb <= "000000";
					when "10101111011100111" => rgb <= "000000";
					when "10101111011101000" => rgb <= "000000";
					when "10101111011101001" => rgb <= "000000";
					when "10101111011101010" => rgb <= "000000";
					when "10101111011101011" => rgb <= "000000";
					when "10101111011101100" => rgb <= "000000";
					when "10101111011101101" => rgb <= "010101";
					when "10101111011101110" => rgb <= "111111";
					when "10101111011101111" => rgb <= "101010";
					when "10101111011110000" => rgb <= "111111";
					when "10101111011110001" => rgb <= "111111";
					when "10101111011110010" => rgb <= "111111";
					when "10101111011110011" => rgb <= "101010";
					when "10101111011110100" => rgb <= "111111";
					when "10101111011110101" => rgb <= "101010";
					when "10101111011110110" => rgb <= "101010";
					when "10101111011110111" => rgb <= "101010";
					when "10101111011111000" => rgb <= "101010";
					when "10101111011111001" => rgb <= "101010";
					when "10101111011111010" => rgb <= "101010";
					when "10101111011111011" => rgb <= "101010";
					when "10101111011111100" => rgb <= "010101";
					when "10101111011111101" => rgb <= "000000";
					when "10101111011111110" => rgb <= "000000";
					when "10101111011111111" => rgb <= "000000";
					when "10101111100000000" => rgb <= "000000";
					when "10101111100000001" => rgb <= "000000";
					when "10101111100000010" => rgb <= "000000";
					when "10101111100000011" => rgb <= "000000";
					when "10101111100000100" => rgb <= "000000";
					when "10101111100000101" => rgb <= "000000";
					when "10101111100000110" => rgb <= "000000";
					when "10101111100000111" => rgb <= "000000";
					when "10101111100001000" => rgb <= "000000";
					when "10101111100001001" => rgb <= "000000";
					when "10101111100001010" => rgb <= "000000";
					when "10101111100001011" => rgb <= "010101";
					when "10101111100001100" => rgb <= "111111";
					when "10101111100001101" => rgb <= "101010";
					when "10101111100001110" => rgb <= "111111";
					when "10101111100001111" => rgb <= "111111";
					when "10101111100010000" => rgb <= "111111";
					when "10101111100010001" => rgb <= "111111";
					when "10101111100010010" => rgb <= "111111";
					when "10101111100010011" => rgb <= "111111";
					when "10101111100010100" => rgb <= "111111";
					when "10101111100010101" => rgb <= "111111";
					when "10101111100010110" => rgb <= "111111";
					when "10101111100010111" => rgb <= "111111";
					when "10101111100011000" => rgb <= "101010";
					when "10101111100011001" => rgb <= "101010";
					when "10101111100011010" => rgb <= "101010";
					when "10101111100011011" => rgb <= "000000";
					when "10101111100011100" => rgb <= "000000";
					when "10101111100011101" => rgb <= "000000";
					when "10101111100011110" => rgb <= "000000";
					when "10101111100011111" => rgb <= "000000";
					when "10101111100100000" => rgb <= "000000";
					when "10101111100100001" => rgb <= "000000";
					when "10101111100100010" => rgb <= "101010";
					when "10101111100100011" => rgb <= "101010";
					when "10101111100100100" => rgb <= "101010";
					when "10101111100100101" => rgb <= "101010";
					when "10101111100100110" => rgb <= "111111";
					when "10101111100100111" => rgb <= "111111";
					when "10101111100101000" => rgb <= "101010";
					when "10101111100101001" => rgb <= "111111";
					when "10101111100101010" => rgb <= "111111";
					when "10101111100101011" => rgb <= "101010";
					when "10101111100101100" => rgb <= "111111";
					when "10101111100101101" => rgb <= "111111";
					when "10101111100101110" => rgb <= "101010";
					when "10101111100101111" => rgb <= "101010";
					when "10101111100110000" => rgb <= "111111";
					when "10101111100110001" => rgb <= "010101";
					when "10101111100110010" => rgb <= "000000";
					when "10101111100110011" => rgb <= "000000";
					when "10101111100110100" => rgb <= "000000";
					when "10101111100110101" => rgb <= "000000";
					when "10101111100110110" => rgb <= "000000";
					when "10101111100110111" => rgb <= "000000";
					when "10101111100111000" => rgb <= "000000";
					when "10101111100111001" => rgb <= "000000";
					when "10101111100111010" => rgb <= "000000";
					when "10101111100111011" => rgb <= "000000";
					when "10101111100111100" => rgb <= "000000";
					when "10101111100111101" => rgb <= "000000";
					when "10101111100111110" => rgb <= "000000";
					when "10101111100111111" => rgb <= "000000";
					when "10110000000000000" => rgb <= "000000";
					when "10110000000000001" => rgb <= "000000";
					when "10110000000000010" => rgb <= "000000";
					when "10110000000000011" => rgb <= "000000";
					when "10110000000000100" => rgb <= "000000";
					when "10110000000000101" => rgb <= "101010";
					when "10110000000000110" => rgb <= "111111";
					when "10110000000000111" => rgb <= "101010";
					when "10110000000001000" => rgb <= "101010";
					when "10110000000001001" => rgb <= "111111";
					when "10110000000001010" => rgb <= "101010";
					when "10110000000001011" => rgb <= "101010";
					when "10110000000001100" => rgb <= "101010";
					when "10110000000001101" => rgb <= "000000";
					when "10110000000001110" => rgb <= "000000";
					when "10110000000001111" => rgb <= "000000";
					when "10110000000010000" => rgb <= "000000";
					when "10110000000010001" => rgb <= "000000";
					when "10110000000010010" => rgb <= "000000";
					when "10110000000010011" => rgb <= "000000";
					when "10110000000010100" => rgb <= "000000";
					when "10110000000010101" => rgb <= "000000";
					when "10110000000010110" => rgb <= "000000";
					when "10110000000010111" => rgb <= "000000";
					when "10110000000011000" => rgb <= "000000";
					when "10110000000011001" => rgb <= "000000";
					when "10110000000011010" => rgb <= "000000";
					when "10110000000011011" => rgb <= "010101";
					when "10110000000011100" => rgb <= "101010";
					when "10110000000011101" => rgb <= "101010";
					when "10110000000011110" => rgb <= "101010";
					when "10110000000011111" => rgb <= "101010";
					when "10110000000100000" => rgb <= "101010";
					when "10110000000100001" => rgb <= "101010";
					when "10110000000100010" => rgb <= "101010";
					when "10110000000100011" => rgb <= "101010";
					when "10110000000100100" => rgb <= "101010";
					when "10110000000100101" => rgb <= "101010";
					when "10110000000100110" => rgb <= "111111";
					when "10110000000100111" => rgb <= "111111";
					when "10110000000101000" => rgb <= "111111";
					when "10110000000101001" => rgb <= "101010";
					when "10110000000101010" => rgb <= "101010";
					when "10110000000101011" => rgb <= "111111";
					when "10110000000101100" => rgb <= "101010";
					when "10110000000101101" => rgb <= "111111";
					when "10110000000101110" => rgb <= "111111";
					when "10110000000101111" => rgb <= "111111";
					when "10110000000110000" => rgb <= "101010";
					when "10110000000110001" => rgb <= "101010";
					when "10110000000110010" => rgb <= "000000";
					when "10110000000110011" => rgb <= "000000";
					when "10110000000110100" => rgb <= "000000";
					when "10110000000110101" => rgb <= "000000";
					when "10110000000110110" => rgb <= "000000";
					when "10110000000110111" => rgb <= "000000";
					when "10110000000111000" => rgb <= "000000";
					when "10110000000111001" => rgb <= "010101";
					when "10110000000111010" => rgb <= "111111";
					when "10110000000111011" => rgb <= "101010";
					when "10110000000111100" => rgb <= "101010";
					when "10110000000111101" => rgb <= "111111";
					when "10110000000111110" => rgb <= "101010";
					when "10110000000111111" => rgb <= "111111";
					when "10110000001000000" => rgb <= "101010";
					when "10110000001000001" => rgb <= "000000";
					when "10110000001000010" => rgb <= "000000";
					when "10110000001000011" => rgb <= "000000";
					when "10110000001000100" => rgb <= "000000";
					when "10110000001000101" => rgb <= "000000";
					when "10110000001000110" => rgb <= "000000";
					when "10110000001000111" => rgb <= "000000";
					when "10110000001001000" => rgb <= "000000";
					when "10110000001001001" => rgb <= "000000";
					when "10110000001001010" => rgb <= "000000";
					when "10110000001001011" => rgb <= "000000";
					when "10110000001001100" => rgb <= "000000";
					when "10110000001001101" => rgb <= "000000";
					when "10110000001001110" => rgb <= "000000";
					when "10110000001001111" => rgb <= "000000";
					when "10110000001010000" => rgb <= "101010";
					when "10110000001010001" => rgb <= "101010";
					when "10110000001010010" => rgb <= "101010";
					when "10110000001010011" => rgb <= "101010";
					when "10110000001010100" => rgb <= "111111";
					when "10110000001010101" => rgb <= "111111";
					when "10110000001010110" => rgb <= "111111";
					when "10110000001010111" => rgb <= "111111";
					when "10110000001011000" => rgb <= "111111";
					when "10110000001011001" => rgb <= "111111";
					when "10110000001011010" => rgb <= "111111";
					when "10110000001011011" => rgb <= "101010";
					when "10110000001011100" => rgb <= "111111";
					when "10110000001011101" => rgb <= "101010";
					when "10110000001011110" => rgb <= "101010";
					when "10110000001011111" => rgb <= "000000";
					when "10110000001100000" => rgb <= "000000";
					when "10110000001100001" => rgb <= "000000";
					when "10110000001100010" => rgb <= "000000";
					when "10110000001100011" => rgb <= "000000";
					when "10110000001100100" => rgb <= "000000";
					when "10110000001100101" => rgb <= "000000";
					when "10110000001100110" => rgb <= "010101";
					when "10110000001100111" => rgb <= "101010";
					when "10110000001101000" => rgb <= "101010";
					when "10110000001101001" => rgb <= "111111";
					when "10110000001101010" => rgb <= "101010";
					when "10110000001101011" => rgb <= "111111";
					when "10110000001101100" => rgb <= "101010";
					when "10110000001101101" => rgb <= "101010";
					when "10110000001101110" => rgb <= "000000";
					when "10110000001101111" => rgb <= "000000";
					when "10110000001110000" => rgb <= "000000";
					when "10110000001110001" => rgb <= "000000";
					when "10110000001110010" => rgb <= "000000";
					when "10110000001110011" => rgb <= "000000";
					when "10110000001110100" => rgb <= "000000";
					when "10110000001110101" => rgb <= "000000";
					when "10110000001110110" => rgb <= "000000";
					when "10110000001110111" => rgb <= "000000";
					when "10110000001111000" => rgb <= "000000";
					when "10110000001111001" => rgb <= "000000";
					when "10110000001111010" => rgb <= "000000";
					when "10110000001111011" => rgb <= "000000";
					when "10110000001111100" => rgb <= "000000";
					when "10110000001111101" => rgb <= "101010";
					when "10110000001111110" => rgb <= "111111";
					when "10110000001111111" => rgb <= "111111";
					when "10110000010000000" => rgb <= "111111";
					when "10110000010000001" => rgb <= "111111";
					when "10110000010000010" => rgb <= "111111";
					when "10110000010000011" => rgb <= "111111";
					when "10110000010000100" => rgb <= "111111";
					when "10110000010000101" => rgb <= "111111";
					when "10110000010000110" => rgb <= "111111";
					when "10110000010000111" => rgb <= "111111";
					when "10110000010001000" => rgb <= "111111";
					when "10110000010001001" => rgb <= "111111";
					when "10110000010001010" => rgb <= "111111";
					when "10110000010001011" => rgb <= "101010";
					when "10110000010001100" => rgb <= "000000";
					when "10110000010001101" => rgb <= "000000";
					when "10110000010001110" => rgb <= "000000";
					when "10110000010001111" => rgb <= "000000";
					when "10110000010010000" => rgb <= "000000";
					when "10110000010010001" => rgb <= "000000";
					when "10110000010010010" => rgb <= "000000";
					when "10110000010010011" => rgb <= "000000";
					when "10110000010010100" => rgb <= "000000";
					when "10110000010010101" => rgb <= "000000";
					when "10110000010010110" => rgb <= "000000";
					when "10110000010010111" => rgb <= "000000";
					when "10110000010011000" => rgb <= "000000";
					when "10110000010011001" => rgb <= "000000";
					when "10110000010011010" => rgb <= "000000";
					when "10110000010011011" => rgb <= "000000";
					when "10110000010011100" => rgb <= "000000";
					when "10110000010011101" => rgb <= "000000";
					when "10110000010011110" => rgb <= "000000";
					when "10110000010011111" => rgb <= "000000";
					when "10110000010100000" => rgb <= "000000";
					when "10110000010100001" => rgb <= "000000";
					when "10110000010100010" => rgb <= "010101";
					when "10110000010100011" => rgb <= "111111";
					when "10110000010100100" => rgb <= "101010";
					when "10110000010100101" => rgb <= "111111";
					when "10110000010100110" => rgb <= "111111";
					when "10110000010100111" => rgb <= "111111";
					when "10110000010101000" => rgb <= "111111";
					when "10110000010101001" => rgb <= "111111";
					when "10110000010101010" => rgb <= "000000";
					when "10110000010101011" => rgb <= "000000";
					when "10110000010101100" => rgb <= "000000";
					when "10110000010101101" => rgb <= "000000";
					when "10110000010101110" => rgb <= "000000";
					when "10110000010101111" => rgb <= "000000";
					when "10110000010110000" => rgb <= "000000";
					when "10110000010110001" => rgb <= "000000";
					when "10110000010110010" => rgb <= "000000";
					when "10110000010110011" => rgb <= "000000";
					when "10110000010110100" => rgb <= "000000";
					when "10110000010110101" => rgb <= "000000";
					when "10110000010110110" => rgb <= "000000";
					when "10110000010110111" => rgb <= "000000";
					when "10110000010111000" => rgb <= "000000";
					when "10110000010111001" => rgb <= "000000";
					when "10110000010111010" => rgb <= "000000";
					when "10110000010111011" => rgb <= "000000";
					when "10110000010111100" => rgb <= "000000";
					when "10110000010111101" => rgb <= "000000";
					when "10110000010111110" => rgb <= "000000";
					when "10110000010111111" => rgb <= "000000";
					when "10110000011000000" => rgb <= "010101";
					when "10110000011000001" => rgb <= "101010";
					when "10110000011000010" => rgb <= "101010";
					when "10110000011000011" => rgb <= "111111";
					when "10110000011000100" => rgb <= "111111";
					when "10110000011000101" => rgb <= "111111";
					when "10110000011000110" => rgb <= "111111";
					when "10110000011000111" => rgb <= "111111";
					when "10110000011001000" => rgb <= "111111";
					when "10110000011001001" => rgb <= "111111";
					when "10110000011001010" => rgb <= "111111";
					when "10110000011001011" => rgb <= "101010";
					when "10110000011001100" => rgb <= "111111";
					when "10110000011001101" => rgb <= "101010";
					when "10110000011001110" => rgb <= "111111";
					when "10110000011001111" => rgb <= "101010";
					when "10110000011010000" => rgb <= "000000";
					when "10110000011010001" => rgb <= "000000";
					when "10110000011010010" => rgb <= "000000";
					when "10110000011010011" => rgb <= "000000";
					when "10110000011010100" => rgb <= "000000";
					when "10110000011010101" => rgb <= "000000";
					when "10110000011010110" => rgb <= "000000";
					when "10110000011010111" => rgb <= "101010";
					when "10110000011011000" => rgb <= "101010";
					when "10110000011011001" => rgb <= "101010";
					when "10110000011011010" => rgb <= "101010";
					when "10110000011011011" => rgb <= "111111";
					when "10110000011011100" => rgb <= "111111";
					when "10110000011011101" => rgb <= "111111";
					when "10110000011011110" => rgb <= "111111";
					when "10110000011011111" => rgb <= "111111";
					when "10110000011100000" => rgb <= "111111";
					when "10110000011100001" => rgb <= "111111";
					when "10110000011100010" => rgb <= "111111";
					when "10110000011100011" => rgb <= "101010";
					when "10110000011100100" => rgb <= "111111";
					when "10110000011100101" => rgb <= "111111";
					when "10110000011100110" => rgb <= "000000";
					when "10110000011100111" => rgb <= "000000";
					when "10110000011101000" => rgb <= "000000";
					when "10110000011101001" => rgb <= "000000";
					when "10110000011101010" => rgb <= "000000";
					when "10110000011101011" => rgb <= "000000";
					when "10110000011101100" => rgb <= "000000";
					when "10110000011101101" => rgb <= "010101";
					when "10110000011101110" => rgb <= "111111";
					when "10110000011101111" => rgb <= "101010";
					when "10110000011110000" => rgb <= "111111";
					when "10110000011110001" => rgb <= "111111";
					when "10110000011110010" => rgb <= "101010";
					when "10110000011110011" => rgb <= "111111";
					when "10110000011110100" => rgb <= "101010";
					when "10110000011110101" => rgb <= "000000";
					when "10110000011110110" => rgb <= "000000";
					when "10110000011110111" => rgb <= "000000";
					when "10110000011111000" => rgb <= "000000";
					when "10110000011111001" => rgb <= "000000";
					when "10110000011111010" => rgb <= "000000";
					when "10110000011111011" => rgb <= "000000";
					when "10110000011111100" => rgb <= "010101";
					when "10110000011111101" => rgb <= "101010";
					when "10110000011111110" => rgb <= "101010";
					when "10110000011111111" => rgb <= "101010";
					when "10110000100000000" => rgb <= "101010";
					when "10110000100000001" => rgb <= "101010";
					when "10110000100000010" => rgb <= "101010";
					when "10110000100000011" => rgb <= "101010";
					when "10110000100000100" => rgb <= "000000";
					when "10110000100000101" => rgb <= "000000";
					when "10110000100000110" => rgb <= "000000";
					when "10110000100000111" => rgb <= "000000";
					when "10110000100001000" => rgb <= "000000";
					when "10110000100001001" => rgb <= "000000";
					when "10110000100001010" => rgb <= "000000";
					when "10110000100001011" => rgb <= "010101";
					when "10110000100001100" => rgb <= "111111";
					when "10110000100001101" => rgb <= "101010";
					when "10110000100001110" => rgb <= "111111";
					when "10110000100001111" => rgb <= "101010";
					when "10110000100010000" => rgb <= "111111";
					when "10110000100010001" => rgb <= "111111";
					when "10110000100010010" => rgb <= "111111";
					when "10110000100010011" => rgb <= "111111";
					when "10110000100010100" => rgb <= "111111";
					when "10110000100010101" => rgb <= "111111";
					when "10110000100010110" => rgb <= "111111";
					when "10110000100010111" => rgb <= "111111";
					when "10110000100011000" => rgb <= "101010";
					when "10110000100011001" => rgb <= "111111";
					when "10110000100011010" => rgb <= "101010";
					when "10110000100011011" => rgb <= "000000";
					when "10110000100011100" => rgb <= "000000";
					when "10110000100011101" => rgb <= "000000";
					when "10110000100011110" => rgb <= "000000";
					when "10110000100011111" => rgb <= "000000";
					when "10110000100100000" => rgb <= "000000";
					when "10110000100100001" => rgb <= "000000";
					when "10110000100100010" => rgb <= "101010";
					when "10110000100100011" => rgb <= "101010";
					when "10110000100100100" => rgb <= "101010";
					when "10110000100100101" => rgb <= "111111";
					when "10110000100100110" => rgb <= "111111";
					when "10110000100100111" => rgb <= "111111";
					when "10110000100101000" => rgb <= "111111";
					when "10110000100101001" => rgb <= "111111";
					when "10110000100101010" => rgb <= "111111";
					when "10110000100101011" => rgb <= "111111";
					when "10110000100101100" => rgb <= "111111";
					when "10110000100101101" => rgb <= "111111";
					when "10110000100101110" => rgb <= "101010";
					when "10110000100101111" => rgb <= "101010";
					when "10110000100110000" => rgb <= "111111";
					when "10110000100110001" => rgb <= "010101";
					when "10110000100110010" => rgb <= "000000";
					when "10110000100110011" => rgb <= "000000";
					when "10110000100110100" => rgb <= "000000";
					when "10110000100110101" => rgb <= "000000";
					when "10110000100110110" => rgb <= "000000";
					when "10110000100110111" => rgb <= "000000";
					when "10110000100111000" => rgb <= "000000";
					when "10110000100111001" => rgb <= "000000";
					when "10110000100111010" => rgb <= "000000";
					when "10110000100111011" => rgb <= "000000";
					when "10110000100111100" => rgb <= "000000";
					when "10110000100111101" => rgb <= "000000";
					when "10110000100111110" => rgb <= "000000";
					when "10110000100111111" => rgb <= "000000";
					when "10110001000000000" => rgb <= "000000";
					when "10110001000000001" => rgb <= "000000";
					when "10110001000000010" => rgb <= "000000";
					when "10110001000000011" => rgb <= "000000";
					when "10110001000000100" => rgb <= "000000";
					when "10110001000000101" => rgb <= "101010";
					when "10110001000000110" => rgb <= "111111";
					when "10110001000000111" => rgb <= "111111";
					when "10110001000001000" => rgb <= "111111";
					when "10110001000001001" => rgb <= "101010";
					when "10110001000001010" => rgb <= "101010";
					when "10110001000001011" => rgb <= "111111";
					when "10110001000001100" => rgb <= "010101";
					when "10110001000001101" => rgb <= "000000";
					when "10110001000001110" => rgb <= "000000";
					when "10110001000001111" => rgb <= "000000";
					when "10110001000010000" => rgb <= "000000";
					when "10110001000010001" => rgb <= "000000";
					when "10110001000010010" => rgb <= "000000";
					when "10110001000010011" => rgb <= "000000";
					when "10110001000010100" => rgb <= "000000";
					when "10110001000010101" => rgb <= "000000";
					when "10110001000010110" => rgb <= "000000";
					when "10110001000010111" => rgb <= "000000";
					when "10110001000011000" => rgb <= "000000";
					when "10110001000011001" => rgb <= "000000";
					when "10110001000011010" => rgb <= "000000";
					when "10110001000011011" => rgb <= "010101";
					when "10110001000011100" => rgb <= "111111";
					when "10110001000011101" => rgb <= "101010";
					when "10110001000011110" => rgb <= "111111";
					when "10110001000011111" => rgb <= "101010";
					when "10110001000100000" => rgb <= "101010";
					when "10110001000100001" => rgb <= "101010";
					when "10110001000100010" => rgb <= "101010";
					when "10110001000100011" => rgb <= "101010";
					when "10110001000100100" => rgb <= "111111";
					when "10110001000100101" => rgb <= "111111";
					when "10110001000100110" => rgb <= "111111";
					when "10110001000100111" => rgb <= "111111";
					when "10110001000101000" => rgb <= "101010";
					when "10110001000101001" => rgb <= "111111";
					when "10110001000101010" => rgb <= "111111";
					when "10110001000101011" => rgb <= "101010";
					when "10110001000101100" => rgb <= "111111";
					when "10110001000101101" => rgb <= "111111";
					when "10110001000101110" => rgb <= "101010";
					when "10110001000101111" => rgb <= "101010";
					when "10110001000110000" => rgb <= "101010";
					when "10110001000110001" => rgb <= "101010";
					when "10110001000110010" => rgb <= "000000";
					when "10110001000110011" => rgb <= "000000";
					when "10110001000110100" => rgb <= "000000";
					when "10110001000110101" => rgb <= "000000";
					when "10110001000110110" => rgb <= "000000";
					when "10110001000110111" => rgb <= "000000";
					when "10110001000111000" => rgb <= "000000";
					when "10110001000111001" => rgb <= "010101";
					when "10110001000111010" => rgb <= "111111";
					when "10110001000111011" => rgb <= "101010";
					when "10110001000111100" => rgb <= "101010";
					when "10110001000111101" => rgb <= "111111";
					when "10110001000111110" => rgb <= "101010";
					when "10110001000111111" => rgb <= "111111";
					when "10110001001000000" => rgb <= "101010";
					when "10110001001000001" => rgb <= "000000";
					when "10110001001000010" => rgb <= "000000";
					when "10110001001000011" => rgb <= "000000";
					when "10110001001000100" => rgb <= "000000";
					when "10110001001000101" => rgb <= "000000";
					when "10110001001000110" => rgb <= "000000";
					when "10110001001000111" => rgb <= "000000";
					when "10110001001001000" => rgb <= "000000";
					when "10110001001001001" => rgb <= "000000";
					when "10110001001001010" => rgb <= "000000";
					when "10110001001001011" => rgb <= "000000";
					when "10110001001001100" => rgb <= "000000";
					when "10110001001001101" => rgb <= "000000";
					when "10110001001001110" => rgb <= "000000";
					when "10110001001001111" => rgb <= "000000";
					when "10110001001010000" => rgb <= "101010";
					when "10110001001010001" => rgb <= "101010";
					when "10110001001010010" => rgb <= "101010";
					when "10110001001010011" => rgb <= "101010";
					when "10110001001010100" => rgb <= "111111";
					when "10110001001010101" => rgb <= "111111";
					when "10110001001010110" => rgb <= "111111";
					when "10110001001010111" => rgb <= "111111";
					when "10110001001011000" => rgb <= "111111";
					when "10110001001011001" => rgb <= "111111";
					when "10110001001011010" => rgb <= "111111";
					when "10110001001011011" => rgb <= "101010";
					when "10110001001011100" => rgb <= "111111";
					when "10110001001011101" => rgb <= "101010";
					when "10110001001011110" => rgb <= "101010";
					when "10110001001011111" => rgb <= "000000";
					when "10110001001100000" => rgb <= "000000";
					when "10110001001100001" => rgb <= "000000";
					when "10110001001100010" => rgb <= "000000";
					when "10110001001100011" => rgb <= "000000";
					when "10110001001100100" => rgb <= "000000";
					when "10110001001100101" => rgb <= "000000";
					when "10110001001100110" => rgb <= "010101";
					when "10110001001100111" => rgb <= "111111";
					when "10110001001101000" => rgb <= "101010";
					when "10110001001101001" => rgb <= "111111";
					when "10110001001101010" => rgb <= "101010";
					when "10110001001101011" => rgb <= "111111";
					when "10110001001101100" => rgb <= "101010";
					when "10110001001101101" => rgb <= "101010";
					when "10110001001101110" => rgb <= "000000";
					when "10110001001101111" => rgb <= "000000";
					when "10110001001110000" => rgb <= "000000";
					when "10110001001110001" => rgb <= "000000";
					when "10110001001110010" => rgb <= "000000";
					when "10110001001110011" => rgb <= "000000";
					when "10110001001110100" => rgb <= "000000";
					when "10110001001110101" => rgb <= "000000";
					when "10110001001110110" => rgb <= "000000";
					when "10110001001110111" => rgb <= "000000";
					when "10110001001111000" => rgb <= "000000";
					when "10110001001111001" => rgb <= "000000";
					when "10110001001111010" => rgb <= "000000";
					when "10110001001111011" => rgb <= "000000";
					when "10110001001111100" => rgb <= "000000";
					when "10110001001111101" => rgb <= "101010";
					when "10110001001111110" => rgb <= "111111";
					when "10110001001111111" => rgb <= "111111";
					when "10110001010000000" => rgb <= "111111";
					when "10110001010000001" => rgb <= "111111";
					when "10110001010000010" => rgb <= "111111";
					when "10110001010000011" => rgb <= "111111";
					when "10110001010000100" => rgb <= "111111";
					when "10110001010000101" => rgb <= "111111";
					when "10110001010000110" => rgb <= "111111";
					when "10110001010000111" => rgb <= "111111";
					when "10110001010001000" => rgb <= "111111";
					when "10110001010001001" => rgb <= "111111";
					when "10110001010001010" => rgb <= "111111";
					when "10110001010001011" => rgb <= "101010";
					when "10110001010001100" => rgb <= "000000";
					when "10110001010001101" => rgb <= "000000";
					when "10110001010001110" => rgb <= "000000";
					when "10110001010001111" => rgb <= "000000";
					when "10110001010010000" => rgb <= "000000";
					when "10110001010010001" => rgb <= "000000";
					when "10110001010010010" => rgb <= "000000";
					when "10110001010010011" => rgb <= "000000";
					when "10110001010010100" => rgb <= "000000";
					when "10110001010010101" => rgb <= "000000";
					when "10110001010010110" => rgb <= "000000";
					when "10110001010010111" => rgb <= "000000";
					when "10110001010011000" => rgb <= "000000";
					when "10110001010011001" => rgb <= "000000";
					when "10110001010011010" => rgb <= "000000";
					when "10110001010011011" => rgb <= "000000";
					when "10110001010011100" => rgb <= "000000";
					when "10110001010011101" => rgb <= "000000";
					when "10110001010011110" => rgb <= "000000";
					when "10110001010011111" => rgb <= "000000";
					when "10110001010100000" => rgb <= "000000";
					when "10110001010100001" => rgb <= "000000";
					when "10110001010100010" => rgb <= "010101";
					when "10110001010100011" => rgb <= "111111";
					when "10110001010100100" => rgb <= "101010";
					when "10110001010100101" => rgb <= "111111";
					when "10110001010100110" => rgb <= "111111";
					when "10110001010100111" => rgb <= "111111";
					when "10110001010101000" => rgb <= "111111";
					when "10110001010101001" => rgb <= "111111";
					when "10110001010101010" => rgb <= "000000";
					when "10110001010101011" => rgb <= "000000";
					when "10110001010101100" => rgb <= "000000";
					when "10110001010101101" => rgb <= "000000";
					when "10110001010101110" => rgb <= "000000";
					when "10110001010101111" => rgb <= "000000";
					when "10110001010110000" => rgb <= "000000";
					when "10110001010110001" => rgb <= "000000";
					when "10110001010110010" => rgb <= "000000";
					when "10110001010110011" => rgb <= "000000";
					when "10110001010110100" => rgb <= "000000";
					when "10110001010110101" => rgb <= "000000";
					when "10110001010110110" => rgb <= "000000";
					when "10110001010110111" => rgb <= "000000";
					when "10110001010111000" => rgb <= "000000";
					when "10110001010111001" => rgb <= "000000";
					when "10110001010111010" => rgb <= "000000";
					when "10110001010111011" => rgb <= "000000";
					when "10110001010111100" => rgb <= "000000";
					when "10110001010111101" => rgb <= "000000";
					when "10110001010111110" => rgb <= "000000";
					when "10110001010111111" => rgb <= "000000";
					when "10110001011000000" => rgb <= "010101";
					when "10110001011000001" => rgb <= "101010";
					when "10110001011000010" => rgb <= "101010";
					when "10110001011000011" => rgb <= "111111";
					when "10110001011000100" => rgb <= "111111";
					when "10110001011000101" => rgb <= "111111";
					when "10110001011000110" => rgb <= "111111";
					when "10110001011000111" => rgb <= "111111";
					when "10110001011001000" => rgb <= "111111";
					when "10110001011001001" => rgb <= "111111";
					when "10110001011001010" => rgb <= "111111";
					when "10110001011001011" => rgb <= "101010";
					when "10110001011001100" => rgb <= "111111";
					when "10110001011001101" => rgb <= "101010";
					when "10110001011001110" => rgb <= "111111";
					when "10110001011001111" => rgb <= "101010";
					when "10110001011010000" => rgb <= "000000";
					when "10110001011010001" => rgb <= "000000";
					when "10110001011010010" => rgb <= "000000";
					when "10110001011010011" => rgb <= "000000";
					when "10110001011010100" => rgb <= "000000";
					when "10110001011010101" => rgb <= "000000";
					when "10110001011010110" => rgb <= "000000";
					when "10110001011010111" => rgb <= "101010";
					when "10110001011011000" => rgb <= "101010";
					when "10110001011011001" => rgb <= "101010";
					when "10110001011011010" => rgb <= "101010";
					when "10110001011011011" => rgb <= "111111";
					when "10110001011011100" => rgb <= "111111";
					when "10110001011011101" => rgb <= "111111";
					when "10110001011011110" => rgb <= "111111";
					when "10110001011011111" => rgb <= "111111";
					when "10110001011100000" => rgb <= "111111";
					when "10110001011100001" => rgb <= "111111";
					when "10110001011100010" => rgb <= "111111";
					when "10110001011100011" => rgb <= "101010";
					when "10110001011100100" => rgb <= "111111";
					when "10110001011100101" => rgb <= "111111";
					when "10110001011100110" => rgb <= "000000";
					when "10110001011100111" => rgb <= "000000";
					when "10110001011101000" => rgb <= "000000";
					when "10110001011101001" => rgb <= "000000";
					when "10110001011101010" => rgb <= "000000";
					when "10110001011101011" => rgb <= "000000";
					when "10110001011101100" => rgb <= "000000";
					when "10110001011101101" => rgb <= "010101";
					when "10110001011101110" => rgb <= "111111";
					when "10110001011101111" => rgb <= "101010";
					when "10110001011110000" => rgb <= "111111";
					when "10110001011110001" => rgb <= "111111";
					when "10110001011110010" => rgb <= "101010";
					when "10110001011110011" => rgb <= "101010";
					when "10110001011110100" => rgb <= "101010";
					when "10110001011110101" => rgb <= "000000";
					when "10110001011110110" => rgb <= "000000";
					when "10110001011110111" => rgb <= "000000";
					when "10110001011111000" => rgb <= "000000";
					when "10110001011111001" => rgb <= "000000";
					when "10110001011111010" => rgb <= "000000";
					when "10110001011111011" => rgb <= "000000";
					when "10110001011111100" => rgb <= "010101";
					when "10110001011111101" => rgb <= "101010";
					when "10110001011111110" => rgb <= "111111";
					when "10110001011111111" => rgb <= "111111";
					when "10110001100000000" => rgb <= "111111";
					when "10110001100000001" => rgb <= "111111";
					when "10110001100000010" => rgb <= "101010";
					when "10110001100000011" => rgb <= "111111";
					when "10110001100000100" => rgb <= "000000";
					when "10110001100000101" => rgb <= "000000";
					when "10110001100000110" => rgb <= "000000";
					when "10110001100000111" => rgb <= "000000";
					when "10110001100001000" => rgb <= "000000";
					when "10110001100001001" => rgb <= "000000";
					when "10110001100001010" => rgb <= "000000";
					when "10110001100001011" => rgb <= "010101";
					when "10110001100001100" => rgb <= "111111";
					when "10110001100001101" => rgb <= "101010";
					when "10110001100001110" => rgb <= "111111";
					when "10110001100001111" => rgb <= "111111";
					when "10110001100010000" => rgb <= "111111";
					when "10110001100010001" => rgb <= "111111";
					when "10110001100010010" => rgb <= "111111";
					when "10110001100010011" => rgb <= "111111";
					when "10110001100010100" => rgb <= "111111";
					when "10110001100010101" => rgb <= "111111";
					when "10110001100010110" => rgb <= "111111";
					when "10110001100010111" => rgb <= "111111";
					when "10110001100011000" => rgb <= "101010";
					when "10110001100011001" => rgb <= "111111";
					when "10110001100011010" => rgb <= "101010";
					when "10110001100011011" => rgb <= "000000";
					when "10110001100011100" => rgb <= "000000";
					when "10110001100011101" => rgb <= "000000";
					when "10110001100011110" => rgb <= "000000";
					when "10110001100011111" => rgb <= "000000";
					when "10110001100100000" => rgb <= "000000";
					when "10110001100100001" => rgb <= "000000";
					when "10110001100100010" => rgb <= "101010";
					when "10110001100100011" => rgb <= "101010";
					when "10110001100100100" => rgb <= "101010";
					when "10110001100100101" => rgb <= "111111";
					when "10110001100100110" => rgb <= "111111";
					when "10110001100100111" => rgb <= "111111";
					when "10110001100101000" => rgb <= "111111";
					when "10110001100101001" => rgb <= "111111";
					when "10110001100101010" => rgb <= "111111";
					when "10110001100101011" => rgb <= "111111";
					when "10110001100101100" => rgb <= "111111";
					when "10110001100101101" => rgb <= "111111";
					when "10110001100101110" => rgb <= "101010";
					when "10110001100101111" => rgb <= "101010";
					when "10110001100110000" => rgb <= "111111";
					when "10110001100110001" => rgb <= "010101";
					when "10110001100110010" => rgb <= "000000";
					when "10110001100110011" => rgb <= "000000";
					when "10110001100110100" => rgb <= "000000";
					when "10110001100110101" => rgb <= "000000";
					when "10110001100110110" => rgb <= "000000";
					when "10110001100110111" => rgb <= "000000";
					when "10110001100111000" => rgb <= "000000";
					when "10110001100111001" => rgb <= "000000";
					when "10110001100111010" => rgb <= "000000";
					when "10110001100111011" => rgb <= "000000";
					when "10110001100111100" => rgb <= "000000";
					when "10110001100111101" => rgb <= "000000";
					when "10110001100111110" => rgb <= "000000";
					when "10110001100111111" => rgb <= "000000";
					when "10110010000000000" => rgb <= "000000";
					when "10110010000000001" => rgb <= "000000";
					when "10110010000000010" => rgb <= "000000";
					when "10110010000000011" => rgb <= "000000";
					when "10110010000000100" => rgb <= "000000";
					when "10110010000000101" => rgb <= "101010";
					when "10110010000000110" => rgb <= "101010";
					when "10110010000000111" => rgb <= "101010";
					when "10110010000001000" => rgb <= "101010";
					when "10110010000001001" => rgb <= "101010";
					when "10110010000001010" => rgb <= "101010";
					when "10110010000001011" => rgb <= "111111";
					when "10110010000001100" => rgb <= "010101";
					when "10110010000001101" => rgb <= "000000";
					when "10110010000001110" => rgb <= "000000";
					when "10110010000001111" => rgb <= "000000";
					when "10110010000010000" => rgb <= "000000";
					when "10110010000010001" => rgb <= "000000";
					when "10110010000010010" => rgb <= "000000";
					when "10110010000010011" => rgb <= "000000";
					when "10110010000010100" => rgb <= "000000";
					when "10110010000010101" => rgb <= "000000";
					when "10110010000010110" => rgb <= "000000";
					when "10110010000010111" => rgb <= "000000";
					when "10110010000011000" => rgb <= "000000";
					when "10110010000011001" => rgb <= "000000";
					when "10110010000011010" => rgb <= "000000";
					when "10110010000011011" => rgb <= "010101";
					when "10110010000011100" => rgb <= "111111";
					when "10110010000011101" => rgb <= "101010";
					when "10110010000011110" => rgb <= "101010";
					when "10110010000011111" => rgb <= "111111";
					when "10110010000100000" => rgb <= "111111";
					when "10110010000100001" => rgb <= "101010";
					when "10110010000100010" => rgb <= "101010";
					when "10110010000100011" => rgb <= "111111";
					when "10110010000100100" => rgb <= "111111";
					when "10110010000100101" => rgb <= "111111";
					when "10110010000100110" => rgb <= "111111";
					when "10110010000100111" => rgb <= "101010";
					when "10110010000101000" => rgb <= "111111";
					when "10110010000101001" => rgb <= "101010";
					when "10110010000101010" => rgb <= "101010";
					when "10110010000101011" => rgb <= "101010";
					when "10110010000101100" => rgb <= "111111";
					when "10110010000101101" => rgb <= "101010";
					when "10110010000101110" => rgb <= "101010";
					when "10110010000101111" => rgb <= "111111";
					when "10110010000110000" => rgb <= "111111";
					when "10110010000110001" => rgb <= "101010";
					when "10110010000110010" => rgb <= "000000";
					when "10110010000110011" => rgb <= "000000";
					when "10110010000110100" => rgb <= "000000";
					when "10110010000110101" => rgb <= "000000";
					when "10110010000110110" => rgb <= "000000";
					when "10110010000110111" => rgb <= "000000";
					when "10110010000111000" => rgb <= "000000";
					when "10110010000111001" => rgb <= "010101";
					when "10110010000111010" => rgb <= "111111";
					when "10110010000111011" => rgb <= "101010";
					when "10110010000111100" => rgb <= "101010";
					when "10110010000111101" => rgb <= "111111";
					when "10110010000111110" => rgb <= "101010";
					when "10110010000111111" => rgb <= "111111";
					when "10110010001000000" => rgb <= "111111";
					when "10110010001000001" => rgb <= "000000";
					when "10110010001000010" => rgb <= "000000";
					when "10110010001000011" => rgb <= "000000";
					when "10110010001000100" => rgb <= "000000";
					when "10110010001000101" => rgb <= "000000";
					when "10110010001000110" => rgb <= "000000";
					when "10110010001000111" => rgb <= "000000";
					when "10110010001001000" => rgb <= "000000";
					when "10110010001001001" => rgb <= "000000";
					when "10110010001001010" => rgb <= "000000";
					when "10110010001001011" => rgb <= "000000";
					when "10110010001001100" => rgb <= "000000";
					when "10110010001001101" => rgb <= "000000";
					when "10110010001001110" => rgb <= "000000";
					when "10110010001001111" => rgb <= "000000";
					when "10110010001010000" => rgb <= "101010";
					when "10110010001010001" => rgb <= "101010";
					when "10110010001010010" => rgb <= "101010";
					when "10110010001010011" => rgb <= "101010";
					when "10110010001010100" => rgb <= "111111";
					when "10110010001010101" => rgb <= "111111";
					when "10110010001010110" => rgb <= "111111";
					when "10110010001010111" => rgb <= "111111";
					when "10110010001011000" => rgb <= "111111";
					when "10110010001011001" => rgb <= "111111";
					when "10110010001011010" => rgb <= "111111";
					when "10110010001011011" => rgb <= "101010";
					when "10110010001011100" => rgb <= "111111";
					when "10110010001011101" => rgb <= "101010";
					when "10110010001011110" => rgb <= "101010";
					when "10110010001011111" => rgb <= "000000";
					when "10110010001100000" => rgb <= "000000";
					when "10110010001100001" => rgb <= "000000";
					when "10110010001100010" => rgb <= "000000";
					when "10110010001100011" => rgb <= "000000";
					when "10110010001100100" => rgb <= "000000";
					when "10110010001100101" => rgb <= "000000";
					when "10110010001100110" => rgb <= "010101";
					when "10110010001100111" => rgb <= "111111";
					when "10110010001101000" => rgb <= "101010";
					when "10110010001101001" => rgb <= "111111";
					when "10110010001101010" => rgb <= "101010";
					when "10110010001101011" => rgb <= "111111";
					when "10110010001101100" => rgb <= "101010";
					when "10110010001101101" => rgb <= "101010";
					when "10110010001101110" => rgb <= "000000";
					when "10110010001101111" => rgb <= "000000";
					when "10110010001110000" => rgb <= "000000";
					when "10110010001110001" => rgb <= "000000";
					when "10110010001110010" => rgb <= "000000";
					when "10110010001110011" => rgb <= "000000";
					when "10110010001110100" => rgb <= "000000";
					when "10110010001110101" => rgb <= "000000";
					when "10110010001110110" => rgb <= "000000";
					when "10110010001110111" => rgb <= "000000";
					when "10110010001111000" => rgb <= "000000";
					when "10110010001111001" => rgb <= "000000";
					when "10110010001111010" => rgb <= "000000";
					when "10110010001111011" => rgb <= "000000";
					when "10110010001111100" => rgb <= "000000";
					when "10110010001111101" => rgb <= "101010";
					when "10110010001111110" => rgb <= "111111";
					when "10110010001111111" => rgb <= "111111";
					when "10110010010000000" => rgb <= "111111";
					when "10110010010000001" => rgb <= "111111";
					when "10110010010000010" => rgb <= "111111";
					when "10110010010000011" => rgb <= "111111";
					when "10110010010000100" => rgb <= "111111";
					when "10110010010000101" => rgb <= "111111";
					when "10110010010000110" => rgb <= "111111";
					when "10110010010000111" => rgb <= "111111";
					when "10110010010001000" => rgb <= "111111";
					when "10110010010001001" => rgb <= "111111";
					when "10110010010001010" => rgb <= "111111";
					when "10110010010001011" => rgb <= "101010";
					when "10110010010001100" => rgb <= "000000";
					when "10110010010001101" => rgb <= "000000";
					when "10110010010001110" => rgb <= "000000";
					when "10110010010001111" => rgb <= "000000";
					when "10110010010010000" => rgb <= "000000";
					when "10110010010010001" => rgb <= "000000";
					when "10110010010010010" => rgb <= "000000";
					when "10110010010010011" => rgb <= "000000";
					when "10110010010010100" => rgb <= "000000";
					when "10110010010010101" => rgb <= "000000";
					when "10110010010010110" => rgb <= "000000";
					when "10110010010010111" => rgb <= "000000";
					when "10110010010011000" => rgb <= "000000";
					when "10110010010011001" => rgb <= "000000";
					when "10110010010011010" => rgb <= "000000";
					when "10110010010011011" => rgb <= "000000";
					when "10110010010011100" => rgb <= "000000";
					when "10110010010011101" => rgb <= "000000";
					when "10110010010011110" => rgb <= "000000";
					when "10110010010011111" => rgb <= "000000";
					when "10110010010100000" => rgb <= "000000";
					when "10110010010100001" => rgb <= "000000";
					when "10110010010100010" => rgb <= "010101";
					when "10110010010100011" => rgb <= "111111";
					when "10110010010100100" => rgb <= "101010";
					when "10110010010100101" => rgb <= "111111";
					when "10110010010100110" => rgb <= "111111";
					when "10110010010100111" => rgb <= "111111";
					when "10110010010101000" => rgb <= "111111";
					when "10110010010101001" => rgb <= "111111";
					when "10110010010101010" => rgb <= "000000";
					when "10110010010101011" => rgb <= "000000";
					when "10110010010101100" => rgb <= "000000";
					when "10110010010101101" => rgb <= "000000";
					when "10110010010101110" => rgb <= "000000";
					when "10110010010101111" => rgb <= "000000";
					when "10110010010110000" => rgb <= "000000";
					when "10110010010110001" => rgb <= "000000";
					when "10110010010110010" => rgb <= "000000";
					when "10110010010110011" => rgb <= "000000";
					when "10110010010110100" => rgb <= "000000";
					when "10110010010110101" => rgb <= "000000";
					when "10110010010110110" => rgb <= "000000";
					when "10110010010110111" => rgb <= "000000";
					when "10110010010111000" => rgb <= "000000";
					when "10110010010111001" => rgb <= "000000";
					when "10110010010111010" => rgb <= "000000";
					when "10110010010111011" => rgb <= "000000";
					when "10110010010111100" => rgb <= "000000";
					when "10110010010111101" => rgb <= "000000";
					when "10110010010111110" => rgb <= "000000";
					when "10110010010111111" => rgb <= "000000";
					when "10110010011000000" => rgb <= "010101";
					when "10110010011000001" => rgb <= "101010";
					when "10110010011000010" => rgb <= "101010";
					when "10110010011000011" => rgb <= "111111";
					when "10110010011000100" => rgb <= "111111";
					when "10110010011000101" => rgb <= "111111";
					when "10110010011000110" => rgb <= "111111";
					when "10110010011000111" => rgb <= "111111";
					when "10110010011001000" => rgb <= "111111";
					when "10110010011001001" => rgb <= "111111";
					when "10110010011001010" => rgb <= "111111";
					when "10110010011001011" => rgb <= "101010";
					when "10110010011001100" => rgb <= "111111";
					when "10110010011001101" => rgb <= "101010";
					when "10110010011001110" => rgb <= "111111";
					when "10110010011001111" => rgb <= "101010";
					when "10110010011010000" => rgb <= "000000";
					when "10110010011010001" => rgb <= "000000";
					when "10110010011010010" => rgb <= "000000";
					when "10110010011010011" => rgb <= "000000";
					when "10110010011010100" => rgb <= "000000";
					when "10110010011010101" => rgb <= "000000";
					when "10110010011010110" => rgb <= "000000";
					when "10110010011010111" => rgb <= "101010";
					when "10110010011011000" => rgb <= "101010";
					when "10110010011011001" => rgb <= "101010";
					when "10110010011011010" => rgb <= "101010";
					when "10110010011011011" => rgb <= "111111";
					when "10110010011011100" => rgb <= "111111";
					when "10110010011011101" => rgb <= "111111";
					when "10110010011011110" => rgb <= "111111";
					when "10110010011011111" => rgb <= "111111";
					when "10110010011100000" => rgb <= "111111";
					when "10110010011100001" => rgb <= "111111";
					when "10110010011100010" => rgb <= "111111";
					when "10110010011100011" => rgb <= "101010";
					when "10110010011100100" => rgb <= "111111";
					when "10110010011100101" => rgb <= "111111";
					when "10110010011100110" => rgb <= "000000";
					when "10110010011100111" => rgb <= "000000";
					when "10110010011101000" => rgb <= "000000";
					when "10110010011101001" => rgb <= "000000";
					when "10110010011101010" => rgb <= "000000";
					when "10110010011101011" => rgb <= "000000";
					when "10110010011101100" => rgb <= "000000";
					when "10110010011101101" => rgb <= "010101";
					when "10110010011101110" => rgb <= "111111";
					when "10110010011101111" => rgb <= "101010";
					when "10110010011110000" => rgb <= "111111";
					when "10110010011110001" => rgb <= "111111";
					when "10110010011110010" => rgb <= "101010";
					when "10110010011110011" => rgb <= "101010";
					when "10110010011110100" => rgb <= "101010";
					when "10110010011110101" => rgb <= "000000";
					when "10110010011110110" => rgb <= "000000";
					when "10110010011110111" => rgb <= "000000";
					when "10110010011111000" => rgb <= "000000";
					when "10110010011111001" => rgb <= "000000";
					when "10110010011111010" => rgb <= "000000";
					when "10110010011111011" => rgb <= "000000";
					when "10110010011111100" => rgb <= "010101";
					when "10110010011111101" => rgb <= "111111";
					when "10110010011111110" => rgb <= "111111";
					when "10110010011111111" => rgb <= "101010";
					when "10110010100000000" => rgb <= "101010";
					when "10110010100000001" => rgb <= "111111";
					when "10110010100000010" => rgb <= "111111";
					when "10110010100000011" => rgb <= "101010";
					when "10110010100000100" => rgb <= "000000";
					when "10110010100000101" => rgb <= "000000";
					when "10110010100000110" => rgb <= "000000";
					when "10110010100000111" => rgb <= "000000";
					when "10110010100001000" => rgb <= "000000";
					when "10110010100001001" => rgb <= "000000";
					when "10110010100001010" => rgb <= "000000";
					when "10110010100001011" => rgb <= "010101";
					when "10110010100001100" => rgb <= "111111";
					when "10110010100001101" => rgb <= "101010";
					when "10110010100001110" => rgb <= "101010";
					when "10110010100001111" => rgb <= "111111";
					when "10110010100010000" => rgb <= "111111";
					when "10110010100010001" => rgb <= "111111";
					when "10110010100010010" => rgb <= "111111";
					when "10110010100010011" => rgb <= "111111";
					when "10110010100010100" => rgb <= "111111";
					when "10110010100010101" => rgb <= "111111";
					when "10110010100010110" => rgb <= "111111";
					when "10110010100010111" => rgb <= "111111";
					when "10110010100011000" => rgb <= "101010";
					when "10110010100011001" => rgb <= "111111";
					when "10110010100011010" => rgb <= "101010";
					when "10110010100011011" => rgb <= "000000";
					when "10110010100011100" => rgb <= "000000";
					when "10110010100011101" => rgb <= "000000";
					when "10110010100011110" => rgb <= "000000";
					when "10110010100011111" => rgb <= "000000";
					when "10110010100100000" => rgb <= "000000";
					when "10110010100100001" => rgb <= "000000";
					when "10110010100100010" => rgb <= "101010";
					when "10110010100100011" => rgb <= "101010";
					when "10110010100100100" => rgb <= "101010";
					when "10110010100100101" => rgb <= "111111";
					when "10110010100100110" => rgb <= "111111";
					when "10110010100100111" => rgb <= "111111";
					when "10110010100101000" => rgb <= "111111";
					when "10110010100101001" => rgb <= "111111";
					when "10110010100101010" => rgb <= "111111";
					when "10110010100101011" => rgb <= "111111";
					when "10110010100101100" => rgb <= "111111";
					when "10110010100101101" => rgb <= "111111";
					when "10110010100101110" => rgb <= "101010";
					when "10110010100101111" => rgb <= "101010";
					when "10110010100110000" => rgb <= "111111";
					when "10110010100110001" => rgb <= "010101";
					when "10110010100110010" => rgb <= "000000";
					when "10110010100110011" => rgb <= "000000";
					when "10110010100110100" => rgb <= "000000";
					when "10110010100110101" => rgb <= "000000";
					when "10110010100110110" => rgb <= "000000";
					when "10110010100110111" => rgb <= "000000";
					when "10110010100111000" => rgb <= "000000";
					when "10110010100111001" => rgb <= "000000";
					when "10110010100111010" => rgb <= "000000";
					when "10110010100111011" => rgb <= "000000";
					when "10110010100111100" => rgb <= "000000";
					when "10110010100111101" => rgb <= "000000";
					when "10110010100111110" => rgb <= "000000";
					when "10110010100111111" => rgb <= "000000";
					when "10110011000000000" => rgb <= "000000";
					when "10110011000000001" => rgb <= "000000";
					when "10110011000000010" => rgb <= "000000";
					when "10110011000000011" => rgb <= "000000";
					when "10110011000000100" => rgb <= "000000";
					when "10110011000000101" => rgb <= "101010";
					when "10110011000000110" => rgb <= "101010";
					when "10110011000000111" => rgb <= "111111";
					when "10110011000001000" => rgb <= "111111";
					when "10110011000001001" => rgb <= "101010";
					when "10110011000001010" => rgb <= "101010";
					when "10110011000001011" => rgb <= "111111";
					when "10110011000001100" => rgb <= "010101";
					when "10110011000001101" => rgb <= "000000";
					when "10110011000001110" => rgb <= "000000";
					when "10110011000001111" => rgb <= "000000";
					when "10110011000010000" => rgb <= "000000";
					when "10110011000010001" => rgb <= "000000";
					when "10110011000010010" => rgb <= "000000";
					when "10110011000010011" => rgb <= "000000";
					when "10110011000010100" => rgb <= "000000";
					when "10110011000010101" => rgb <= "000000";
					when "10110011000010110" => rgb <= "000000";
					when "10110011000010111" => rgb <= "000000";
					when "10110011000011000" => rgb <= "000000";
					when "10110011000011001" => rgb <= "000000";
					when "10110011000011010" => rgb <= "000000";
					when "10110011000011011" => rgb <= "010101";
					when "10110011000011100" => rgb <= "111111";
					when "10110011000011101" => rgb <= "111111";
					when "10110011000011110" => rgb <= "101010";
					when "10110011000011111" => rgb <= "111111";
					when "10110011000100000" => rgb <= "101010";
					when "10110011000100001" => rgb <= "101010";
					when "10110011000100010" => rgb <= "101010";
					when "10110011000100011" => rgb <= "101010";
					when "10110011000100100" => rgb <= "111111";
					when "10110011000100101" => rgb <= "111111";
					when "10110011000100110" => rgb <= "101010";
					when "10110011000100111" => rgb <= "101010";
					when "10110011000101000" => rgb <= "111111";
					when "10110011000101001" => rgb <= "101010";
					when "10110011000101010" => rgb <= "101010";
					when "10110011000101011" => rgb <= "111111";
					when "10110011000101100" => rgb <= "111111";
					when "10110011000101101" => rgb <= "101010";
					when "10110011000101110" => rgb <= "101010";
					when "10110011000101111" => rgb <= "101010";
					when "10110011000110000" => rgb <= "111111";
					when "10110011000110001" => rgb <= "101010";
					when "10110011000110010" => rgb <= "000000";
					when "10110011000110011" => rgb <= "000000";
					when "10110011000110100" => rgb <= "000000";
					when "10110011000110101" => rgb <= "000000";
					when "10110011000110110" => rgb <= "000000";
					when "10110011000110111" => rgb <= "000000";
					when "10110011000111000" => rgb <= "000000";
					when "10110011000111001" => rgb <= "010101";
					when "10110011000111010" => rgb <= "111111";
					when "10110011000111011" => rgb <= "101010";
					when "10110011000111100" => rgb <= "111111";
					when "10110011000111101" => rgb <= "111111";
					when "10110011000111110" => rgb <= "101010";
					when "10110011000111111" => rgb <= "111111";
					when "10110011001000000" => rgb <= "101010";
					when "10110011001000001" => rgb <= "000000";
					when "10110011001000010" => rgb <= "000000";
					when "10110011001000011" => rgb <= "000000";
					when "10110011001000100" => rgb <= "000000";
					when "10110011001000101" => rgb <= "000000";
					when "10110011001000110" => rgb <= "000000";
					when "10110011001000111" => rgb <= "000000";
					when "10110011001001000" => rgb <= "000000";
					when "10110011001001001" => rgb <= "000000";
					when "10110011001001010" => rgb <= "000000";
					when "10110011001001011" => rgb <= "000000";
					when "10110011001001100" => rgb <= "000000";
					when "10110011001001101" => rgb <= "000000";
					when "10110011001001110" => rgb <= "000000";
					when "10110011001001111" => rgb <= "000000";
					when "10110011001010000" => rgb <= "101010";
					when "10110011001010001" => rgb <= "101010";
					when "10110011001010010" => rgb <= "101010";
					when "10110011001010011" => rgb <= "101010";
					when "10110011001010100" => rgb <= "111111";
					when "10110011001010101" => rgb <= "111111";
					when "10110011001010110" => rgb <= "111111";
					when "10110011001010111" => rgb <= "111111";
					when "10110011001011000" => rgb <= "111111";
					when "10110011001011001" => rgb <= "111111";
					when "10110011001011010" => rgb <= "111111";
					when "10110011001011011" => rgb <= "101010";
					when "10110011001011100" => rgb <= "111111";
					when "10110011001011101" => rgb <= "101010";
					when "10110011001011110" => rgb <= "101010";
					when "10110011001011111" => rgb <= "000000";
					when "10110011001100000" => rgb <= "000000";
					when "10110011001100001" => rgb <= "000000";
					when "10110011001100010" => rgb <= "000000";
					when "10110011001100011" => rgb <= "000000";
					when "10110011001100100" => rgb <= "000000";
					when "10110011001100101" => rgb <= "000000";
					when "10110011001100110" => rgb <= "010101";
					when "10110011001100111" => rgb <= "111111";
					when "10110011001101000" => rgb <= "101010";
					when "10110011001101001" => rgb <= "111111";
					when "10110011001101010" => rgb <= "101010";
					when "10110011001101011" => rgb <= "111111";
					when "10110011001101100" => rgb <= "101010";
					when "10110011001101101" => rgb <= "101010";
					when "10110011001101110" => rgb <= "000000";
					when "10110011001101111" => rgb <= "000000";
					when "10110011001110000" => rgb <= "000000";
					when "10110011001110001" => rgb <= "000000";
					when "10110011001110010" => rgb <= "000000";
					when "10110011001110011" => rgb <= "000000";
					when "10110011001110100" => rgb <= "000000";
					when "10110011001110101" => rgb <= "000000";
					when "10110011001110110" => rgb <= "000000";
					when "10110011001110111" => rgb <= "000000";
					when "10110011001111000" => rgb <= "000000";
					when "10110011001111001" => rgb <= "000000";
					when "10110011001111010" => rgb <= "000000";
					when "10110011001111011" => rgb <= "000000";
					when "10110011001111100" => rgb <= "000000";
					when "10110011001111101" => rgb <= "101010";
					when "10110011001111110" => rgb <= "111111";
					when "10110011001111111" => rgb <= "111111";
					when "10110011010000000" => rgb <= "111111";
					when "10110011010000001" => rgb <= "111111";
					when "10110011010000010" => rgb <= "111111";
					when "10110011010000011" => rgb <= "111111";
					when "10110011010000100" => rgb <= "111111";
					when "10110011010000101" => rgb <= "111111";
					when "10110011010000110" => rgb <= "111111";
					when "10110011010000111" => rgb <= "111111";
					when "10110011010001000" => rgb <= "111111";
					when "10110011010001001" => rgb <= "111111";
					when "10110011010001010" => rgb <= "111111";
					when "10110011010001011" => rgb <= "101010";
					when "10110011010001100" => rgb <= "000000";
					when "10110011010001101" => rgb <= "000000";
					when "10110011010001110" => rgb <= "000000";
					when "10110011010001111" => rgb <= "000000";
					when "10110011010010000" => rgb <= "000000";
					when "10110011010010001" => rgb <= "000000";
					when "10110011010010010" => rgb <= "000000";
					when "10110011010010011" => rgb <= "000000";
					when "10110011010010100" => rgb <= "000000";
					when "10110011010010101" => rgb <= "000000";
					when "10110011010010110" => rgb <= "000000";
					when "10110011010010111" => rgb <= "000000";
					when "10110011010011000" => rgb <= "000000";
					when "10110011010011001" => rgb <= "000000";
					when "10110011010011010" => rgb <= "000000";
					when "10110011010011011" => rgb <= "000000";
					when "10110011010011100" => rgb <= "000000";
					when "10110011010011101" => rgb <= "000000";
					when "10110011010011110" => rgb <= "000000";
					when "10110011010011111" => rgb <= "000000";
					when "10110011010100000" => rgb <= "000000";
					when "10110011010100001" => rgb <= "000000";
					when "10110011010100010" => rgb <= "010101";
					when "10110011010100011" => rgb <= "111111";
					when "10110011010100100" => rgb <= "101010";
					when "10110011010100101" => rgb <= "111111";
					when "10110011010100110" => rgb <= "111111";
					when "10110011010100111" => rgb <= "111111";
					when "10110011010101000" => rgb <= "111111";
					when "10110011010101001" => rgb <= "111111";
					when "10110011010101010" => rgb <= "000000";
					when "10110011010101011" => rgb <= "000000";
					when "10110011010101100" => rgb <= "000000";
					when "10110011010101101" => rgb <= "000000";
					when "10110011010101110" => rgb <= "000000";
					when "10110011010101111" => rgb <= "000000";
					when "10110011010110000" => rgb <= "000000";
					when "10110011010110001" => rgb <= "000000";
					when "10110011010110010" => rgb <= "000000";
					when "10110011010110011" => rgb <= "000000";
					when "10110011010110100" => rgb <= "000000";
					when "10110011010110101" => rgb <= "000000";
					when "10110011010110110" => rgb <= "000000";
					when "10110011010110111" => rgb <= "000000";
					when "10110011010111000" => rgb <= "000000";
					when "10110011010111001" => rgb <= "000000";
					when "10110011010111010" => rgb <= "000000";
					when "10110011010111011" => rgb <= "000000";
					when "10110011010111100" => rgb <= "000000";
					when "10110011010111101" => rgb <= "000000";
					when "10110011010111110" => rgb <= "000000";
					when "10110011010111111" => rgb <= "000000";
					when "10110011011000000" => rgb <= "010101";
					when "10110011011000001" => rgb <= "101010";
					when "10110011011000010" => rgb <= "101010";
					when "10110011011000011" => rgb <= "111111";
					when "10110011011000100" => rgb <= "111111";
					when "10110011011000101" => rgb <= "111111";
					when "10110011011000110" => rgb <= "111111";
					when "10110011011000111" => rgb <= "111111";
					when "10110011011001000" => rgb <= "111111";
					when "10110011011001001" => rgb <= "111111";
					when "10110011011001010" => rgb <= "111111";
					when "10110011011001011" => rgb <= "101010";
					when "10110011011001100" => rgb <= "111111";
					when "10110011011001101" => rgb <= "101010";
					when "10110011011001110" => rgb <= "111111";
					when "10110011011001111" => rgb <= "101010";
					when "10110011011010000" => rgb <= "000000";
					when "10110011011010001" => rgb <= "000000";
					when "10110011011010010" => rgb <= "000000";
					when "10110011011010011" => rgb <= "000000";
					when "10110011011010100" => rgb <= "000000";
					when "10110011011010101" => rgb <= "000000";
					when "10110011011010110" => rgb <= "000000";
					when "10110011011010111" => rgb <= "101010";
					when "10110011011011000" => rgb <= "101010";
					when "10110011011011001" => rgb <= "101010";
					when "10110011011011010" => rgb <= "101010";
					when "10110011011011011" => rgb <= "111111";
					when "10110011011011100" => rgb <= "111111";
					when "10110011011011101" => rgb <= "111111";
					when "10110011011011110" => rgb <= "111111";
					when "10110011011011111" => rgb <= "111111";
					when "10110011011100000" => rgb <= "111111";
					when "10110011011100001" => rgb <= "111111";
					when "10110011011100010" => rgb <= "111111";
					when "10110011011100011" => rgb <= "101010";
					when "10110011011100100" => rgb <= "111111";
					when "10110011011100101" => rgb <= "111111";
					when "10110011011100110" => rgb <= "000000";
					when "10110011011100111" => rgb <= "000000";
					when "10110011011101000" => rgb <= "000000";
					when "10110011011101001" => rgb <= "000000";
					when "10110011011101010" => rgb <= "000000";
					when "10110011011101011" => rgb <= "000000";
					when "10110011011101100" => rgb <= "000000";
					when "10110011011101101" => rgb <= "010101";
					when "10110011011101110" => rgb <= "111111";
					when "10110011011101111" => rgb <= "101010";
					when "10110011011110000" => rgb <= "111111";
					when "10110011011110001" => rgb <= "111111";
					when "10110011011110010" => rgb <= "101010";
					when "10110011011110011" => rgb <= "111111";
					when "10110011011110100" => rgb <= "101010";
					when "10110011011110101" => rgb <= "000000";
					when "10110011011110110" => rgb <= "000000";
					when "10110011011110111" => rgb <= "000000";
					when "10110011011111000" => rgb <= "000000";
					when "10110011011111001" => rgb <= "000000";
					when "10110011011111010" => rgb <= "000000";
					when "10110011011111011" => rgb <= "000000";
					when "10110011011111100" => rgb <= "010101";
					when "10110011011111101" => rgb <= "111111";
					when "10110011011111110" => rgb <= "101010";
					when "10110011011111111" => rgb <= "111111";
					when "10110011100000000" => rgb <= "111111";
					when "10110011100000001" => rgb <= "101010";
					when "10110011100000010" => rgb <= "101010";
					when "10110011100000011" => rgb <= "111111";
					when "10110011100000100" => rgb <= "000000";
					when "10110011100000101" => rgb <= "000000";
					when "10110011100000110" => rgb <= "000000";
					when "10110011100000111" => rgb <= "000000";
					when "10110011100001000" => rgb <= "000000";
					when "10110011100001001" => rgb <= "000000";
					when "10110011100001010" => rgb <= "000000";
					when "10110011100001011" => rgb <= "010101";
					when "10110011100001100" => rgb <= "111111";
					when "10110011100001101" => rgb <= "111111";
					when "10110011100001110" => rgb <= "101010";
					when "10110011100001111" => rgb <= "101010";
					when "10110011100010000" => rgb <= "111111";
					when "10110011100010001" => rgb <= "111111";
					when "10110011100010010" => rgb <= "111111";
					when "10110011100010011" => rgb <= "111111";
					when "10110011100010100" => rgb <= "111111";
					when "10110011100010101" => rgb <= "111111";
					when "10110011100010110" => rgb <= "111111";
					when "10110011100010111" => rgb <= "111111";
					when "10110011100011000" => rgb <= "101010";
					when "10110011100011001" => rgb <= "111111";
					when "10110011100011010" => rgb <= "101010";
					when "10110011100011011" => rgb <= "000000";
					when "10110011100011100" => rgb <= "000000";
					when "10110011100011101" => rgb <= "000000";
					when "10110011100011110" => rgb <= "000000";
					when "10110011100011111" => rgb <= "000000";
					when "10110011100100000" => rgb <= "000000";
					when "10110011100100001" => rgb <= "000000";
					when "10110011100100010" => rgb <= "101010";
					when "10110011100100011" => rgb <= "101010";
					when "10110011100100100" => rgb <= "101010";
					when "10110011100100101" => rgb <= "111111";
					when "10110011100100110" => rgb <= "111111";
					when "10110011100100111" => rgb <= "111111";
					when "10110011100101000" => rgb <= "111111";
					when "10110011100101001" => rgb <= "111111";
					when "10110011100101010" => rgb <= "111111";
					when "10110011100101011" => rgb <= "111111";
					when "10110011100101100" => rgb <= "111111";
					when "10110011100101101" => rgb <= "111111";
					when "10110011100101110" => rgb <= "101010";
					when "10110011100101111" => rgb <= "101010";
					when "10110011100110000" => rgb <= "111111";
					when "10110011100110001" => rgb <= "010101";
					when "10110011100110010" => rgb <= "000000";
					when "10110011100110011" => rgb <= "000000";
					when "10110011100110100" => rgb <= "000000";
					when "10110011100110101" => rgb <= "000000";
					when "10110011100110110" => rgb <= "000000";
					when "10110011100110111" => rgb <= "000000";
					when "10110011100111000" => rgb <= "000000";
					when "10110011100111001" => rgb <= "000000";
					when "10110011100111010" => rgb <= "000000";
					when "10110011100111011" => rgb <= "000000";
					when "10110011100111100" => rgb <= "000000";
					when "10110011100111101" => rgb <= "000000";
					when "10110011100111110" => rgb <= "000000";
					when "10110011100111111" => rgb <= "000000";
					when "10110100000000000" => rgb <= "000000";
					when "10110100000000001" => rgb <= "000000";
					when "10110100000000010" => rgb <= "000000";
					when "10110100000000011" => rgb <= "000000";
					when "10110100000000100" => rgb <= "000000";
					when "10110100000000101" => rgb <= "101010";
					when "10110100000000110" => rgb <= "111111";
					when "10110100000000111" => rgb <= "111111";
					when "10110100000001000" => rgb <= "111111";
					when "10110100000001001" => rgb <= "101010";
					when "10110100000001010" => rgb <= "111111";
					when "10110100000001011" => rgb <= "101010";
					when "10110100000001100" => rgb <= "101010";
					when "10110100000001101" => rgb <= "000000";
					when "10110100000001110" => rgb <= "000000";
					when "10110100000001111" => rgb <= "000000";
					when "10110100000010000" => rgb <= "000000";
					when "10110100000010001" => rgb <= "000000";
					when "10110100000010010" => rgb <= "000000";
					when "10110100000010011" => rgb <= "000000";
					when "10110100000010100" => rgb <= "000000";
					when "10110100000010101" => rgb <= "000000";
					when "10110100000010110" => rgb <= "000000";
					when "10110100000010111" => rgb <= "000000";
					when "10110100000011000" => rgb <= "000000";
					when "10110100000011001" => rgb <= "000000";
					when "10110100000011010" => rgb <= "000000";
					when "10110100000011011" => rgb <= "010101";
					when "10110100000011100" => rgb <= "111111";
					when "10110100000011101" => rgb <= "101010";
					when "10110100000011110" => rgb <= "101010";
					when "10110100000011111" => rgb <= "111111";
					when "10110100000100000" => rgb <= "111111";
					when "10110100000100001" => rgb <= "111111";
					when "10110100000100010" => rgb <= "111111";
					when "10110100000100011" => rgb <= "111111";
					when "10110100000100100" => rgb <= "111111";
					when "10110100000100101" => rgb <= "111111";
					when "10110100000100110" => rgb <= "111111";
					when "10110100000100111" => rgb <= "111111";
					when "10110100000101000" => rgb <= "111111";
					when "10110100000101001" => rgb <= "111111";
					when "10110100000101010" => rgb <= "111111";
					when "10110100000101011" => rgb <= "101010";
					when "10110100000101100" => rgb <= "101010";
					when "10110100000101101" => rgb <= "111111";
					when "10110100000101110" => rgb <= "111111";
					when "10110100000101111" => rgb <= "101010";
					when "10110100000110000" => rgb <= "101010";
					when "10110100000110001" => rgb <= "111111";
					when "10110100000110010" => rgb <= "000000";
					when "10110100000110011" => rgb <= "000000";
					when "10110100000110100" => rgb <= "000000";
					when "10110100000110101" => rgb <= "000000";
					when "10110100000110110" => rgb <= "000000";
					when "10110100000110111" => rgb <= "000000";
					when "10110100000111000" => rgb <= "000000";
					when "10110100000111001" => rgb <= "010101";
					when "10110100000111010" => rgb <= "111111";
					when "10110100000111011" => rgb <= "101010";
					when "10110100000111100" => rgb <= "111111";
					when "10110100000111101" => rgb <= "111111";
					when "10110100000111110" => rgb <= "101010";
					when "10110100000111111" => rgb <= "111111";
					when "10110100001000000" => rgb <= "101010";
					when "10110100001000001" => rgb <= "000000";
					when "10110100001000010" => rgb <= "000000";
					when "10110100001000011" => rgb <= "000000";
					when "10110100001000100" => rgb <= "000000";
					when "10110100001000101" => rgb <= "000000";
					when "10110100001000110" => rgb <= "000000";
					when "10110100001000111" => rgb <= "000000";
					when "10110100001001000" => rgb <= "000000";
					when "10110100001001001" => rgb <= "000000";
					when "10110100001001010" => rgb <= "000000";
					when "10110100001001011" => rgb <= "000000";
					when "10110100001001100" => rgb <= "000000";
					when "10110100001001101" => rgb <= "000000";
					when "10110100001001110" => rgb <= "000000";
					when "10110100001001111" => rgb <= "000000";
					when "10110100001010000" => rgb <= "101010";
					when "10110100001010001" => rgb <= "101010";
					when "10110100001010010" => rgb <= "101010";
					when "10110100001010011" => rgb <= "101010";
					when "10110100001010100" => rgb <= "111111";
					when "10110100001010101" => rgb <= "111111";
					when "10110100001010110" => rgb <= "111111";
					when "10110100001010111" => rgb <= "111111";
					when "10110100001011000" => rgb <= "111111";
					when "10110100001011001" => rgb <= "111111";
					when "10110100001011010" => rgb <= "111111";
					when "10110100001011011" => rgb <= "101010";
					when "10110100001011100" => rgb <= "111111";
					when "10110100001011101" => rgb <= "101010";
					when "10110100001011110" => rgb <= "101010";
					when "10110100001011111" => rgb <= "000000";
					when "10110100001100000" => rgb <= "000000";
					when "10110100001100001" => rgb <= "000000";
					when "10110100001100010" => rgb <= "000000";
					when "10110100001100011" => rgb <= "000000";
					when "10110100001100100" => rgb <= "000000";
					when "10110100001100101" => rgb <= "000000";
					when "10110100001100110" => rgb <= "010101";
					when "10110100001100111" => rgb <= "111111";
					when "10110100001101000" => rgb <= "101010";
					when "10110100001101001" => rgb <= "111111";
					when "10110100001101010" => rgb <= "101010";
					when "10110100001101011" => rgb <= "111111";
					when "10110100001101100" => rgb <= "101010";
					when "10110100001101101" => rgb <= "101010";
					when "10110100001101110" => rgb <= "000000";
					when "10110100001101111" => rgb <= "000000";
					when "10110100001110000" => rgb <= "000000";
					when "10110100001110001" => rgb <= "000000";
					when "10110100001110010" => rgb <= "000000";
					when "10110100001110011" => rgb <= "000000";
					when "10110100001110100" => rgb <= "000000";
					when "10110100001110101" => rgb <= "000000";
					when "10110100001110110" => rgb <= "000000";
					when "10110100001110111" => rgb <= "000000";
					when "10110100001111000" => rgb <= "000000";
					when "10110100001111001" => rgb <= "000000";
					when "10110100001111010" => rgb <= "000000";
					when "10110100001111011" => rgb <= "000000";
					when "10110100001111100" => rgb <= "000000";
					when "10110100001111101" => rgb <= "101010";
					when "10110100001111110" => rgb <= "111111";
					when "10110100001111111" => rgb <= "111111";
					when "10110100010000000" => rgb <= "111111";
					when "10110100010000001" => rgb <= "111111";
					when "10110100010000010" => rgb <= "111111";
					when "10110100010000011" => rgb <= "111111";
					when "10110100010000100" => rgb <= "111111";
					when "10110100010000101" => rgb <= "111111";
					when "10110100010000110" => rgb <= "111111";
					when "10110100010000111" => rgb <= "111111";
					when "10110100010001000" => rgb <= "111111";
					when "10110100010001001" => rgb <= "111111";
					when "10110100010001010" => rgb <= "111111";
					when "10110100010001011" => rgb <= "101010";
					when "10110100010001100" => rgb <= "000000";
					when "10110100010001101" => rgb <= "000000";
					when "10110100010001110" => rgb <= "000000";
					when "10110100010001111" => rgb <= "000000";
					when "10110100010010000" => rgb <= "000000";
					when "10110100010010001" => rgb <= "000000";
					when "10110100010010010" => rgb <= "000000";
					when "10110100010010011" => rgb <= "000000";
					when "10110100010010100" => rgb <= "000000";
					when "10110100010010101" => rgb <= "000000";
					when "10110100010010110" => rgb <= "000000";
					when "10110100010010111" => rgb <= "000000";
					when "10110100010011000" => rgb <= "000000";
					when "10110100010011001" => rgb <= "000000";
					when "10110100010011010" => rgb <= "000000";
					when "10110100010011011" => rgb <= "000000";
					when "10110100010011100" => rgb <= "000000";
					when "10110100010011101" => rgb <= "000000";
					when "10110100010011110" => rgb <= "000000";
					when "10110100010011111" => rgb <= "000000";
					when "10110100010100000" => rgb <= "000000";
					when "10110100010100001" => rgb <= "000000";
					when "10110100010100010" => rgb <= "010101";
					when "10110100010100011" => rgb <= "111111";
					when "10110100010100100" => rgb <= "101010";
					when "10110100010100101" => rgb <= "111111";
					when "10110100010100110" => rgb <= "111111";
					when "10110100010100111" => rgb <= "111111";
					when "10110100010101000" => rgb <= "111111";
					when "10110100010101001" => rgb <= "111111";
					when "10110100010101010" => rgb <= "000000";
					when "10110100010101011" => rgb <= "000000";
					when "10110100010101100" => rgb <= "000000";
					when "10110100010101101" => rgb <= "000000";
					when "10110100010101110" => rgb <= "000000";
					when "10110100010101111" => rgb <= "000000";
					when "10110100010110000" => rgb <= "000000";
					when "10110100010110001" => rgb <= "000000";
					when "10110100010110010" => rgb <= "000000";
					when "10110100010110011" => rgb <= "000000";
					when "10110100010110100" => rgb <= "000000";
					when "10110100010110101" => rgb <= "000000";
					when "10110100010110110" => rgb <= "000000";
					when "10110100010110111" => rgb <= "000000";
					when "10110100010111000" => rgb <= "000000";
					when "10110100010111001" => rgb <= "000000";
					when "10110100010111010" => rgb <= "000000";
					when "10110100010111011" => rgb <= "000000";
					when "10110100010111100" => rgb <= "000000";
					when "10110100010111101" => rgb <= "000000";
					when "10110100010111110" => rgb <= "000000";
					when "10110100010111111" => rgb <= "000000";
					when "10110100011000000" => rgb <= "010101";
					when "10110100011000001" => rgb <= "101010";
					when "10110100011000010" => rgb <= "101010";
					when "10110100011000011" => rgb <= "111111";
					when "10110100011000100" => rgb <= "111111";
					when "10110100011000101" => rgb <= "111111";
					when "10110100011000110" => rgb <= "111111";
					when "10110100011000111" => rgb <= "111111";
					when "10110100011001000" => rgb <= "111111";
					when "10110100011001001" => rgb <= "111111";
					when "10110100011001010" => rgb <= "111111";
					when "10110100011001011" => rgb <= "101010";
					when "10110100011001100" => rgb <= "111111";
					when "10110100011001101" => rgb <= "101010";
					when "10110100011001110" => rgb <= "111111";
					when "10110100011001111" => rgb <= "101010";
					when "10110100011010000" => rgb <= "000000";
					when "10110100011010001" => rgb <= "000000";
					when "10110100011010010" => rgb <= "000000";
					when "10110100011010011" => rgb <= "000000";
					when "10110100011010100" => rgb <= "000000";
					when "10110100011010101" => rgb <= "000000";
					when "10110100011010110" => rgb <= "000000";
					when "10110100011010111" => rgb <= "101010";
					when "10110100011011000" => rgb <= "101010";
					when "10110100011011001" => rgb <= "101010";
					when "10110100011011010" => rgb <= "101010";
					when "10110100011011011" => rgb <= "111111";
					when "10110100011011100" => rgb <= "111111";
					when "10110100011011101" => rgb <= "111111";
					when "10110100011011110" => rgb <= "111111";
					when "10110100011011111" => rgb <= "111111";
					when "10110100011100000" => rgb <= "111111";
					when "10110100011100001" => rgb <= "111111";
					when "10110100011100010" => rgb <= "111111";
					when "10110100011100011" => rgb <= "101010";
					when "10110100011100100" => rgb <= "111111";
					when "10110100011100101" => rgb <= "111111";
					when "10110100011100110" => rgb <= "000000";
					when "10110100011100111" => rgb <= "000000";
					when "10110100011101000" => rgb <= "000000";
					when "10110100011101001" => rgb <= "000000";
					when "10110100011101010" => rgb <= "000000";
					when "10110100011101011" => rgb <= "000000";
					when "10110100011101100" => rgb <= "000000";
					when "10110100011101101" => rgb <= "010101";
					when "10110100011101110" => rgb <= "111111";
					when "10110100011101111" => rgb <= "101010";
					when "10110100011110000" => rgb <= "111111";
					when "10110100011110001" => rgb <= "111111";
					when "10110100011110010" => rgb <= "101010";
					when "10110100011110011" => rgb <= "101010";
					when "10110100011110100" => rgb <= "101010";
					when "10110100011110101" => rgb <= "000000";
					when "10110100011110110" => rgb <= "000000";
					when "10110100011110111" => rgb <= "000000";
					when "10110100011111000" => rgb <= "000000";
					when "10110100011111001" => rgb <= "000000";
					when "10110100011111010" => rgb <= "000000";
					when "10110100011111011" => rgb <= "000000";
					when "10110100011111100" => rgb <= "010101";
					when "10110100011111101" => rgb <= "111111";
					when "10110100011111110" => rgb <= "101010";
					when "10110100011111111" => rgb <= "111111";
					when "10110100100000000" => rgb <= "111111";
					when "10110100100000001" => rgb <= "101010";
					when "10110100100000010" => rgb <= "111111";
					when "10110100100000011" => rgb <= "101010";
					when "10110100100000100" => rgb <= "000000";
					when "10110100100000101" => rgb <= "000000";
					when "10110100100000110" => rgb <= "000000";
					when "10110100100000111" => rgb <= "000000";
					when "10110100100001000" => rgb <= "000000";
					when "10110100100001001" => rgb <= "000000";
					when "10110100100001010" => rgb <= "000000";
					when "10110100100001011" => rgb <= "010101";
					when "10110100100001100" => rgb <= "101010";
					when "10110100100001101" => rgb <= "111111";
					when "10110100100001110" => rgb <= "111111";
					when "10110100100001111" => rgb <= "111111";
					when "10110100100010000" => rgb <= "111111";
					when "10110100100010001" => rgb <= "111111";
					when "10110100100010010" => rgb <= "111111";
					when "10110100100010011" => rgb <= "111111";
					when "10110100100010100" => rgb <= "111111";
					when "10110100100010101" => rgb <= "111111";
					when "10110100100010110" => rgb <= "111111";
					when "10110100100010111" => rgb <= "111111";
					when "10110100100011000" => rgb <= "101010";
					when "10110100100011001" => rgb <= "111111";
					when "10110100100011010" => rgb <= "101010";
					when "10110100100011011" => rgb <= "000000";
					when "10110100100011100" => rgb <= "000000";
					when "10110100100011101" => rgb <= "000000";
					when "10110100100011110" => rgb <= "000000";
					when "10110100100011111" => rgb <= "000000";
					when "10110100100100000" => rgb <= "000000";
					when "10110100100100001" => rgb <= "000000";
					when "10110100100100010" => rgb <= "101010";
					when "10110100100100011" => rgb <= "101010";
					when "10110100100100100" => rgb <= "101010";
					when "10110100100100101" => rgb <= "111111";
					when "10110100100100110" => rgb <= "111111";
					when "10110100100100111" => rgb <= "111111";
					when "10110100100101000" => rgb <= "111111";
					when "10110100100101001" => rgb <= "111111";
					when "10110100100101010" => rgb <= "111111";
					when "10110100100101011" => rgb <= "111111";
					when "10110100100101100" => rgb <= "111111";
					when "10110100100101101" => rgb <= "111111";
					when "10110100100101110" => rgb <= "101010";
					when "10110100100101111" => rgb <= "101010";
					when "10110100100110000" => rgb <= "111111";
					when "10110100100110001" => rgb <= "010101";
					when "10110100100110010" => rgb <= "000000";
					when "10110100100110011" => rgb <= "000000";
					when "10110100100110100" => rgb <= "000000";
					when "10110100100110101" => rgb <= "000000";
					when "10110100100110110" => rgb <= "000000";
					when "10110100100110111" => rgb <= "000000";
					when "10110100100111000" => rgb <= "000000";
					when "10110100100111001" => rgb <= "000000";
					when "10110100100111010" => rgb <= "000000";
					when "10110100100111011" => rgb <= "000000";
					when "10110100100111100" => rgb <= "000000";
					when "10110100100111101" => rgb <= "000000";
					when "10110100100111110" => rgb <= "000000";
					when "10110100100111111" => rgb <= "000000";
					when "10110101000000000" => rgb <= "000000";
					when "10110101000000001" => rgb <= "000000";
					when "10110101000000010" => rgb <= "000000";
					when "10110101000000011" => rgb <= "000000";
					when "10110101000000100" => rgb <= "000000";
					when "10110101000000101" => rgb <= "101010";
					when "10110101000000110" => rgb <= "101010";
					when "10110101000000111" => rgb <= "101010";
					when "10110101000001000" => rgb <= "101010";
					when "10110101000001001" => rgb <= "101010";
					when "10110101000001010" => rgb <= "101010";
					when "10110101000001011" => rgb <= "111111";
					when "10110101000001100" => rgb <= "101010";
					when "10110101000001101" => rgb <= "000000";
					when "10110101000001110" => rgb <= "000000";
					when "10110101000001111" => rgb <= "000000";
					when "10110101000010000" => rgb <= "000000";
					when "10110101000010001" => rgb <= "000000";
					when "10110101000010010" => rgb <= "000000";
					when "10110101000010011" => rgb <= "000000";
					when "10110101000010100" => rgb <= "000000";
					when "10110101000010101" => rgb <= "000000";
					when "10110101000010110" => rgb <= "000000";
					when "10110101000010111" => rgb <= "000000";
					when "10110101000011000" => rgb <= "000000";
					when "10110101000011001" => rgb <= "000000";
					when "10110101000011010" => rgb <= "000000";
					when "10110101000011011" => rgb <= "010101";
					when "10110101000011100" => rgb <= "111111";
					when "10110101000011101" => rgb <= "111111";
					when "10110101000011110" => rgb <= "111111";
					when "10110101000011111" => rgb <= "111111";
					when "10110101000100000" => rgb <= "111111";
					when "10110101000100001" => rgb <= "111111";
					when "10110101000100010" => rgb <= "111111";
					when "10110101000100011" => rgb <= "111111";
					when "10110101000100100" => rgb <= "111111";
					when "10110101000100101" => rgb <= "111111";
					when "10110101000100110" => rgb <= "111111";
					when "10110101000100111" => rgb <= "101010";
					when "10110101000101000" => rgb <= "111111";
					when "10110101000101001" => rgb <= "101010";
					when "10110101000101010" => rgb <= "101010";
					when "10110101000101011" => rgb <= "111111";
					when "10110101000101100" => rgb <= "101010";
					when "10110101000101101" => rgb <= "101010";
					when "10110101000101110" => rgb <= "101010";
					when "10110101000101111" => rgb <= "101010";
					when "10110101000110000" => rgb <= "101010";
					when "10110101000110001" => rgb <= "101010";
					when "10110101000110010" => rgb <= "000000";
					when "10110101000110011" => rgb <= "000000";
					when "10110101000110100" => rgb <= "000000";
					when "10110101000110101" => rgb <= "000000";
					when "10110101000110110" => rgb <= "000000";
					when "10110101000110111" => rgb <= "000000";
					when "10110101000111000" => rgb <= "000000";
					when "10110101000111001" => rgb <= "010101";
					when "10110101000111010" => rgb <= "111111";
					when "10110101000111011" => rgb <= "101010";
					when "10110101000111100" => rgb <= "111111";
					when "10110101000111101" => rgb <= "111111";
					when "10110101000111110" => rgb <= "101010";
					when "10110101000111111" => rgb <= "111111";
					when "10110101001000000" => rgb <= "101010";
					when "10110101001000001" => rgb <= "000000";
					when "10110101001000010" => rgb <= "000000";
					when "10110101001000011" => rgb <= "000000";
					when "10110101001000100" => rgb <= "000000";
					when "10110101001000101" => rgb <= "000000";
					when "10110101001000110" => rgb <= "000000";
					when "10110101001000111" => rgb <= "000000";
					when "10110101001001000" => rgb <= "000000";
					when "10110101001001001" => rgb <= "000000";
					when "10110101001001010" => rgb <= "000000";
					when "10110101001001011" => rgb <= "000000";
					when "10110101001001100" => rgb <= "000000";
					when "10110101001001101" => rgb <= "000000";
					when "10110101001001110" => rgb <= "000000";
					when "10110101001001111" => rgb <= "000000";
					when "10110101001010000" => rgb <= "101010";
					when "10110101001010001" => rgb <= "101010";
					when "10110101001010010" => rgb <= "101010";
					when "10110101001010011" => rgb <= "101010";
					when "10110101001010100" => rgb <= "111111";
					when "10110101001010101" => rgb <= "111111";
					when "10110101001010110" => rgb <= "111111";
					when "10110101001010111" => rgb <= "111111";
					when "10110101001011000" => rgb <= "111111";
					when "10110101001011001" => rgb <= "111111";
					when "10110101001011010" => rgb <= "111111";
					when "10110101001011011" => rgb <= "101010";
					when "10110101001011100" => rgb <= "111111";
					when "10110101001011101" => rgb <= "101010";
					when "10110101001011110" => rgb <= "101010";
					when "10110101001011111" => rgb <= "000000";
					when "10110101001100000" => rgb <= "000000";
					when "10110101001100001" => rgb <= "000000";
					when "10110101001100010" => rgb <= "000000";
					when "10110101001100011" => rgb <= "000000";
					when "10110101001100100" => rgb <= "000000";
					when "10110101001100101" => rgb <= "000000";
					when "10110101001100110" => rgb <= "010101";
					when "10110101001100111" => rgb <= "111111";
					when "10110101001101000" => rgb <= "101010";
					when "10110101001101001" => rgb <= "111111";
					when "10110101001101010" => rgb <= "101010";
					when "10110101001101011" => rgb <= "111111";
					when "10110101001101100" => rgb <= "101010";
					when "10110101001101101" => rgb <= "101010";
					when "10110101001101110" => rgb <= "000000";
					when "10110101001101111" => rgb <= "000000";
					when "10110101001110000" => rgb <= "000000";
					when "10110101001110001" => rgb <= "000000";
					when "10110101001110010" => rgb <= "000000";
					when "10110101001110011" => rgb <= "000000";
					when "10110101001110100" => rgb <= "000000";
					when "10110101001110101" => rgb <= "000000";
					when "10110101001110110" => rgb <= "000000";
					when "10110101001110111" => rgb <= "000000";
					when "10110101001111000" => rgb <= "000000";
					when "10110101001111001" => rgb <= "000000";
					when "10110101001111010" => rgb <= "000000";
					when "10110101001111011" => rgb <= "000000";
					when "10110101001111100" => rgb <= "000000";
					when "10110101001111101" => rgb <= "101010";
					when "10110101001111110" => rgb <= "111111";
					when "10110101001111111" => rgb <= "111111";
					when "10110101010000000" => rgb <= "111111";
					when "10110101010000001" => rgb <= "111111";
					when "10110101010000010" => rgb <= "111111";
					when "10110101010000011" => rgb <= "111111";
					when "10110101010000100" => rgb <= "111111";
					when "10110101010000101" => rgb <= "111111";
					when "10110101010000110" => rgb <= "111111";
					when "10110101010000111" => rgb <= "111111";
					when "10110101010001000" => rgb <= "111111";
					when "10110101010001001" => rgb <= "111111";
					when "10110101010001010" => rgb <= "111111";
					when "10110101010001011" => rgb <= "101010";
					when "10110101010001100" => rgb <= "000000";
					when "10110101010001101" => rgb <= "000000";
					when "10110101010001110" => rgb <= "000000";
					when "10110101010001111" => rgb <= "000000";
					when "10110101010010000" => rgb <= "000000";
					when "10110101010010001" => rgb <= "000000";
					when "10110101010010010" => rgb <= "000000";
					when "10110101010010011" => rgb <= "000000";
					when "10110101010010100" => rgb <= "000000";
					when "10110101010010101" => rgb <= "000000";
					when "10110101010010110" => rgb <= "000000";
					when "10110101010010111" => rgb <= "000000";
					when "10110101010011000" => rgb <= "000000";
					when "10110101010011001" => rgb <= "000000";
					when "10110101010011010" => rgb <= "000000";
					when "10110101010011011" => rgb <= "000000";
					when "10110101010011100" => rgb <= "000000";
					when "10110101010011101" => rgb <= "000000";
					when "10110101010011110" => rgb <= "000000";
					when "10110101010011111" => rgb <= "000000";
					when "10110101010100000" => rgb <= "000000";
					when "10110101010100001" => rgb <= "000000";
					when "10110101010100010" => rgb <= "010101";
					when "10110101010100011" => rgb <= "111111";
					when "10110101010100100" => rgb <= "101010";
					when "10110101010100101" => rgb <= "111111";
					when "10110101010100110" => rgb <= "111111";
					when "10110101010100111" => rgb <= "111111";
					when "10110101010101000" => rgb <= "111111";
					when "10110101010101001" => rgb <= "111111";
					when "10110101010101010" => rgb <= "000000";
					when "10110101010101011" => rgb <= "000000";
					when "10110101010101100" => rgb <= "000000";
					when "10110101010101101" => rgb <= "000000";
					when "10110101010101110" => rgb <= "000000";
					when "10110101010101111" => rgb <= "000000";
					when "10110101010110000" => rgb <= "000000";
					when "10110101010110001" => rgb <= "000000";
					when "10110101010110010" => rgb <= "000000";
					when "10110101010110011" => rgb <= "000000";
					when "10110101010110100" => rgb <= "000000";
					when "10110101010110101" => rgb <= "000000";
					when "10110101010110110" => rgb <= "000000";
					when "10110101010110111" => rgb <= "000000";
					when "10110101010111000" => rgb <= "000000";
					when "10110101010111001" => rgb <= "000000";
					when "10110101010111010" => rgb <= "000000";
					when "10110101010111011" => rgb <= "000000";
					when "10110101010111100" => rgb <= "000000";
					when "10110101010111101" => rgb <= "000000";
					when "10110101010111110" => rgb <= "000000";
					when "10110101010111111" => rgb <= "000000";
					when "10110101011000000" => rgb <= "010101";
					when "10110101011000001" => rgb <= "101010";
					when "10110101011000010" => rgb <= "101010";
					when "10110101011000011" => rgb <= "111111";
					when "10110101011000100" => rgb <= "111111";
					when "10110101011000101" => rgb <= "111111";
					when "10110101011000110" => rgb <= "111111";
					when "10110101011000111" => rgb <= "111111";
					when "10110101011001000" => rgb <= "111111";
					when "10110101011001001" => rgb <= "111111";
					when "10110101011001010" => rgb <= "111111";
					when "10110101011001011" => rgb <= "101010";
					when "10110101011001100" => rgb <= "111111";
					when "10110101011001101" => rgb <= "101010";
					when "10110101011001110" => rgb <= "111111";
					when "10110101011001111" => rgb <= "101010";
					when "10110101011010000" => rgb <= "000000";
					when "10110101011010001" => rgb <= "000000";
					when "10110101011010010" => rgb <= "000000";
					when "10110101011010011" => rgb <= "000000";
					when "10110101011010100" => rgb <= "000000";
					when "10110101011010101" => rgb <= "000000";
					when "10110101011010110" => rgb <= "000000";
					when "10110101011010111" => rgb <= "101010";
					when "10110101011011000" => rgb <= "101010";
					when "10110101011011001" => rgb <= "101010";
					when "10110101011011010" => rgb <= "101010";
					when "10110101011011011" => rgb <= "111111";
					when "10110101011011100" => rgb <= "111111";
					when "10110101011011101" => rgb <= "111111";
					when "10110101011011110" => rgb <= "111111";
					when "10110101011011111" => rgb <= "111111";
					when "10110101011100000" => rgb <= "111111";
					when "10110101011100001" => rgb <= "111111";
					when "10110101011100010" => rgb <= "111111";
					when "10110101011100011" => rgb <= "101010";
					when "10110101011100100" => rgb <= "111111";
					when "10110101011100101" => rgb <= "111111";
					when "10110101011100110" => rgb <= "000000";
					when "10110101011100111" => rgb <= "000000";
					when "10110101011101000" => rgb <= "000000";
					when "10110101011101001" => rgb <= "000000";
					when "10110101011101010" => rgb <= "000000";
					when "10110101011101011" => rgb <= "000000";
					when "10110101011101100" => rgb <= "000000";
					when "10110101011101101" => rgb <= "010101";
					when "10110101011101110" => rgb <= "111111";
					when "10110101011101111" => rgb <= "101010";
					when "10110101011110000" => rgb <= "111111";
					when "10110101011110001" => rgb <= "111111";
					when "10110101011110010" => rgb <= "101010";
					when "10110101011110011" => rgb <= "111111";
					when "10110101011110100" => rgb <= "101010";
					when "10110101011110101" => rgb <= "000000";
					when "10110101011110110" => rgb <= "000000";
					when "10110101011110111" => rgb <= "000000";
					when "10110101011111000" => rgb <= "000000";
					when "10110101011111001" => rgb <= "000000";
					when "10110101011111010" => rgb <= "000000";
					when "10110101011111011" => rgb <= "000000";
					when "10110101011111100" => rgb <= "010101";
					when "10110101011111101" => rgb <= "111111";
					when "10110101011111110" => rgb <= "101010";
					when "10110101011111111" => rgb <= "101010";
					when "10110101100000000" => rgb <= "101010";
					when "10110101100000001" => rgb <= "101010";
					when "10110101100000010" => rgb <= "111111";
					when "10110101100000011" => rgb <= "101010";
					when "10110101100000100" => rgb <= "000000";
					when "10110101100000101" => rgb <= "000000";
					when "10110101100000110" => rgb <= "000000";
					when "10110101100000111" => rgb <= "000000";
					when "10110101100001000" => rgb <= "000000";
					when "10110101100001001" => rgb <= "000000";
					when "10110101100001010" => rgb <= "000000";
					when "10110101100001011" => rgb <= "010101";
					when "10110101100001100" => rgb <= "101010";
					when "10110101100001101" => rgb <= "101010";
					when "10110101100001110" => rgb <= "101010";
					when "10110101100001111" => rgb <= "111111";
					when "10110101100010000" => rgb <= "111111";
					when "10110101100010001" => rgb <= "111111";
					when "10110101100010010" => rgb <= "111111";
					when "10110101100010011" => rgb <= "111111";
					when "10110101100010100" => rgb <= "111111";
					when "10110101100010101" => rgb <= "111111";
					when "10110101100010110" => rgb <= "111111";
					when "10110101100010111" => rgb <= "111111";
					when "10110101100011000" => rgb <= "101010";
					when "10110101100011001" => rgb <= "111111";
					when "10110101100011010" => rgb <= "101010";
					when "10110101100011011" => rgb <= "000000";
					when "10110101100011100" => rgb <= "000000";
					when "10110101100011101" => rgb <= "000000";
					when "10110101100011110" => rgb <= "000000";
					when "10110101100011111" => rgb <= "000000";
					when "10110101100100000" => rgb <= "000000";
					when "10110101100100001" => rgb <= "000000";
					when "10110101100100010" => rgb <= "101010";
					when "10110101100100011" => rgb <= "101010";
					when "10110101100100100" => rgb <= "101010";
					when "10110101100100101" => rgb <= "111111";
					when "10110101100100110" => rgb <= "111111";
					when "10110101100100111" => rgb <= "111111";
					when "10110101100101000" => rgb <= "111111";
					when "10110101100101001" => rgb <= "111111";
					when "10110101100101010" => rgb <= "111111";
					when "10110101100101011" => rgb <= "111111";
					when "10110101100101100" => rgb <= "111111";
					when "10110101100101101" => rgb <= "111111";
					when "10110101100101110" => rgb <= "101010";
					when "10110101100101111" => rgb <= "101010";
					when "10110101100110000" => rgb <= "111111";
					when "10110101100110001" => rgb <= "010101";
					when "10110101100110010" => rgb <= "000000";
					when "10110101100110011" => rgb <= "000000";
					when "10110101100110100" => rgb <= "000000";
					when "10110101100110101" => rgb <= "000000";
					when "10110101100110110" => rgb <= "000000";
					when "10110101100110111" => rgb <= "000000";
					when "10110101100111000" => rgb <= "000000";
					when "10110101100111001" => rgb <= "000000";
					when "10110101100111010" => rgb <= "000000";
					when "10110101100111011" => rgb <= "000000";
					when "10110101100111100" => rgb <= "000000";
					when "10110101100111101" => rgb <= "000000";
					when "10110101100111110" => rgb <= "000000";
					when "10110101100111111" => rgb <= "000000";
					when "10110110000000000" => rgb <= "000000";
					when "10110110000000001" => rgb <= "000000";
					when "10110110000000010" => rgb <= "000000";
					when "10110110000000011" => rgb <= "000000";
					when "10110110000000100" => rgb <= "000000";
					when "10110110000000101" => rgb <= "101010";
					when "10110110000000110" => rgb <= "111111";
					when "10110110000000111" => rgb <= "111111";
					when "10110110000001000" => rgb <= "101010";
					when "10110110000001001" => rgb <= "111111";
					when "10110110000001010" => rgb <= "101010";
					when "10110110000001011" => rgb <= "111111";
					when "10110110000001100" => rgb <= "010101";
					when "10110110000001101" => rgb <= "000000";
					when "10110110000001110" => rgb <= "000000";
					when "10110110000001111" => rgb <= "000000";
					when "10110110000010000" => rgb <= "000000";
					when "10110110000010001" => rgb <= "000000";
					when "10110110000010010" => rgb <= "000000";
					when "10110110000010011" => rgb <= "000000";
					when "10110110000010100" => rgb <= "000000";
					when "10110110000010101" => rgb <= "000000";
					when "10110110000010110" => rgb <= "000000";
					when "10110110000010111" => rgb <= "000000";
					when "10110110000011000" => rgb <= "000000";
					when "10110110000011001" => rgb <= "000000";
					when "10110110000011010" => rgb <= "000000";
					when "10110110000011011" => rgb <= "010101";
					when "10110110000011100" => rgb <= "101010";
					when "10110110000011101" => rgb <= "111111";
					when "10110110000011110" => rgb <= "111111";
					when "10110110000011111" => rgb <= "101010";
					when "10110110000100000" => rgb <= "111111";
					when "10110110000100001" => rgb <= "111111";
					when "10110110000100010" => rgb <= "111111";
					when "10110110000100011" => rgb <= "111111";
					when "10110110000100100" => rgb <= "111111";
					when "10110110000100101" => rgb <= "111111";
					when "10110110000100110" => rgb <= "101010";
					when "10110110000100111" => rgb <= "101010";
					when "10110110000101000" => rgb <= "101010";
					when "10110110000101001" => rgb <= "101010";
					when "10110110000101010" => rgb <= "111111";
					when "10110110000101011" => rgb <= "101010";
					when "10110110000101100" => rgb <= "111111";
					when "10110110000101101" => rgb <= "101010";
					when "10110110000101110" => rgb <= "101010";
					when "10110110000101111" => rgb <= "111111";
					when "10110110000110000" => rgb <= "111111";
					when "10110110000110001" => rgb <= "101010";
					when "10110110000110010" => rgb <= "000000";
					when "10110110000110011" => rgb <= "000000";
					when "10110110000110100" => rgb <= "000000";
					when "10110110000110101" => rgb <= "000000";
					when "10110110000110110" => rgb <= "000000";
					when "10110110000110111" => rgb <= "000000";
					when "10110110000111000" => rgb <= "000000";
					when "10110110000111001" => rgb <= "010101";
					when "10110110000111010" => rgb <= "111111";
					when "10110110000111011" => rgb <= "101010";
					when "10110110000111100" => rgb <= "111111";
					when "10110110000111101" => rgb <= "111111";
					when "10110110000111110" => rgb <= "111111";
					when "10110110000111111" => rgb <= "111111";
					when "10110110001000000" => rgb <= "101010";
					when "10110110001000001" => rgb <= "000000";
					when "10110110001000010" => rgb <= "000000";
					when "10110110001000011" => rgb <= "000000";
					when "10110110001000100" => rgb <= "000000";
					when "10110110001000101" => rgb <= "000000";
					when "10110110001000110" => rgb <= "000000";
					when "10110110001000111" => rgb <= "000000";
					when "10110110001001000" => rgb <= "000000";
					when "10110110001001001" => rgb <= "000000";
					when "10110110001001010" => rgb <= "000000";
					when "10110110001001011" => rgb <= "000000";
					when "10110110001001100" => rgb <= "000000";
					when "10110110001001101" => rgb <= "000000";
					when "10110110001001110" => rgb <= "000000";
					when "10110110001001111" => rgb <= "000000";
					when "10110110001010000" => rgb <= "101010";
					when "10110110001010001" => rgb <= "101010";
					when "10110110001010010" => rgb <= "101010";
					when "10110110001010011" => rgb <= "101010";
					when "10110110001010100" => rgb <= "111111";
					when "10110110001010101" => rgb <= "111111";
					when "10110110001010110" => rgb <= "111111";
					when "10110110001010111" => rgb <= "111111";
					when "10110110001011000" => rgb <= "111111";
					when "10110110001011001" => rgb <= "111111";
					when "10110110001011010" => rgb <= "111111";
					when "10110110001011011" => rgb <= "101010";
					when "10110110001011100" => rgb <= "111111";
					when "10110110001011101" => rgb <= "101010";
					when "10110110001011110" => rgb <= "101010";
					when "10110110001011111" => rgb <= "000000";
					when "10110110001100000" => rgb <= "000000";
					when "10110110001100001" => rgb <= "000000";
					when "10110110001100010" => rgb <= "000000";
					when "10110110001100011" => rgb <= "000000";
					when "10110110001100100" => rgb <= "000000";
					when "10110110001100101" => rgb <= "000000";
					when "10110110001100110" => rgb <= "010101";
					when "10110110001100111" => rgb <= "101010";
					when "10110110001101000" => rgb <= "101010";
					when "10110110001101001" => rgb <= "111111";
					when "10110110001101010" => rgb <= "101010";
					when "10110110001101011" => rgb <= "111111";
					when "10110110001101100" => rgb <= "101010";
					when "10110110001101101" => rgb <= "101010";
					when "10110110001101110" => rgb <= "000000";
					when "10110110001101111" => rgb <= "000000";
					when "10110110001110000" => rgb <= "000000";
					when "10110110001110001" => rgb <= "000000";
					when "10110110001110010" => rgb <= "000000";
					when "10110110001110011" => rgb <= "000000";
					when "10110110001110100" => rgb <= "000000";
					when "10110110001110101" => rgb <= "000000";
					when "10110110001110110" => rgb <= "000000";
					when "10110110001110111" => rgb <= "000000";
					when "10110110001111000" => rgb <= "000000";
					when "10110110001111001" => rgb <= "000000";
					when "10110110001111010" => rgb <= "000000";
					when "10110110001111011" => rgb <= "000000";
					when "10110110001111100" => rgb <= "000000";
					when "10110110001111101" => rgb <= "101010";
					when "10110110001111110" => rgb <= "111111";
					when "10110110001111111" => rgb <= "111111";
					when "10110110010000000" => rgb <= "111111";
					when "10110110010000001" => rgb <= "111111";
					when "10110110010000010" => rgb <= "111111";
					when "10110110010000011" => rgb <= "111111";
					when "10110110010000100" => rgb <= "111111";
					when "10110110010000101" => rgb <= "111111";
					when "10110110010000110" => rgb <= "111111";
					when "10110110010000111" => rgb <= "111111";
					when "10110110010001000" => rgb <= "111111";
					when "10110110010001001" => rgb <= "111111";
					when "10110110010001010" => rgb <= "111111";
					when "10110110010001011" => rgb <= "101010";
					when "10110110010001100" => rgb <= "000000";
					when "10110110010001101" => rgb <= "000000";
					when "10110110010001110" => rgb <= "000000";
					when "10110110010001111" => rgb <= "000000";
					when "10110110010010000" => rgb <= "000000";
					when "10110110010010001" => rgb <= "000000";
					when "10110110010010010" => rgb <= "000000";
					when "10110110010010011" => rgb <= "000000";
					when "10110110010010100" => rgb <= "000000";
					when "10110110010010101" => rgb <= "000000";
					when "10110110010010110" => rgb <= "000000";
					when "10110110010010111" => rgb <= "000000";
					when "10110110010011000" => rgb <= "000000";
					when "10110110010011001" => rgb <= "000000";
					when "10110110010011010" => rgb <= "000000";
					when "10110110010011011" => rgb <= "000000";
					when "10110110010011100" => rgb <= "000000";
					when "10110110010011101" => rgb <= "000000";
					when "10110110010011110" => rgb <= "000000";
					when "10110110010011111" => rgb <= "000000";
					when "10110110010100000" => rgb <= "000000";
					when "10110110010100001" => rgb <= "000000";
					when "10110110010100010" => rgb <= "010101";
					when "10110110010100011" => rgb <= "111111";
					when "10110110010100100" => rgb <= "101010";
					when "10110110010100101" => rgb <= "111111";
					when "10110110010100110" => rgb <= "111111";
					when "10110110010100111" => rgb <= "111111";
					when "10110110010101000" => rgb <= "111111";
					when "10110110010101001" => rgb <= "111111";
					when "10110110010101010" => rgb <= "000000";
					when "10110110010101011" => rgb <= "000000";
					when "10110110010101100" => rgb <= "000000";
					when "10110110010101101" => rgb <= "000000";
					when "10110110010101110" => rgb <= "000000";
					when "10110110010101111" => rgb <= "000000";
					when "10110110010110000" => rgb <= "000000";
					when "10110110010110001" => rgb <= "000000";
					when "10110110010110010" => rgb <= "000000";
					when "10110110010110011" => rgb <= "000000";
					when "10110110010110100" => rgb <= "000000";
					when "10110110010110101" => rgb <= "000000";
					when "10110110010110110" => rgb <= "000000";
					when "10110110010110111" => rgb <= "000000";
					when "10110110010111000" => rgb <= "000000";
					when "10110110010111001" => rgb <= "000000";
					when "10110110010111010" => rgb <= "000000";
					when "10110110010111011" => rgb <= "000000";
					when "10110110010111100" => rgb <= "000000";
					when "10110110010111101" => rgb <= "000000";
					when "10110110010111110" => rgb <= "000000";
					when "10110110010111111" => rgb <= "000000";
					when "10110110011000000" => rgb <= "010101";
					when "10110110011000001" => rgb <= "101010";
					when "10110110011000010" => rgb <= "101010";
					when "10110110011000011" => rgb <= "111111";
					when "10110110011000100" => rgb <= "111111";
					when "10110110011000101" => rgb <= "111111";
					when "10110110011000110" => rgb <= "111111";
					when "10110110011000111" => rgb <= "111111";
					when "10110110011001000" => rgb <= "111111";
					when "10110110011001001" => rgb <= "111111";
					when "10110110011001010" => rgb <= "111111";
					when "10110110011001011" => rgb <= "101010";
					when "10110110011001100" => rgb <= "111111";
					when "10110110011001101" => rgb <= "101010";
					when "10110110011001110" => rgb <= "111111";
					when "10110110011001111" => rgb <= "101010";
					when "10110110011010000" => rgb <= "000000";
					when "10110110011010001" => rgb <= "000000";
					when "10110110011010010" => rgb <= "000000";
					when "10110110011010011" => rgb <= "000000";
					when "10110110011010100" => rgb <= "000000";
					when "10110110011010101" => rgb <= "000000";
					when "10110110011010110" => rgb <= "000000";
					when "10110110011010111" => rgb <= "101010";
					when "10110110011011000" => rgb <= "101010";
					when "10110110011011001" => rgb <= "101010";
					when "10110110011011010" => rgb <= "101010";
					when "10110110011011011" => rgb <= "111111";
					when "10110110011011100" => rgb <= "111111";
					when "10110110011011101" => rgb <= "111111";
					when "10110110011011110" => rgb <= "111111";
					when "10110110011011111" => rgb <= "111111";
					when "10110110011100000" => rgb <= "111111";
					when "10110110011100001" => rgb <= "111111";
					when "10110110011100010" => rgb <= "111111";
					when "10110110011100011" => rgb <= "101010";
					when "10110110011100100" => rgb <= "111111";
					when "10110110011100101" => rgb <= "111111";
					when "10110110011100110" => rgb <= "000000";
					when "10110110011100111" => rgb <= "000000";
					when "10110110011101000" => rgb <= "000000";
					when "10110110011101001" => rgb <= "000000";
					when "10110110011101010" => rgb <= "000000";
					when "10110110011101011" => rgb <= "000000";
					when "10110110011101100" => rgb <= "000000";
					when "10110110011101101" => rgb <= "010101";
					when "10110110011101110" => rgb <= "111111";
					when "10110110011101111" => rgb <= "101010";
					when "10110110011110000" => rgb <= "111111";
					when "10110110011110001" => rgb <= "111111";
					when "10110110011110010" => rgb <= "111111";
					when "10110110011110011" => rgb <= "111111";
					when "10110110011110100" => rgb <= "101010";
					when "10110110011110101" => rgb <= "000000";
					when "10110110011110110" => rgb <= "000000";
					when "10110110011110111" => rgb <= "000000";
					when "10110110011111000" => rgb <= "000000";
					when "10110110011111001" => rgb <= "000000";
					when "10110110011111010" => rgb <= "000000";
					when "10110110011111011" => rgb <= "000000";
					when "10110110011111100" => rgb <= "010101";
					when "10110110011111101" => rgb <= "101010";
					when "10110110011111110" => rgb <= "111111";
					when "10110110011111111" => rgb <= "111111";
					when "10110110100000000" => rgb <= "111111";
					when "10110110100000001" => rgb <= "111111";
					when "10110110100000010" => rgb <= "111111";
					when "10110110100000011" => rgb <= "101010";
					when "10110110100000100" => rgb <= "000000";
					when "10110110100000101" => rgb <= "000000";
					when "10110110100000110" => rgb <= "000000";
					when "10110110100000111" => rgb <= "000000";
					when "10110110100001000" => rgb <= "000000";
					when "10110110100001001" => rgb <= "000000";
					when "10110110100001010" => rgb <= "000000";
					when "10110110100001011" => rgb <= "010101";
					when "10110110100001100" => rgb <= "101010";
					when "10110110100001101" => rgb <= "111111";
					when "10110110100001110" => rgb <= "111111";
					when "10110110100001111" => rgb <= "101010";
					when "10110110100010000" => rgb <= "111111";
					when "10110110100010001" => rgb <= "111111";
					when "10110110100010010" => rgb <= "111111";
					when "10110110100010011" => rgb <= "111111";
					when "10110110100010100" => rgb <= "111111";
					when "10110110100010101" => rgb <= "111111";
					when "10110110100010110" => rgb <= "111111";
					when "10110110100010111" => rgb <= "111111";
					when "10110110100011000" => rgb <= "101010";
					when "10110110100011001" => rgb <= "111111";
					when "10110110100011010" => rgb <= "101010";
					when "10110110100011011" => rgb <= "000000";
					when "10110110100011100" => rgb <= "000000";
					when "10110110100011101" => rgb <= "000000";
					when "10110110100011110" => rgb <= "000000";
					when "10110110100011111" => rgb <= "000000";
					when "10110110100100000" => rgb <= "000000";
					when "10110110100100001" => rgb <= "000000";
					when "10110110100100010" => rgb <= "101010";
					when "10110110100100011" => rgb <= "101010";
					when "10110110100100100" => rgb <= "101010";
					when "10110110100100101" => rgb <= "111111";
					when "10110110100100110" => rgb <= "111111";
					when "10110110100100111" => rgb <= "111111";
					when "10110110100101000" => rgb <= "111111";
					when "10110110100101001" => rgb <= "111111";
					when "10110110100101010" => rgb <= "111111";
					when "10110110100101011" => rgb <= "111111";
					when "10110110100101100" => rgb <= "111111";
					when "10110110100101101" => rgb <= "111111";
					when "10110110100101110" => rgb <= "101010";
					when "10110110100101111" => rgb <= "101010";
					when "10110110100110000" => rgb <= "111111";
					when "10110110100110001" => rgb <= "010101";
					when "10110110100110010" => rgb <= "000000";
					when "10110110100110011" => rgb <= "000000";
					when "10110110100110100" => rgb <= "000000";
					when "10110110100110101" => rgb <= "000000";
					when "10110110100110110" => rgb <= "000000";
					when "10110110100110111" => rgb <= "000000";
					when "10110110100111000" => rgb <= "000000";
					when "10110110100111001" => rgb <= "000000";
					when "10110110100111010" => rgb <= "000000";
					when "10110110100111011" => rgb <= "000000";
					when "10110110100111100" => rgb <= "000000";
					when "10110110100111101" => rgb <= "000000";
					when "10110110100111110" => rgb <= "000000";
					when "10110110100111111" => rgb <= "000000";
					when "10110111000000000" => rgb <= "000000";
					when "10110111000000001" => rgb <= "000000";
					when "10110111000000010" => rgb <= "000000";
					when "10110111000000011" => rgb <= "000000";
					when "10110111000000100" => rgb <= "000000";
					when "10110111000000101" => rgb <= "010101";
					when "10110111000000110" => rgb <= "010101";
					when "10110111000000111" => rgb <= "010101";
					when "10110111000001000" => rgb <= "010101";
					when "10110111000001001" => rgb <= "010101";
					when "10110111000001010" => rgb <= "010101";
					when "10110111000001011" => rgb <= "010101";
					when "10110111000001100" => rgb <= "010101";
					when "10110111000001101" => rgb <= "010101";
					when "10110111000001110" => rgb <= "010101";
					when "10110111000001111" => rgb <= "010101";
					when "10110111000010000" => rgb <= "010101";
					when "10110111000010001" => rgb <= "010101";
					when "10110111000010010" => rgb <= "010101";
					when "10110111000010011" => rgb <= "010101";
					when "10110111000010100" => rgb <= "010101";
					when "10110111000010101" => rgb <= "010101";
					when "10110111000010110" => rgb <= "010101";
					when "10110111000010111" => rgb <= "010101";
					when "10110111000011000" => rgb <= "010101";
					when "10110111000011001" => rgb <= "010101";
					when "10110111000011010" => rgb <= "010101";
					when "10110111000011011" => rgb <= "101010";
					when "10110111000011100" => rgb <= "111111";
					when "10110111000011101" => rgb <= "101010";
					when "10110111000011110" => rgb <= "111111";
					when "10110111000011111" => rgb <= "111111";
					when "10110111000100000" => rgb <= "111111";
					when "10110111000100001" => rgb <= "111111";
					when "10110111000100010" => rgb <= "111111";
					when "10110111000100011" => rgb <= "111111";
					when "10110111000100100" => rgb <= "111111";
					when "10110111000100101" => rgb <= "111111";
					when "10110111000100110" => rgb <= "111111";
					when "10110111000100111" => rgb <= "111111";
					when "10110111000101000" => rgb <= "101010";
					when "10110111000101001" => rgb <= "101010";
					when "10110111000101010" => rgb <= "101010";
					when "10110111000101011" => rgb <= "010101";
					when "10110111000101100" => rgb <= "010101";
					when "10110111000101101" => rgb <= "010101";
					when "10110111000101110" => rgb <= "010101";
					when "10110111000101111" => rgb <= "010101";
					when "10110111000110000" => rgb <= "010101";
					when "10110111000110001" => rgb <= "010101";
					when "10110111000110010" => rgb <= "000000";
					when "10110111000110011" => rgb <= "000000";
					when "10110111000110100" => rgb <= "000000";
					when "10110111000110101" => rgb <= "000000";
					when "10110111000110110" => rgb <= "000000";
					when "10110111000110111" => rgb <= "000000";
					when "10110111000111000" => rgb <= "000000";
					when "10110111000111001" => rgb <= "010101";
					when "10110111000111010" => rgb <= "111111";
					when "10110111000111011" => rgb <= "101010";
					when "10110111000111100" => rgb <= "111111";
					when "10110111000111101" => rgb <= "111111";
					when "10110111000111110" => rgb <= "111111";
					when "10110111000111111" => rgb <= "111111";
					when "10110111001000000" => rgb <= "101010";
					when "10110111001000001" => rgb <= "000000";
					when "10110111001000010" => rgb <= "000000";
					when "10110111001000011" => rgb <= "000000";
					when "10110111001000100" => rgb <= "000000";
					when "10110111001000101" => rgb <= "000000";
					when "10110111001000110" => rgb <= "000000";
					when "10110111001000111" => rgb <= "000000";
					when "10110111001001000" => rgb <= "000000";
					when "10110111001001001" => rgb <= "000000";
					when "10110111001001010" => rgb <= "000000";
					when "10110111001001011" => rgb <= "000000";
					when "10110111001001100" => rgb <= "000000";
					when "10110111001001101" => rgb <= "000000";
					when "10110111001001110" => rgb <= "000000";
					when "10110111001001111" => rgb <= "000000";
					when "10110111001010000" => rgb <= "101010";
					when "10110111001010001" => rgb <= "101010";
					when "10110111001010010" => rgb <= "101010";
					when "10110111001010011" => rgb <= "101010";
					when "10110111001010100" => rgb <= "111111";
					when "10110111001010101" => rgb <= "111111";
					when "10110111001010110" => rgb <= "111111";
					when "10110111001010111" => rgb <= "111111";
					when "10110111001011000" => rgb <= "111111";
					when "10110111001011001" => rgb <= "111111";
					when "10110111001011010" => rgb <= "111111";
					when "10110111001011011" => rgb <= "101010";
					when "10110111001011100" => rgb <= "111111";
					when "10110111001011101" => rgb <= "101010";
					when "10110111001011110" => rgb <= "101010";
					when "10110111001011111" => rgb <= "000000";
					when "10110111001100000" => rgb <= "000000";
					when "10110111001100001" => rgb <= "000000";
					when "10110111001100010" => rgb <= "000000";
					when "10110111001100011" => rgb <= "000000";
					when "10110111001100100" => rgb <= "000000";
					when "10110111001100101" => rgb <= "000000";
					when "10110111001100110" => rgb <= "010101";
					when "10110111001100111" => rgb <= "111111";
					when "10110111001101000" => rgb <= "101010";
					when "10110111001101001" => rgb <= "111111";
					when "10110111001101010" => rgb <= "101010";
					when "10110111001101011" => rgb <= "111111";
					when "10110111001101100" => rgb <= "101010";
					when "10110111001101101" => rgb <= "101010";
					when "10110111001101110" => rgb <= "000000";
					when "10110111001101111" => rgb <= "000000";
					when "10110111001110000" => rgb <= "000000";
					when "10110111001110001" => rgb <= "000000";
					when "10110111001110010" => rgb <= "000000";
					when "10110111001110011" => rgb <= "000000";
					when "10110111001110100" => rgb <= "000000";
					when "10110111001110101" => rgb <= "000000";
					when "10110111001110110" => rgb <= "000000";
					when "10110111001110111" => rgb <= "000000";
					when "10110111001111000" => rgb <= "000000";
					when "10110111001111001" => rgb <= "000000";
					when "10110111001111010" => rgb <= "000000";
					when "10110111001111011" => rgb <= "000000";
					when "10110111001111100" => rgb <= "000000";
					when "10110111001111101" => rgb <= "101010";
					when "10110111001111110" => rgb <= "111111";
					when "10110111001111111" => rgb <= "111111";
					when "10110111010000000" => rgb <= "111111";
					when "10110111010000001" => rgb <= "111111";
					when "10110111010000010" => rgb <= "111111";
					when "10110111010000011" => rgb <= "111111";
					when "10110111010000100" => rgb <= "111111";
					when "10110111010000101" => rgb <= "111111";
					when "10110111010000110" => rgb <= "111111";
					when "10110111010000111" => rgb <= "111111";
					when "10110111010001000" => rgb <= "111111";
					when "10110111010001001" => rgb <= "111111";
					when "10110111010001010" => rgb <= "111111";
					when "10110111010001011" => rgb <= "101010";
					when "10110111010001100" => rgb <= "000000";
					when "10110111010001101" => rgb <= "000000";
					when "10110111010001110" => rgb <= "000000";
					when "10110111010001111" => rgb <= "000000";
					when "10110111010010000" => rgb <= "000000";
					when "10110111010010001" => rgb <= "000000";
					when "10110111010010010" => rgb <= "000000";
					when "10110111010010011" => rgb <= "000000";
					when "10110111010010100" => rgb <= "000000";
					when "10110111010010101" => rgb <= "000000";
					when "10110111010010110" => rgb <= "000000";
					when "10110111010010111" => rgb <= "000000";
					when "10110111010011000" => rgb <= "000000";
					when "10110111010011001" => rgb <= "000000";
					when "10110111010011010" => rgb <= "000000";
					when "10110111010011011" => rgb <= "000000";
					when "10110111010011100" => rgb <= "000000";
					when "10110111010011101" => rgb <= "000000";
					when "10110111010011110" => rgb <= "000000";
					when "10110111010011111" => rgb <= "000000";
					when "10110111010100000" => rgb <= "000000";
					when "10110111010100001" => rgb <= "000000";
					when "10110111010100010" => rgb <= "010101";
					when "10110111010100011" => rgb <= "111111";
					when "10110111010100100" => rgb <= "101010";
					when "10110111010100101" => rgb <= "111111";
					when "10110111010100110" => rgb <= "111111";
					when "10110111010100111" => rgb <= "111111";
					when "10110111010101000" => rgb <= "111111";
					when "10110111010101001" => rgb <= "111111";
					when "10110111010101010" => rgb <= "000000";
					when "10110111010101011" => rgb <= "000000";
					when "10110111010101100" => rgb <= "000000";
					when "10110111010101101" => rgb <= "000000";
					when "10110111010101110" => rgb <= "000000";
					when "10110111010101111" => rgb <= "000000";
					when "10110111010110000" => rgb <= "000000";
					when "10110111010110001" => rgb <= "000000";
					when "10110111010110010" => rgb <= "010101";
					when "10110111010110011" => rgb <= "010101";
					when "10110111010110100" => rgb <= "010101";
					when "10110111010110101" => rgb <= "010101";
					when "10110111010110110" => rgb <= "010101";
					when "10110111010110111" => rgb <= "010101";
					when "10110111010111000" => rgb <= "010101";
					when "10110111010111001" => rgb <= "000000";
					when "10110111010111010" => rgb <= "000000";
					when "10110111010111011" => rgb <= "000000";
					when "10110111010111100" => rgb <= "000000";
					when "10110111010111101" => rgb <= "000000";
					when "10110111010111110" => rgb <= "000000";
					when "10110111010111111" => rgb <= "000000";
					when "10110111011000000" => rgb <= "010101";
					when "10110111011000001" => rgb <= "101010";
					when "10110111011000010" => rgb <= "101010";
					when "10110111011000011" => rgb <= "111111";
					when "10110111011000100" => rgb <= "111111";
					when "10110111011000101" => rgb <= "111111";
					when "10110111011000110" => rgb <= "111111";
					when "10110111011000111" => rgb <= "111111";
					when "10110111011001000" => rgb <= "111111";
					when "10110111011001001" => rgb <= "111111";
					when "10110111011001010" => rgb <= "111111";
					when "10110111011001011" => rgb <= "101010";
					when "10110111011001100" => rgb <= "111111";
					when "10110111011001101" => rgb <= "101010";
					when "10110111011001110" => rgb <= "111111";
					when "10110111011001111" => rgb <= "101010";
					when "10110111011010000" => rgb <= "000000";
					when "10110111011010001" => rgb <= "000000";
					when "10110111011010010" => rgb <= "000000";
					when "10110111011010011" => rgb <= "000000";
					when "10110111011010100" => rgb <= "000000";
					when "10110111011010101" => rgb <= "000000";
					when "10110111011010110" => rgb <= "000000";
					when "10110111011010111" => rgb <= "101010";
					when "10110111011011000" => rgb <= "101010";
					when "10110111011011001" => rgb <= "101010";
					when "10110111011011010" => rgb <= "101010";
					when "10110111011011011" => rgb <= "111111";
					when "10110111011011100" => rgb <= "111111";
					when "10110111011011101" => rgb <= "111111";
					when "10110111011011110" => rgb <= "111111";
					when "10110111011011111" => rgb <= "111111";
					when "10110111011100000" => rgb <= "111111";
					when "10110111011100001" => rgb <= "111111";
					when "10110111011100010" => rgb <= "111111";
					when "10110111011100011" => rgb <= "101010";
					when "10110111011100100" => rgb <= "111111";
					when "10110111011100101" => rgb <= "111111";
					when "10110111011100110" => rgb <= "000000";
					when "10110111011100111" => rgb <= "000000";
					when "10110111011101000" => rgb <= "000000";
					when "10110111011101001" => rgb <= "000000";
					when "10110111011101010" => rgb <= "000000";
					when "10110111011101011" => rgb <= "000000";
					when "10110111011101100" => rgb <= "000000";
					when "10110111011101101" => rgb <= "010101";
					when "10110111011101110" => rgb <= "111111";
					when "10110111011101111" => rgb <= "101010";
					when "10110111011110000" => rgb <= "111111";
					when "10110111011110001" => rgb <= "111111";
					when "10110111011110010" => rgb <= "101010";
					when "10110111011110011" => rgb <= "111111";
					when "10110111011110100" => rgb <= "101010";
					when "10110111011110101" => rgb <= "000000";
					when "10110111011110110" => rgb <= "000000";
					when "10110111011110111" => rgb <= "000000";
					when "10110111011111000" => rgb <= "000000";
					when "10110111011111001" => rgb <= "000000";
					when "10110111011111010" => rgb <= "000000";
					when "10110111011111011" => rgb <= "000000";
					when "10110111011111100" => rgb <= "000000";
					when "10110111011111101" => rgb <= "010101";
					when "10110111011111110" => rgb <= "010101";
					when "10110111011111111" => rgb <= "010101";
					when "10110111100000000" => rgb <= "010101";
					when "10110111100000001" => rgb <= "010101";
					when "10110111100000010" => rgb <= "010101";
					when "10110111100000011" => rgb <= "010101";
					when "10110111100000100" => rgb <= "010101";
					when "10110111100000101" => rgb <= "010101";
					when "10110111100000110" => rgb <= "010101";
					when "10110111100000111" => rgb <= "010101";
					when "10110111100001000" => rgb <= "010101";
					when "10110111100001001" => rgb <= "010101";
					when "10110111100001010" => rgb <= "010101";
					when "10110111100001011" => rgb <= "101010";
					when "10110111100001100" => rgb <= "111111";
					when "10110111100001101" => rgb <= "101010";
					when "10110111100001110" => rgb <= "111111";
					when "10110111100001111" => rgb <= "111111";
					when "10110111100010000" => rgb <= "111111";
					when "10110111100010001" => rgb <= "111111";
					when "10110111100010010" => rgb <= "111111";
					when "10110111100010011" => rgb <= "111111";
					when "10110111100010100" => rgb <= "111111";
					when "10110111100010101" => rgb <= "111111";
					when "10110111100010110" => rgb <= "111111";
					when "10110111100010111" => rgb <= "111111";
					when "10110111100011000" => rgb <= "101010";
					when "10110111100011001" => rgb <= "111111";
					when "10110111100011010" => rgb <= "101010";
					when "10110111100011011" => rgb <= "000000";
					when "10110111100011100" => rgb <= "000000";
					when "10110111100011101" => rgb <= "000000";
					when "10110111100011110" => rgb <= "000000";
					when "10110111100011111" => rgb <= "000000";
					when "10110111100100000" => rgb <= "000000";
					when "10110111100100001" => rgb <= "000000";
					when "10110111100100010" => rgb <= "101010";
					when "10110111100100011" => rgb <= "101010";
					when "10110111100100100" => rgb <= "101010";
					when "10110111100100101" => rgb <= "111111";
					when "10110111100100110" => rgb <= "111111";
					when "10110111100100111" => rgb <= "111111";
					when "10110111100101000" => rgb <= "111111";
					when "10110111100101001" => rgb <= "111111";
					when "10110111100101010" => rgb <= "111111";
					when "10110111100101011" => rgb <= "111111";
					when "10110111100101100" => rgb <= "111111";
					when "10110111100101101" => rgb <= "111111";
					when "10110111100101110" => rgb <= "101010";
					when "10110111100101111" => rgb <= "101010";
					when "10110111100110000" => rgb <= "111111";
					when "10110111100110001" => rgb <= "010101";
					when "10110111100110010" => rgb <= "000000";
					when "10110111100110011" => rgb <= "000000";
					when "10110111100110100" => rgb <= "000000";
					when "10110111100110101" => rgb <= "000000";
					when "10110111100110110" => rgb <= "000000";
					when "10110111100110111" => rgb <= "000000";
					when "10110111100111000" => rgb <= "000000";
					when "10110111100111001" => rgb <= "000000";
					when "10110111100111010" => rgb <= "000000";
					when "10110111100111011" => rgb <= "000000";
					when "10110111100111100" => rgb <= "000000";
					when "10110111100111101" => rgb <= "000000";
					when "10110111100111110" => rgb <= "000000";
					when "10110111100111111" => rgb <= "000000";
					when "10111000000000000" => rgb <= "000000";
					when "10111000000000001" => rgb <= "000000";
					when "10111000000000010" => rgb <= "000000";
					when "10111000000000011" => rgb <= "000000";
					when "10111000000000100" => rgb <= "000000";
					when "10111000000000101" => rgb <= "000000";
					when "10111000000000110" => rgb <= "000000";
					when "10111000000000111" => rgb <= "000000";
					when "10111000000001000" => rgb <= "000000";
					when "10111000000001001" => rgb <= "000000";
					when "10111000000001010" => rgb <= "000000";
					when "10111000000001011" => rgb <= "000000";
					when "10111000000001100" => rgb <= "010101";
					when "10111000000001101" => rgb <= "101010";
					when "10111000000001110" => rgb <= "111111";
					when "10111000000001111" => rgb <= "111111";
					when "10111000000010000" => rgb <= "101010";
					when "10111000000010001" => rgb <= "101010";
					when "10111000000010010" => rgb <= "101010";
					when "10111000000010011" => rgb <= "111111";
					when "10111000000010100" => rgb <= "111111";
					when "10111000000010101" => rgb <= "111111";
					when "10111000000010110" => rgb <= "111111";
					when "10111000000010111" => rgb <= "111111";
					when "10111000000011000" => rgb <= "111111";
					when "10111000000011001" => rgb <= "111111";
					when "10111000000011010" => rgb <= "111111";
					when "10111000000011011" => rgb <= "111111";
					when "10111000000011100" => rgb <= "101010";
					when "10111000000011101" => rgb <= "101010";
					when "10111000000011110" => rgb <= "101010";
					when "10111000000011111" => rgb <= "101010";
					when "10111000000100000" => rgb <= "111111";
					when "10111000000100001" => rgb <= "111111";
					when "10111000000100010" => rgb <= "111111";
					when "10111000000100011" => rgb <= "111111";
					when "10111000000100100" => rgb <= "111111";
					when "10111000000100101" => rgb <= "111111";
					when "10111000000100110" => rgb <= "101010";
					when "10111000000100111" => rgb <= "101010";
					when "10111000000101000" => rgb <= "101010";
					when "10111000000101001" => rgb <= "111111";
					when "10111000000101010" => rgb <= "101010";
					when "10111000000101011" => rgb <= "000000";
					when "10111000000101100" => rgb <= "000000";
					when "10111000000101101" => rgb <= "000000";
					when "10111000000101110" => rgb <= "000000";
					when "10111000000101111" => rgb <= "000000";
					when "10111000000110000" => rgb <= "000000";
					when "10111000000110001" => rgb <= "000000";
					when "10111000000110010" => rgb <= "000000";
					when "10111000000110011" => rgb <= "000000";
					when "10111000000110100" => rgb <= "000000";
					when "10111000000110101" => rgb <= "000000";
					when "10111000000110110" => rgb <= "000000";
					when "10111000000110111" => rgb <= "000000";
					when "10111000000111000" => rgb <= "000000";
					when "10111000000111001" => rgb <= "010101";
					when "10111000000111010" => rgb <= "101010";
					when "10111000000111011" => rgb <= "101010";
					when "10111000000111100" => rgb <= "101010";
					when "10111000000111101" => rgb <= "111111";
					when "10111000000111110" => rgb <= "111111";
					when "10111000000111111" => rgb <= "111111";
					when "10111000001000000" => rgb <= "101010";
					when "10111000001000001" => rgb <= "000000";
					when "10111000001000010" => rgb <= "000000";
					when "10111000001000011" => rgb <= "000000";
					when "10111000001000100" => rgb <= "000000";
					when "10111000001000101" => rgb <= "000000";
					when "10111000001000110" => rgb <= "000000";
					when "10111000001000111" => rgb <= "000000";
					when "10111000001001000" => rgb <= "000000";
					when "10111000001001001" => rgb <= "000000";
					when "10111000001001010" => rgb <= "000000";
					when "10111000001001011" => rgb <= "000000";
					when "10111000001001100" => rgb <= "000000";
					when "10111000001001101" => rgb <= "000000";
					when "10111000001001110" => rgb <= "000000";
					when "10111000001001111" => rgb <= "000000";
					when "10111000001010000" => rgb <= "101010";
					when "10111000001010001" => rgb <= "101010";
					when "10111000001010010" => rgb <= "101010";
					when "10111000001010011" => rgb <= "101010";
					when "10111000001010100" => rgb <= "111111";
					when "10111000001010101" => rgb <= "111111";
					when "10111000001010110" => rgb <= "101010";
					when "10111000001010111" => rgb <= "111111";
					when "10111000001011000" => rgb <= "111111";
					when "10111000001011001" => rgb <= "111111";
					when "10111000001011010" => rgb <= "111111";
					when "10111000001011011" => rgb <= "101010";
					when "10111000001011100" => rgb <= "111111";
					when "10111000001011101" => rgb <= "101010";
					when "10111000001011110" => rgb <= "101010";
					when "10111000001011111" => rgb <= "000000";
					when "10111000001100000" => rgb <= "000000";
					when "10111000001100001" => rgb <= "000000";
					when "10111000001100010" => rgb <= "000000";
					when "10111000001100011" => rgb <= "000000";
					when "10111000001100100" => rgb <= "000000";
					when "10111000001100101" => rgb <= "000000";
					when "10111000001100110" => rgb <= "010101";
					when "10111000001100111" => rgb <= "111111";
					when "10111000001101000" => rgb <= "101010";
					when "10111000001101001" => rgb <= "111111";
					when "10111000001101010" => rgb <= "101010";
					when "10111000001101011" => rgb <= "111111";
					when "10111000001101100" => rgb <= "101010";
					when "10111000001101101" => rgb <= "101010";
					when "10111000001101110" => rgb <= "000000";
					when "10111000001101111" => rgb <= "000000";
					when "10111000001110000" => rgb <= "000000";
					when "10111000001110001" => rgb <= "000000";
					when "10111000001110010" => rgb <= "000000";
					when "10111000001110011" => rgb <= "000000";
					when "10111000001110100" => rgb <= "000000";
					when "10111000001110101" => rgb <= "000000";
					when "10111000001110110" => rgb <= "000000";
					when "10111000001110111" => rgb <= "000000";
					when "10111000001111000" => rgb <= "000000";
					when "10111000001111001" => rgb <= "000000";
					when "10111000001111010" => rgb <= "000000";
					when "10111000001111011" => rgb <= "000000";
					when "10111000001111100" => rgb <= "000000";
					when "10111000001111101" => rgb <= "101010";
					when "10111000001111110" => rgb <= "111111";
					when "10111000001111111" => rgb <= "111111";
					when "10111000010000000" => rgb <= "111111";
					when "10111000010000001" => rgb <= "111111";
					when "10111000010000010" => rgb <= "111111";
					when "10111000010000011" => rgb <= "111111";
					when "10111000010000100" => rgb <= "111111";
					when "10111000010000101" => rgb <= "111111";
					when "10111000010000110" => rgb <= "111111";
					when "10111000010000111" => rgb <= "111111";
					when "10111000010001000" => rgb <= "111111";
					when "10111000010001001" => rgb <= "111111";
					when "10111000010001010" => rgb <= "111111";
					when "10111000010001011" => rgb <= "101010";
					when "10111000010001100" => rgb <= "000000";
					when "10111000010001101" => rgb <= "000000";
					when "10111000010001110" => rgb <= "000000";
					when "10111000010001111" => rgb <= "000000";
					when "10111000010010000" => rgb <= "000000";
					when "10111000010010001" => rgb <= "000000";
					when "10111000010010010" => rgb <= "000000";
					when "10111000010010011" => rgb <= "000000";
					when "10111000010010100" => rgb <= "000000";
					when "10111000010010101" => rgb <= "000000";
					when "10111000010010110" => rgb <= "000000";
					when "10111000010010111" => rgb <= "000000";
					when "10111000010011000" => rgb <= "000000";
					when "10111000010011001" => rgb <= "000000";
					when "10111000010011010" => rgb <= "000000";
					when "10111000010011011" => rgb <= "000000";
					when "10111000010011100" => rgb <= "000000";
					when "10111000010011101" => rgb <= "000000";
					when "10111000010011110" => rgb <= "000000";
					when "10111000010011111" => rgb <= "000000";
					when "10111000010100000" => rgb <= "000000";
					when "10111000010100001" => rgb <= "000000";
					when "10111000010100010" => rgb <= "010101";
					when "10111000010100011" => rgb <= "111111";
					when "10111000010100100" => rgb <= "101010";
					when "10111000010100101" => rgb <= "111111";
					when "10111000010100110" => rgb <= "111111";
					when "10111000010100111" => rgb <= "111111";
					when "10111000010101000" => rgb <= "111111";
					when "10111000010101001" => rgb <= "111111";
					when "10111000010101010" => rgb <= "000000";
					when "10111000010101011" => rgb <= "000000";
					when "10111000010101100" => rgb <= "000000";
					when "10111000010101101" => rgb <= "000000";
					when "10111000010101110" => rgb <= "000000";
					when "10111000010101111" => rgb <= "000000";
					when "10111000010110000" => rgb <= "000000";
					when "10111000010110001" => rgb <= "010101";
					when "10111000010110010" => rgb <= "111111";
					when "10111000010110011" => rgb <= "101010";
					when "10111000010110100" => rgb <= "111111";
					when "10111000010110101" => rgb <= "111111";
					when "10111000010110110" => rgb <= "101010";
					when "10111000010110111" => rgb <= "111111";
					when "10111000010111000" => rgb <= "101010";
					when "10111000010111001" => rgb <= "000000";
					when "10111000010111010" => rgb <= "000000";
					when "10111000010111011" => rgb <= "000000";
					when "10111000010111100" => rgb <= "000000";
					when "10111000010111101" => rgb <= "000000";
					when "10111000010111110" => rgb <= "000000";
					when "10111000010111111" => rgb <= "000000";
					when "10111000011000000" => rgb <= "010101";
					when "10111000011000001" => rgb <= "111111";
					when "10111000011000010" => rgb <= "101010";
					when "10111000011000011" => rgb <= "111111";
					when "10111000011000100" => rgb <= "101010";
					when "10111000011000101" => rgb <= "101010";
					when "10111000011000110" => rgb <= "111111";
					when "10111000011000111" => rgb <= "111111";
					when "10111000011001000" => rgb <= "111111";
					when "10111000011001001" => rgb <= "111111";
					when "10111000011001010" => rgb <= "111111";
					when "10111000011001011" => rgb <= "101010";
					when "10111000011001100" => rgb <= "111111";
					when "10111000011001101" => rgb <= "101010";
					when "10111000011001110" => rgb <= "111111";
					when "10111000011001111" => rgb <= "101010";
					when "10111000011010000" => rgb <= "000000";
					when "10111000011010001" => rgb <= "000000";
					when "10111000011010010" => rgb <= "000000";
					when "10111000011010011" => rgb <= "000000";
					when "10111000011010100" => rgb <= "000000";
					when "10111000011010101" => rgb <= "000000";
					when "10111000011010110" => rgb <= "000000";
					when "10111000011010111" => rgb <= "101010";
					when "10111000011011000" => rgb <= "101010";
					when "10111000011011001" => rgb <= "101010";
					when "10111000011011010" => rgb <= "101010";
					when "10111000011011011" => rgb <= "111111";
					when "10111000011011100" => rgb <= "111111";
					when "10111000011011101" => rgb <= "111111";
					when "10111000011011110" => rgb <= "111111";
					when "10111000011011111" => rgb <= "111111";
					when "10111000011100000" => rgb <= "111111";
					when "10111000011100001" => rgb <= "111111";
					when "10111000011100010" => rgb <= "111111";
					when "10111000011100011" => rgb <= "101010";
					when "10111000011100100" => rgb <= "111111";
					when "10111000011100101" => rgb <= "111111";
					when "10111000011100110" => rgb <= "000000";
					when "10111000011100111" => rgb <= "000000";
					when "10111000011101000" => rgb <= "000000";
					when "10111000011101001" => rgb <= "000000";
					when "10111000011101010" => rgb <= "000000";
					when "10111000011101011" => rgb <= "000000";
					when "10111000011101100" => rgb <= "000000";
					when "10111000011101101" => rgb <= "010101";
					when "10111000011101110" => rgb <= "111111";
					when "10111000011101111" => rgb <= "101010";
					when "10111000011110000" => rgb <= "111111";
					when "10111000011110001" => rgb <= "111111";
					when "10111000011110010" => rgb <= "111111";
					when "10111000011110011" => rgb <= "101010";
					when "10111000011110100" => rgb <= "101010";
					when "10111000011110101" => rgb <= "000000";
					when "10111000011110110" => rgb <= "000000";
					when "10111000011110111" => rgb <= "000000";
					when "10111000011111000" => rgb <= "000000";
					when "10111000011111001" => rgb <= "000000";
					when "10111000011111010" => rgb <= "000000";
					when "10111000011111011" => rgb <= "000000";
					when "10111000011111100" => rgb <= "000000";
					when "10111000011111101" => rgb <= "000000";
					when "10111000011111110" => rgb <= "000000";
					when "10111000011111111" => rgb <= "000000";
					when "10111000100000000" => rgb <= "000000";
					when "10111000100000001" => rgb <= "000000";
					when "10111000100000010" => rgb <= "000000";
					when "10111000100000011" => rgb <= "000000";
					when "10111000100000100" => rgb <= "101010";
					when "10111000100000101" => rgb <= "111111";
					when "10111000100000110" => rgb <= "101010";
					when "10111000100000111" => rgb <= "111111";
					when "10111000100001000" => rgb <= "111111";
					when "10111000100001001" => rgb <= "101010";
					when "10111000100001010" => rgb <= "111111";
					when "10111000100001011" => rgb <= "101010";
					when "10111000100001100" => rgb <= "101010";
					when "10111000100001101" => rgb <= "111111";
					when "10111000100001110" => rgb <= "111111";
					when "10111000100001111" => rgb <= "101010";
					when "10111000100010000" => rgb <= "111111";
					when "10111000100010001" => rgb <= "111111";
					when "10111000100010010" => rgb <= "111111";
					when "10111000100010011" => rgb <= "111111";
					when "10111000100010100" => rgb <= "111111";
					when "10111000100010101" => rgb <= "111111";
					when "10111000100010110" => rgb <= "111111";
					when "10111000100010111" => rgb <= "111111";
					when "10111000100011000" => rgb <= "101010";
					when "10111000100011001" => rgb <= "111111";
					when "10111000100011010" => rgb <= "101010";
					when "10111000100011011" => rgb <= "000000";
					when "10111000100011100" => rgb <= "000000";
					when "10111000100011101" => rgb <= "000000";
					when "10111000100011110" => rgb <= "000000";
					when "10111000100011111" => rgb <= "000000";
					when "10111000100100000" => rgb <= "000000";
					when "10111000100100001" => rgb <= "000000";
					when "10111000100100010" => rgb <= "101010";
					when "10111000100100011" => rgb <= "101010";
					when "10111000100100100" => rgb <= "101010";
					when "10111000100100101" => rgb <= "111111";
					when "10111000100100110" => rgb <= "111111";
					when "10111000100100111" => rgb <= "111111";
					when "10111000100101000" => rgb <= "111111";
					when "10111000100101001" => rgb <= "111111";
					when "10111000100101010" => rgb <= "111111";
					when "10111000100101011" => rgb <= "111111";
					when "10111000100101100" => rgb <= "111111";
					when "10111000100101101" => rgb <= "111111";
					when "10111000100101110" => rgb <= "101010";
					when "10111000100101111" => rgb <= "101010";
					when "10111000100110000" => rgb <= "111111";
					when "10111000100110001" => rgb <= "010101";
					when "10111000100110010" => rgb <= "000000";
					when "10111000100110011" => rgb <= "000000";
					when "10111000100110100" => rgb <= "000000";
					when "10111000100110101" => rgb <= "000000";
					when "10111000100110110" => rgb <= "000000";
					when "10111000100110111" => rgb <= "000000";
					when "10111000100111000" => rgb <= "000000";
					when "10111000100111001" => rgb <= "000000";
					when "10111000100111010" => rgb <= "000000";
					when "10111000100111011" => rgb <= "000000";
					when "10111000100111100" => rgb <= "000000";
					when "10111000100111101" => rgb <= "000000";
					when "10111000100111110" => rgb <= "000000";
					when "10111000100111111" => rgb <= "000000";
					when "10111001000000000" => rgb <= "000000";
					when "10111001000000001" => rgb <= "000000";
					when "10111001000000010" => rgb <= "000000";
					when "10111001000000011" => rgb <= "000000";
					when "10111001000000100" => rgb <= "000000";
					when "10111001000000101" => rgb <= "000000";
					when "10111001000000110" => rgb <= "000000";
					when "10111001000000111" => rgb <= "000000";
					when "10111001000001000" => rgb <= "000000";
					when "10111001000001001" => rgb <= "000000";
					when "10111001000001010" => rgb <= "000000";
					when "10111001000001011" => rgb <= "000000";
					when "10111001000001100" => rgb <= "010101";
					when "10111001000001101" => rgb <= "111111";
					when "10111001000001110" => rgb <= "101010";
					when "10111001000001111" => rgb <= "101010";
					when "10111001000010000" => rgb <= "101010";
					when "10111001000010001" => rgb <= "111111";
					when "10111001000010010" => rgb <= "101010";
					when "10111001000010011" => rgb <= "101010";
					when "10111001000010100" => rgb <= "101010";
					when "10111001000010101" => rgb <= "101010";
					when "10111001000010110" => rgb <= "101010";
					when "10111001000010111" => rgb <= "101010";
					when "10111001000011000" => rgb <= "101010";
					when "10111001000011001" => rgb <= "101010";
					when "10111001000011010" => rgb <= "101010";
					when "10111001000011011" => rgb <= "101010";
					when "10111001000011100" => rgb <= "101010";
					when "10111001000011101" => rgb <= "111111";
					when "10111001000011110" => rgb <= "111111";
					when "10111001000011111" => rgb <= "111111";
					when "10111001000100000" => rgb <= "101010";
					when "10111001000100001" => rgb <= "111111";
					when "10111001000100010" => rgb <= "101010";
					when "10111001000100011" => rgb <= "111111";
					when "10111001000100100" => rgb <= "101010";
					when "10111001000100101" => rgb <= "101010";
					when "10111001000100110" => rgb <= "111111";
					when "10111001000100111" => rgb <= "111111";
					when "10111001000101000" => rgb <= "101010";
					when "10111001000101001" => rgb <= "101010";
					when "10111001000101010" => rgb <= "101010";
					when "10111001000101011" => rgb <= "000000";
					when "10111001000101100" => rgb <= "000000";
					when "10111001000101101" => rgb <= "000000";
					when "10111001000101110" => rgb <= "000000";
					when "10111001000101111" => rgb <= "000000";
					when "10111001000110000" => rgb <= "000000";
					when "10111001000110001" => rgb <= "000000";
					when "10111001000110010" => rgb <= "000000";
					when "10111001000110011" => rgb <= "000000";
					when "10111001000110100" => rgb <= "000000";
					when "10111001000110101" => rgb <= "000000";
					when "10111001000110110" => rgb <= "000000";
					when "10111001000110111" => rgb <= "000000";
					when "10111001000111000" => rgb <= "000000";
					when "10111001000111001" => rgb <= "010101";
					when "10111001000111010" => rgb <= "111111";
					when "10111001000111011" => rgb <= "101010";
					when "10111001000111100" => rgb <= "111111";
					when "10111001000111101" => rgb <= "111111";
					when "10111001000111110" => rgb <= "111111";
					when "10111001000111111" => rgb <= "111111";
					when "10111001001000000" => rgb <= "101010";
					when "10111001001000001" => rgb <= "000000";
					when "10111001001000010" => rgb <= "000000";
					when "10111001001000011" => rgb <= "000000";
					when "10111001001000100" => rgb <= "000000";
					when "10111001001000101" => rgb <= "000000";
					when "10111001001000110" => rgb <= "000000";
					when "10111001001000111" => rgb <= "000000";
					when "10111001001001000" => rgb <= "000000";
					when "10111001001001001" => rgb <= "000000";
					when "10111001001001010" => rgb <= "000000";
					when "10111001001001011" => rgb <= "000000";
					when "10111001001001100" => rgb <= "000000";
					when "10111001001001101" => rgb <= "000000";
					when "10111001001001110" => rgb <= "000000";
					when "10111001001001111" => rgb <= "000000";
					when "10111001001010000" => rgb <= "101010";
					when "10111001001010001" => rgb <= "101010";
					when "10111001001010010" => rgb <= "101010";
					when "10111001001010011" => rgb <= "101010";
					when "10111001001010100" => rgb <= "111111";
					when "10111001001010101" => rgb <= "111111";
					when "10111001001010110" => rgb <= "101010";
					when "10111001001010111" => rgb <= "111111";
					when "10111001001011000" => rgb <= "111111";
					when "10111001001011001" => rgb <= "111111";
					when "10111001001011010" => rgb <= "111111";
					when "10111001001011011" => rgb <= "101010";
					when "10111001001011100" => rgb <= "111111";
					when "10111001001011101" => rgb <= "101010";
					when "10111001001011110" => rgb <= "101010";
					when "10111001001011111" => rgb <= "000000";
					when "10111001001100000" => rgb <= "000000";
					when "10111001001100001" => rgb <= "000000";
					when "10111001001100010" => rgb <= "000000";
					when "10111001001100011" => rgb <= "000000";
					when "10111001001100100" => rgb <= "000000";
					when "10111001001100101" => rgb <= "000000";
					when "10111001001100110" => rgb <= "010101";
					when "10111001001100111" => rgb <= "111111";
					when "10111001001101000" => rgb <= "101010";
					when "10111001001101001" => rgb <= "111111";
					when "10111001001101010" => rgb <= "101010";
					when "10111001001101011" => rgb <= "111111";
					when "10111001001101100" => rgb <= "101010";
					when "10111001001101101" => rgb <= "101010";
					when "10111001001101110" => rgb <= "000000";
					when "10111001001101111" => rgb <= "000000";
					when "10111001001110000" => rgb <= "000000";
					when "10111001001110001" => rgb <= "000000";
					when "10111001001110010" => rgb <= "000000";
					when "10111001001110011" => rgb <= "000000";
					when "10111001001110100" => rgb <= "000000";
					when "10111001001110101" => rgb <= "000000";
					when "10111001001110110" => rgb <= "000000";
					when "10111001001110111" => rgb <= "000000";
					when "10111001001111000" => rgb <= "000000";
					when "10111001001111001" => rgb <= "000000";
					when "10111001001111010" => rgb <= "000000";
					when "10111001001111011" => rgb <= "000000";
					when "10111001001111100" => rgb <= "000000";
					when "10111001001111101" => rgb <= "101010";
					when "10111001001111110" => rgb <= "111111";
					when "10111001001111111" => rgb <= "111111";
					when "10111001010000000" => rgb <= "111111";
					when "10111001010000001" => rgb <= "111111";
					when "10111001010000010" => rgb <= "111111";
					when "10111001010000011" => rgb <= "111111";
					when "10111001010000100" => rgb <= "111111";
					when "10111001010000101" => rgb <= "111111";
					when "10111001010000110" => rgb <= "111111";
					when "10111001010000111" => rgb <= "111111";
					when "10111001010001000" => rgb <= "111111";
					when "10111001010001001" => rgb <= "111111";
					when "10111001010001010" => rgb <= "111111";
					when "10111001010001011" => rgb <= "101010";
					when "10111001010001100" => rgb <= "000000";
					when "10111001010001101" => rgb <= "000000";
					when "10111001010001110" => rgb <= "000000";
					when "10111001010001111" => rgb <= "000000";
					when "10111001010010000" => rgb <= "000000";
					when "10111001010010001" => rgb <= "000000";
					when "10111001010010010" => rgb <= "000000";
					when "10111001010010011" => rgb <= "000000";
					when "10111001010010100" => rgb <= "000000";
					when "10111001010010101" => rgb <= "000000";
					when "10111001010010110" => rgb <= "000000";
					when "10111001010010111" => rgb <= "000000";
					when "10111001010011000" => rgb <= "000000";
					when "10111001010011001" => rgb <= "000000";
					when "10111001010011010" => rgb <= "000000";
					when "10111001010011011" => rgb <= "000000";
					when "10111001010011100" => rgb <= "000000";
					when "10111001010011101" => rgb <= "000000";
					when "10111001010011110" => rgb <= "000000";
					when "10111001010011111" => rgb <= "000000";
					when "10111001010100000" => rgb <= "000000";
					when "10111001010100001" => rgb <= "000000";
					when "10111001010100010" => rgb <= "010101";
					when "10111001010100011" => rgb <= "111111";
					when "10111001010100100" => rgb <= "101010";
					when "10111001010100101" => rgb <= "111111";
					when "10111001010100110" => rgb <= "111111";
					when "10111001010100111" => rgb <= "111111";
					when "10111001010101000" => rgb <= "111111";
					when "10111001010101001" => rgb <= "111111";
					when "10111001010101010" => rgb <= "000000";
					when "10111001010101011" => rgb <= "000000";
					when "10111001010101100" => rgb <= "000000";
					when "10111001010101101" => rgb <= "000000";
					when "10111001010101110" => rgb <= "000000";
					when "10111001010101111" => rgb <= "000000";
					when "10111001010110000" => rgb <= "000000";
					when "10111001010110001" => rgb <= "010101";
					when "10111001010110010" => rgb <= "101010";
					when "10111001010110011" => rgb <= "101010";
					when "10111001010110100" => rgb <= "101010";
					when "10111001010110101" => rgb <= "101010";
					when "10111001010110110" => rgb <= "101010";
					when "10111001010110111" => rgb <= "111111";
					when "10111001010111000" => rgb <= "101010";
					when "10111001010111001" => rgb <= "000000";
					when "10111001010111010" => rgb <= "000000";
					when "10111001010111011" => rgb <= "000000";
					when "10111001010111100" => rgb <= "000000";
					when "10111001010111101" => rgb <= "000000";
					when "10111001010111110" => rgb <= "000000";
					when "10111001010111111" => rgb <= "000000";
					when "10111001011000000" => rgb <= "010101";
					when "10111001011000001" => rgb <= "111111";
					when "10111001011000010" => rgb <= "101010";
					when "10111001011000011" => rgb <= "111111";
					when "10111001011000100" => rgb <= "101010";
					when "10111001011000101" => rgb <= "101010";
					when "10111001011000110" => rgb <= "111111";
					when "10111001011000111" => rgb <= "111111";
					when "10111001011001000" => rgb <= "111111";
					when "10111001011001001" => rgb <= "111111";
					when "10111001011001010" => rgb <= "111111";
					when "10111001011001011" => rgb <= "101010";
					when "10111001011001100" => rgb <= "111111";
					when "10111001011001101" => rgb <= "101010";
					when "10111001011001110" => rgb <= "111111";
					when "10111001011001111" => rgb <= "101010";
					when "10111001011010000" => rgb <= "000000";
					when "10111001011010001" => rgb <= "000000";
					when "10111001011010010" => rgb <= "000000";
					when "10111001011010011" => rgb <= "000000";
					when "10111001011010100" => rgb <= "000000";
					when "10111001011010101" => rgb <= "000000";
					when "10111001011010110" => rgb <= "000000";
					when "10111001011010111" => rgb <= "101010";
					when "10111001011011000" => rgb <= "101010";
					when "10111001011011001" => rgb <= "101010";
					when "10111001011011010" => rgb <= "101010";
					when "10111001011011011" => rgb <= "111111";
					when "10111001011011100" => rgb <= "111111";
					when "10111001011011101" => rgb <= "111111";
					when "10111001011011110" => rgb <= "111111";
					when "10111001011011111" => rgb <= "111111";
					when "10111001011100000" => rgb <= "111111";
					when "10111001011100001" => rgb <= "111111";
					when "10111001011100010" => rgb <= "111111";
					when "10111001011100011" => rgb <= "101010";
					when "10111001011100100" => rgb <= "111111";
					when "10111001011100101" => rgb <= "111111";
					when "10111001011100110" => rgb <= "000000";
					when "10111001011100111" => rgb <= "000000";
					when "10111001011101000" => rgb <= "000000";
					when "10111001011101001" => rgb <= "000000";
					when "10111001011101010" => rgb <= "000000";
					when "10111001011101011" => rgb <= "000000";
					when "10111001011101100" => rgb <= "000000";
					when "10111001011101101" => rgb <= "010101";
					when "10111001011101110" => rgb <= "111111";
					when "10111001011101111" => rgb <= "101010";
					when "10111001011110000" => rgb <= "111111";
					when "10111001011110001" => rgb <= "111111";
					when "10111001011110010" => rgb <= "111111";
					when "10111001011110011" => rgb <= "101010";
					when "10111001011110100" => rgb <= "101010";
					when "10111001011110101" => rgb <= "000000";
					when "10111001011110110" => rgb <= "000000";
					when "10111001011110111" => rgb <= "000000";
					when "10111001011111000" => rgb <= "000000";
					when "10111001011111001" => rgb <= "000000";
					when "10111001011111010" => rgb <= "000000";
					when "10111001011111011" => rgb <= "000000";
					when "10111001011111100" => rgb <= "000000";
					when "10111001011111101" => rgb <= "000000";
					when "10111001011111110" => rgb <= "000000";
					when "10111001011111111" => rgb <= "000000";
					when "10111001100000000" => rgb <= "000000";
					when "10111001100000001" => rgb <= "000000";
					when "10111001100000010" => rgb <= "000000";
					when "10111001100000011" => rgb <= "000000";
					when "10111001100000100" => rgb <= "101010";
					when "10111001100000101" => rgb <= "111111";
					when "10111001100000110" => rgb <= "101010";
					when "10111001100000111" => rgb <= "101010";
					when "10111001100001000" => rgb <= "101010";
					when "10111001100001001" => rgb <= "101010";
					when "10111001100001010" => rgb <= "101010";
					when "10111001100001011" => rgb <= "111111";
					when "10111001100001100" => rgb <= "111111";
					when "10111001100001101" => rgb <= "101010";
					when "10111001100001110" => rgb <= "101010";
					when "10111001100001111" => rgb <= "111111";
					when "10111001100010000" => rgb <= "111111";
					when "10111001100010001" => rgb <= "111111";
					when "10111001100010010" => rgb <= "111111";
					when "10111001100010011" => rgb <= "111111";
					when "10111001100010100" => rgb <= "111111";
					when "10111001100010101" => rgb <= "111111";
					when "10111001100010110" => rgb <= "111111";
					when "10111001100010111" => rgb <= "111111";
					when "10111001100011000" => rgb <= "101010";
					when "10111001100011001" => rgb <= "111111";
					when "10111001100011010" => rgb <= "101010";
					when "10111001100011011" => rgb <= "000000";
					when "10111001100011100" => rgb <= "000000";
					when "10111001100011101" => rgb <= "000000";
					when "10111001100011110" => rgb <= "000000";
					when "10111001100011111" => rgb <= "000000";
					when "10111001100100000" => rgb <= "000000";
					when "10111001100100001" => rgb <= "000000";
					when "10111001100100010" => rgb <= "101010";
					when "10111001100100011" => rgb <= "101010";
					when "10111001100100100" => rgb <= "101010";
					when "10111001100100101" => rgb <= "111111";
					when "10111001100100110" => rgb <= "111111";
					when "10111001100100111" => rgb <= "111111";
					when "10111001100101000" => rgb <= "111111";
					when "10111001100101001" => rgb <= "111111";
					when "10111001100101010" => rgb <= "111111";
					when "10111001100101011" => rgb <= "111111";
					when "10111001100101100" => rgb <= "111111";
					when "10111001100101101" => rgb <= "111111";
					when "10111001100101110" => rgb <= "101010";
					when "10111001100101111" => rgb <= "101010";
					when "10111001100110000" => rgb <= "111111";
					when "10111001100110001" => rgb <= "010101";
					when "10111001100110010" => rgb <= "000000";
					when "10111001100110011" => rgb <= "000000";
					when "10111001100110100" => rgb <= "000000";
					when "10111001100110101" => rgb <= "000000";
					when "10111001100110110" => rgb <= "000000";
					when "10111001100110111" => rgb <= "000000";
					when "10111001100111000" => rgb <= "000000";
					when "10111001100111001" => rgb <= "000000";
					when "10111001100111010" => rgb <= "000000";
					when "10111001100111011" => rgb <= "000000";
					when "10111001100111100" => rgb <= "000000";
					when "10111001100111101" => rgb <= "000000";
					when "10111001100111110" => rgb <= "000000";
					when "10111001100111111" => rgb <= "000000";
					when "10111010000000000" => rgb <= "000000";
					when "10111010000000001" => rgb <= "000000";
					when "10111010000000010" => rgb <= "000000";
					when "10111010000000011" => rgb <= "000000";
					when "10111010000000100" => rgb <= "000000";
					when "10111010000000101" => rgb <= "000000";
					when "10111010000000110" => rgb <= "000000";
					when "10111010000000111" => rgb <= "000000";
					when "10111010000001000" => rgb <= "000000";
					when "10111010000001001" => rgb <= "000000";
					when "10111010000001010" => rgb <= "000000";
					when "10111010000001011" => rgb <= "000000";
					when "10111010000001100" => rgb <= "010101";
					when "10111010000001101" => rgb <= "101010";
					when "10111010000001110" => rgb <= "101010";
					when "10111010000001111" => rgb <= "111111";
					when "10111010000010000" => rgb <= "111111";
					when "10111010000010001" => rgb <= "111111";
					when "10111010000010010" => rgb <= "101010";
					when "10111010000010011" => rgb <= "111111";
					when "10111010000010100" => rgb <= "101010";
					when "10111010000010101" => rgb <= "111111";
					when "10111010000010110" => rgb <= "111111";
					when "10111010000010111" => rgb <= "101010";
					when "10111010000011000" => rgb <= "101010";
					when "10111010000011001" => rgb <= "101010";
					when "10111010000011010" => rgb <= "101010";
					when "10111010000011011" => rgb <= "101010";
					when "10111010000011100" => rgb <= "101010";
					when "10111010000011101" => rgb <= "111111";
					when "10111010000011110" => rgb <= "111111";
					when "10111010000011111" => rgb <= "111111";
					when "10111010000100000" => rgb <= "111111";
					when "10111010000100001" => rgb <= "111111";
					when "10111010000100010" => rgb <= "101010";
					when "10111010000100011" => rgb <= "111111";
					when "10111010000100100" => rgb <= "101010";
					when "10111010000100101" => rgb <= "101010";
					when "10111010000100110" => rgb <= "111111";
					when "10111010000100111" => rgb <= "111111";
					when "10111010000101000" => rgb <= "101010";
					when "10111010000101001" => rgb <= "111111";
					when "10111010000101010" => rgb <= "101010";
					when "10111010000101011" => rgb <= "000000";
					when "10111010000101100" => rgb <= "000000";
					when "10111010000101101" => rgb <= "000000";
					when "10111010000101110" => rgb <= "000000";
					when "10111010000101111" => rgb <= "000000";
					when "10111010000110000" => rgb <= "000000";
					when "10111010000110001" => rgb <= "000000";
					when "10111010000110010" => rgb <= "000000";
					when "10111010000110011" => rgb <= "000000";
					when "10111010000110100" => rgb <= "000000";
					when "10111010000110101" => rgb <= "000000";
					when "10111010000110110" => rgb <= "000000";
					when "10111010000110111" => rgb <= "000000";
					when "10111010000111000" => rgb <= "000000";
					when "10111010000111001" => rgb <= "010101";
					when "10111010000111010" => rgb <= "111111";
					when "10111010000111011" => rgb <= "101010";
					when "10111010000111100" => rgb <= "111111";
					when "10111010000111101" => rgb <= "111111";
					when "10111010000111110" => rgb <= "111111";
					when "10111010000111111" => rgb <= "111111";
					when "10111010001000000" => rgb <= "101010";
					when "10111010001000001" => rgb <= "000000";
					when "10111010001000010" => rgb <= "000000";
					when "10111010001000011" => rgb <= "000000";
					when "10111010001000100" => rgb <= "000000";
					when "10111010001000101" => rgb <= "000000";
					when "10111010001000110" => rgb <= "000000";
					when "10111010001000111" => rgb <= "000000";
					when "10111010001001000" => rgb <= "000000";
					when "10111010001001001" => rgb <= "000000";
					when "10111010001001010" => rgb <= "000000";
					when "10111010001001011" => rgb <= "000000";
					when "10111010001001100" => rgb <= "000000";
					when "10111010001001101" => rgb <= "000000";
					when "10111010001001110" => rgb <= "000000";
					when "10111010001001111" => rgb <= "000000";
					when "10111010001010000" => rgb <= "101010";
					when "10111010001010001" => rgb <= "101010";
					when "10111010001010010" => rgb <= "101010";
					when "10111010001010011" => rgb <= "101010";
					when "10111010001010100" => rgb <= "111111";
					when "10111010001010101" => rgb <= "111111";
					when "10111010001010110" => rgb <= "101010";
					when "10111010001010111" => rgb <= "111111";
					when "10111010001011000" => rgb <= "111111";
					when "10111010001011001" => rgb <= "111111";
					when "10111010001011010" => rgb <= "111111";
					when "10111010001011011" => rgb <= "101010";
					when "10111010001011100" => rgb <= "111111";
					when "10111010001011101" => rgb <= "101010";
					when "10111010001011110" => rgb <= "101010";
					when "10111010001011111" => rgb <= "000000";
					when "10111010001100000" => rgb <= "000000";
					when "10111010001100001" => rgb <= "000000";
					when "10111010001100010" => rgb <= "000000";
					when "10111010001100011" => rgb <= "000000";
					when "10111010001100100" => rgb <= "000000";
					when "10111010001100101" => rgb <= "000000";
					when "10111010001100110" => rgb <= "010101";
					when "10111010001100111" => rgb <= "111111";
					when "10111010001101000" => rgb <= "101010";
					when "10111010001101001" => rgb <= "111111";
					when "10111010001101010" => rgb <= "101010";
					when "10111010001101011" => rgb <= "111111";
					when "10111010001101100" => rgb <= "101010";
					when "10111010001101101" => rgb <= "101010";
					when "10111010001101110" => rgb <= "000000";
					when "10111010001101111" => rgb <= "000000";
					when "10111010001110000" => rgb <= "000000";
					when "10111010001110001" => rgb <= "000000";
					when "10111010001110010" => rgb <= "000000";
					when "10111010001110011" => rgb <= "000000";
					when "10111010001110100" => rgb <= "000000";
					when "10111010001110101" => rgb <= "000000";
					when "10111010001110110" => rgb <= "000000";
					when "10111010001110111" => rgb <= "000000";
					when "10111010001111000" => rgb <= "000000";
					when "10111010001111001" => rgb <= "000000";
					when "10111010001111010" => rgb <= "000000";
					when "10111010001111011" => rgb <= "000000";
					when "10111010001111100" => rgb <= "000000";
					when "10111010001111101" => rgb <= "101010";
					when "10111010001111110" => rgb <= "111111";
					when "10111010001111111" => rgb <= "111111";
					when "10111010010000000" => rgb <= "111111";
					when "10111010010000001" => rgb <= "111111";
					when "10111010010000010" => rgb <= "111111";
					when "10111010010000011" => rgb <= "111111";
					when "10111010010000100" => rgb <= "111111";
					when "10111010010000101" => rgb <= "111111";
					when "10111010010000110" => rgb <= "111111";
					when "10111010010000111" => rgb <= "111111";
					when "10111010010001000" => rgb <= "111111";
					when "10111010010001001" => rgb <= "111111";
					when "10111010010001010" => rgb <= "111111";
					when "10111010010001011" => rgb <= "101010";
					when "10111010010001100" => rgb <= "000000";
					when "10111010010001101" => rgb <= "000000";
					when "10111010010001110" => rgb <= "000000";
					when "10111010010001111" => rgb <= "000000";
					when "10111010010010000" => rgb <= "000000";
					when "10111010010010001" => rgb <= "000000";
					when "10111010010010010" => rgb <= "000000";
					when "10111010010010011" => rgb <= "000000";
					when "10111010010010100" => rgb <= "000000";
					when "10111010010010101" => rgb <= "000000";
					when "10111010010010110" => rgb <= "000000";
					when "10111010010010111" => rgb <= "000000";
					when "10111010010011000" => rgb <= "000000";
					when "10111010010011001" => rgb <= "000000";
					when "10111010010011010" => rgb <= "000000";
					when "10111010010011011" => rgb <= "000000";
					when "10111010010011100" => rgb <= "000000";
					when "10111010010011101" => rgb <= "000000";
					when "10111010010011110" => rgb <= "000000";
					when "10111010010011111" => rgb <= "000000";
					when "10111010010100000" => rgb <= "000000";
					when "10111010010100001" => rgb <= "000000";
					when "10111010010100010" => rgb <= "010101";
					when "10111010010100011" => rgb <= "111111";
					when "10111010010100100" => rgb <= "101010";
					when "10111010010100101" => rgb <= "111111";
					when "10111010010100110" => rgb <= "111111";
					when "10111010010100111" => rgb <= "111111";
					when "10111010010101000" => rgb <= "111111";
					when "10111010010101001" => rgb <= "111111";
					when "10111010010101010" => rgb <= "000000";
					when "10111010010101011" => rgb <= "000000";
					when "10111010010101100" => rgb <= "000000";
					when "10111010010101101" => rgb <= "000000";
					when "10111010010101110" => rgb <= "000000";
					when "10111010010101111" => rgb <= "000000";
					when "10111010010110000" => rgb <= "000000";
					when "10111010010110001" => rgb <= "010101";
					when "10111010010110010" => rgb <= "101010";
					when "10111010010110011" => rgb <= "101010";
					when "10111010010110100" => rgb <= "101010";
					when "10111010010110101" => rgb <= "101010";
					when "10111010010110110" => rgb <= "101010";
					when "10111010010110111" => rgb <= "111111";
					when "10111010010111000" => rgb <= "101010";
					when "10111010010111001" => rgb <= "000000";
					when "10111010010111010" => rgb <= "000000";
					when "10111010010111011" => rgb <= "000000";
					when "10111010010111100" => rgb <= "000000";
					when "10111010010111101" => rgb <= "000000";
					when "10111010010111110" => rgb <= "000000";
					when "10111010010111111" => rgb <= "000000";
					when "10111010011000000" => rgb <= "010101";
					when "10111010011000001" => rgb <= "101010";
					when "10111010011000010" => rgb <= "101010";
					when "10111010011000011" => rgb <= "111111";
					when "10111010011000100" => rgb <= "101010";
					when "10111010011000101" => rgb <= "101010";
					when "10111010011000110" => rgb <= "111111";
					when "10111010011000111" => rgb <= "111111";
					when "10111010011001000" => rgb <= "111111";
					when "10111010011001001" => rgb <= "111111";
					when "10111010011001010" => rgb <= "111111";
					when "10111010011001011" => rgb <= "101010";
					when "10111010011001100" => rgb <= "111111";
					when "10111010011001101" => rgb <= "101010";
					when "10111010011001110" => rgb <= "111111";
					when "10111010011001111" => rgb <= "101010";
					when "10111010011010000" => rgb <= "000000";
					when "10111010011010001" => rgb <= "000000";
					when "10111010011010010" => rgb <= "000000";
					when "10111010011010011" => rgb <= "000000";
					when "10111010011010100" => rgb <= "000000";
					when "10111010011010101" => rgb <= "000000";
					when "10111010011010110" => rgb <= "000000";
					when "10111010011010111" => rgb <= "101010";
					when "10111010011011000" => rgb <= "101010";
					when "10111010011011001" => rgb <= "101010";
					when "10111010011011010" => rgb <= "101010";
					when "10111010011011011" => rgb <= "111111";
					when "10111010011011100" => rgb <= "111111";
					when "10111010011011101" => rgb <= "111111";
					when "10111010011011110" => rgb <= "111111";
					when "10111010011011111" => rgb <= "111111";
					when "10111010011100000" => rgb <= "111111";
					when "10111010011100001" => rgb <= "111111";
					when "10111010011100010" => rgb <= "111111";
					when "10111010011100011" => rgb <= "101010";
					when "10111010011100100" => rgb <= "111111";
					when "10111010011100101" => rgb <= "111111";
					when "10111010011100110" => rgb <= "000000";
					when "10111010011100111" => rgb <= "000000";
					when "10111010011101000" => rgb <= "000000";
					when "10111010011101001" => rgb <= "000000";
					when "10111010011101010" => rgb <= "000000";
					when "10111010011101011" => rgb <= "000000";
					when "10111010011101100" => rgb <= "000000";
					when "10111010011101101" => rgb <= "010101";
					when "10111010011101110" => rgb <= "111111";
					when "10111010011101111" => rgb <= "101010";
					when "10111010011110000" => rgb <= "111111";
					when "10111010011110001" => rgb <= "111111";
					when "10111010011110010" => rgb <= "111111";
					when "10111010011110011" => rgb <= "101010";
					when "10111010011110100" => rgb <= "101010";
					when "10111010011110101" => rgb <= "000000";
					when "10111010011110110" => rgb <= "000000";
					when "10111010011110111" => rgb <= "000000";
					when "10111010011111000" => rgb <= "000000";
					when "10111010011111001" => rgb <= "000000";
					when "10111010011111010" => rgb <= "000000";
					when "10111010011111011" => rgb <= "000000";
					when "10111010011111100" => rgb <= "000000";
					when "10111010011111101" => rgb <= "000000";
					when "10111010011111110" => rgb <= "000000";
					when "10111010011111111" => rgb <= "000000";
					when "10111010100000000" => rgb <= "000000";
					when "10111010100000001" => rgb <= "000000";
					when "10111010100000010" => rgb <= "000000";
					when "10111010100000011" => rgb <= "000000";
					when "10111010100000100" => rgb <= "101010";
					when "10111010100000101" => rgb <= "111111";
					when "10111010100000110" => rgb <= "101010";
					when "10111010100000111" => rgb <= "111111";
					when "10111010100001000" => rgb <= "101010";
					when "10111010100001001" => rgb <= "111111";
					when "10111010100001010" => rgb <= "101010";
					when "10111010100001011" => rgb <= "101010";
					when "10111010100001100" => rgb <= "111111";
					when "10111010100001101" => rgb <= "111111";
					when "10111010100001110" => rgb <= "101010";
					when "10111010100001111" => rgb <= "101010";
					when "10111010100010000" => rgb <= "111111";
					when "10111010100010001" => rgb <= "111111";
					when "10111010100010010" => rgb <= "111111";
					when "10111010100010011" => rgb <= "111111";
					when "10111010100010100" => rgb <= "111111";
					when "10111010100010101" => rgb <= "111111";
					when "10111010100010110" => rgb <= "111111";
					when "10111010100010111" => rgb <= "111111";
					when "10111010100011000" => rgb <= "101010";
					when "10111010100011001" => rgb <= "111111";
					when "10111010100011010" => rgb <= "101010";
					when "10111010100011011" => rgb <= "000000";
					when "10111010100011100" => rgb <= "000000";
					when "10111010100011101" => rgb <= "000000";
					when "10111010100011110" => rgb <= "000000";
					when "10111010100011111" => rgb <= "000000";
					when "10111010100100000" => rgb <= "000000";
					when "10111010100100001" => rgb <= "000000";
					when "10111010100100010" => rgb <= "101010";
					when "10111010100100011" => rgb <= "101010";
					when "10111010100100100" => rgb <= "101010";
					when "10111010100100101" => rgb <= "111111";
					when "10111010100100110" => rgb <= "111111";
					when "10111010100100111" => rgb <= "111111";
					when "10111010100101000" => rgb <= "111111";
					when "10111010100101001" => rgb <= "111111";
					when "10111010100101010" => rgb <= "111111";
					when "10111010100101011" => rgb <= "111111";
					when "10111010100101100" => rgb <= "111111";
					when "10111010100101101" => rgb <= "111111";
					when "10111010100101110" => rgb <= "101010";
					when "10111010100101111" => rgb <= "101010";
					when "10111010100110000" => rgb <= "111111";
					when "10111010100110001" => rgb <= "010101";
					when "10111010100110010" => rgb <= "000000";
					when "10111010100110011" => rgb <= "000000";
					when "10111010100110100" => rgb <= "000000";
					when "10111010100110101" => rgb <= "000000";
					when "10111010100110110" => rgb <= "000000";
					when "10111010100110111" => rgb <= "000000";
					when "10111010100111000" => rgb <= "000000";
					when "10111010100111001" => rgb <= "000000";
					when "10111010100111010" => rgb <= "000000";
					when "10111010100111011" => rgb <= "000000";
					when "10111010100111100" => rgb <= "000000";
					when "10111010100111101" => rgb <= "000000";
					when "10111010100111110" => rgb <= "000000";
					when "10111010100111111" => rgb <= "000000";
					when "10111011000000000" => rgb <= "000000";
					when "10111011000000001" => rgb <= "000000";
					when "10111011000000010" => rgb <= "000000";
					when "10111011000000011" => rgb <= "000000";
					when "10111011000000100" => rgb <= "000000";
					when "10111011000000101" => rgb <= "000000";
					when "10111011000000110" => rgb <= "000000";
					when "10111011000000111" => rgb <= "000000";
					when "10111011000001000" => rgb <= "000000";
					when "10111011000001001" => rgb <= "000000";
					when "10111011000001010" => rgb <= "000000";
					when "10111011000001011" => rgb <= "000000";
					when "10111011000001100" => rgb <= "010101";
					when "10111011000001101" => rgb <= "111111";
					when "10111011000001110" => rgb <= "111111";
					when "10111011000001111" => rgb <= "101010";
					when "10111011000010000" => rgb <= "101010";
					when "10111011000010001" => rgb <= "101010";
					when "10111011000010010" => rgb <= "111111";
					when "10111011000010011" => rgb <= "101010";
					when "10111011000010100" => rgb <= "111111";
					when "10111011000010101" => rgb <= "101010";
					when "10111011000010110" => rgb <= "111111";
					when "10111011000010111" => rgb <= "111111";
					when "10111011000011000" => rgb <= "111111";
					when "10111011000011001" => rgb <= "111111";
					when "10111011000011010" => rgb <= "111111";
					when "10111011000011011" => rgb <= "111111";
					when "10111011000011100" => rgb <= "111111";
					when "10111011000011101" => rgb <= "111111";
					when "10111011000011110" => rgb <= "111111";
					when "10111011000011111" => rgb <= "111111";
					when "10111011000100000" => rgb <= "111111";
					when "10111011000100001" => rgb <= "101010";
					when "10111011000100010" => rgb <= "111111";
					when "10111011000100011" => rgb <= "101010";
					when "10111011000100100" => rgb <= "111111";
					when "10111011000100101" => rgb <= "111111";
					when "10111011000100110" => rgb <= "101010";
					when "10111011000100111" => rgb <= "101010";
					when "10111011000101000" => rgb <= "101010";
					when "10111011000101001" => rgb <= "111111";
					when "10111011000101010" => rgb <= "101010";
					when "10111011000101011" => rgb <= "000000";
					when "10111011000101100" => rgb <= "000000";
					when "10111011000101101" => rgb <= "000000";
					when "10111011000101110" => rgb <= "000000";
					when "10111011000101111" => rgb <= "000000";
					when "10111011000110000" => rgb <= "000000";
					when "10111011000110001" => rgb <= "000000";
					when "10111011000110010" => rgb <= "000000";
					when "10111011000110011" => rgb <= "000000";
					when "10111011000110100" => rgb <= "000000";
					when "10111011000110101" => rgb <= "000000";
					when "10111011000110110" => rgb <= "000000";
					when "10111011000110111" => rgb <= "000000";
					when "10111011000111000" => rgb <= "000000";
					when "10111011000111001" => rgb <= "010101";
					when "10111011000111010" => rgb <= "111111";
					when "10111011000111011" => rgb <= "101010";
					when "10111011000111100" => rgb <= "111111";
					when "10111011000111101" => rgb <= "111111";
					when "10111011000111110" => rgb <= "111111";
					when "10111011000111111" => rgb <= "111111";
					when "10111011001000000" => rgb <= "101010";
					when "10111011001000001" => rgb <= "000000";
					when "10111011001000010" => rgb <= "000000";
					when "10111011001000011" => rgb <= "000000";
					when "10111011001000100" => rgb <= "000000";
					when "10111011001000101" => rgb <= "000000";
					when "10111011001000110" => rgb <= "000000";
					when "10111011001000111" => rgb <= "000000";
					when "10111011001001000" => rgb <= "000000";
					when "10111011001001001" => rgb <= "000000";
					when "10111011001001010" => rgb <= "000000";
					when "10111011001001011" => rgb <= "000000";
					when "10111011001001100" => rgb <= "000000";
					when "10111011001001101" => rgb <= "000000";
					when "10111011001001110" => rgb <= "000000";
					when "10111011001001111" => rgb <= "000000";
					when "10111011001010000" => rgb <= "101010";
					when "10111011001010001" => rgb <= "101010";
					when "10111011001010010" => rgb <= "101010";
					when "10111011001010011" => rgb <= "101010";
					when "10111011001010100" => rgb <= "111111";
					when "10111011001010101" => rgb <= "111111";
					when "10111011001010110" => rgb <= "101010";
					when "10111011001010111" => rgb <= "111111";
					when "10111011001011000" => rgb <= "111111";
					when "10111011001011001" => rgb <= "111111";
					when "10111011001011010" => rgb <= "111111";
					when "10111011001011011" => rgb <= "101010";
					when "10111011001011100" => rgb <= "111111";
					when "10111011001011101" => rgb <= "101010";
					when "10111011001011110" => rgb <= "101010";
					when "10111011001011111" => rgb <= "000000";
					when "10111011001100000" => rgb <= "000000";
					when "10111011001100001" => rgb <= "000000";
					when "10111011001100010" => rgb <= "000000";
					when "10111011001100011" => rgb <= "000000";
					when "10111011001100100" => rgb <= "000000";
					when "10111011001100101" => rgb <= "000000";
					when "10111011001100110" => rgb <= "010101";
					when "10111011001100111" => rgb <= "111111";
					when "10111011001101000" => rgb <= "101010";
					when "10111011001101001" => rgb <= "111111";
					when "10111011001101010" => rgb <= "101010";
					when "10111011001101011" => rgb <= "111111";
					when "10111011001101100" => rgb <= "101010";
					when "10111011001101101" => rgb <= "101010";
					when "10111011001101110" => rgb <= "000000";
					when "10111011001101111" => rgb <= "000000";
					when "10111011001110000" => rgb <= "000000";
					when "10111011001110001" => rgb <= "000000";
					when "10111011001110010" => rgb <= "000000";
					when "10111011001110011" => rgb <= "000000";
					when "10111011001110100" => rgb <= "000000";
					when "10111011001110101" => rgb <= "000000";
					when "10111011001110110" => rgb <= "000000";
					when "10111011001110111" => rgb <= "000000";
					when "10111011001111000" => rgb <= "000000";
					when "10111011001111001" => rgb <= "000000";
					when "10111011001111010" => rgb <= "000000";
					when "10111011001111011" => rgb <= "000000";
					when "10111011001111100" => rgb <= "000000";
					when "10111011001111101" => rgb <= "101010";
					when "10111011001111110" => rgb <= "111111";
					when "10111011001111111" => rgb <= "111111";
					when "10111011010000000" => rgb <= "111111";
					when "10111011010000001" => rgb <= "111111";
					when "10111011010000010" => rgb <= "111111";
					when "10111011010000011" => rgb <= "111111";
					when "10111011010000100" => rgb <= "111111";
					when "10111011010000101" => rgb <= "111111";
					when "10111011010000110" => rgb <= "111111";
					when "10111011010000111" => rgb <= "111111";
					when "10111011010001000" => rgb <= "111111";
					when "10111011010001001" => rgb <= "111111";
					when "10111011010001010" => rgb <= "111111";
					when "10111011010001011" => rgb <= "101010";
					when "10111011010001100" => rgb <= "000000";
					when "10111011010001101" => rgb <= "000000";
					when "10111011010001110" => rgb <= "000000";
					when "10111011010001111" => rgb <= "000000";
					when "10111011010010000" => rgb <= "000000";
					when "10111011010010001" => rgb <= "000000";
					when "10111011010010010" => rgb <= "000000";
					when "10111011010010011" => rgb <= "000000";
					when "10111011010010100" => rgb <= "000000";
					when "10111011010010101" => rgb <= "000000";
					when "10111011010010110" => rgb <= "000000";
					when "10111011010010111" => rgb <= "000000";
					when "10111011010011000" => rgb <= "000000";
					when "10111011010011001" => rgb <= "000000";
					when "10111011010011010" => rgb <= "000000";
					when "10111011010011011" => rgb <= "000000";
					when "10111011010011100" => rgb <= "000000";
					when "10111011010011101" => rgb <= "000000";
					when "10111011010011110" => rgb <= "000000";
					when "10111011010011111" => rgb <= "000000";
					when "10111011010100000" => rgb <= "000000";
					when "10111011010100001" => rgb <= "000000";
					when "10111011010100010" => rgb <= "010101";
					when "10111011010100011" => rgb <= "111111";
					when "10111011010100100" => rgb <= "101010";
					when "10111011010100101" => rgb <= "111111";
					when "10111011010100110" => rgb <= "111111";
					when "10111011010100111" => rgb <= "111111";
					when "10111011010101000" => rgb <= "111111";
					when "10111011010101001" => rgb <= "111111";
					when "10111011010101010" => rgb <= "000000";
					when "10111011010101011" => rgb <= "000000";
					when "10111011010101100" => rgb <= "000000";
					when "10111011010101101" => rgb <= "000000";
					when "10111011010101110" => rgb <= "000000";
					when "10111011010101111" => rgb <= "000000";
					when "10111011010110000" => rgb <= "000000";
					when "10111011010110001" => rgb <= "010101";
					when "10111011010110010" => rgb <= "101010";
					when "10111011010110011" => rgb <= "101010";
					when "10111011010110100" => rgb <= "111111";
					when "10111011010110101" => rgb <= "111111";
					when "10111011010110110" => rgb <= "101010";
					when "10111011010110111" => rgb <= "111111";
					when "10111011010111000" => rgb <= "101010";
					when "10111011010111001" => rgb <= "000000";
					when "10111011010111010" => rgb <= "000000";
					when "10111011010111011" => rgb <= "000000";
					when "10111011010111100" => rgb <= "000000";
					when "10111011010111101" => rgb <= "000000";
					when "10111011010111110" => rgb <= "000000";
					when "10111011010111111" => rgb <= "000000";
					when "10111011011000000" => rgb <= "010101";
					when "10111011011000001" => rgb <= "101010";
					when "10111011011000010" => rgb <= "101010";
					when "10111011011000011" => rgb <= "111111";
					when "10111011011000100" => rgb <= "111111";
					when "10111011011000101" => rgb <= "101010";
					when "10111011011000110" => rgb <= "111111";
					when "10111011011000111" => rgb <= "101010";
					when "10111011011001000" => rgb <= "111111";
					when "10111011011001001" => rgb <= "111111";
					when "10111011011001010" => rgb <= "111111";
					when "10111011011001011" => rgb <= "101010";
					when "10111011011001100" => rgb <= "111111";
					when "10111011011001101" => rgb <= "101010";
					when "10111011011001110" => rgb <= "111111";
					when "10111011011001111" => rgb <= "101010";
					when "10111011011010000" => rgb <= "000000";
					when "10111011011010001" => rgb <= "000000";
					when "10111011011010010" => rgb <= "000000";
					when "10111011011010011" => rgb <= "000000";
					when "10111011011010100" => rgb <= "000000";
					when "10111011011010101" => rgb <= "000000";
					when "10111011011010110" => rgb <= "000000";
					when "10111011011010111" => rgb <= "101010";
					when "10111011011011000" => rgb <= "101010";
					when "10111011011011001" => rgb <= "101010";
					when "10111011011011010" => rgb <= "101010";
					when "10111011011011011" => rgb <= "111111";
					when "10111011011011100" => rgb <= "111111";
					when "10111011011011101" => rgb <= "111111";
					when "10111011011011110" => rgb <= "111111";
					when "10111011011011111" => rgb <= "111111";
					when "10111011011100000" => rgb <= "111111";
					when "10111011011100001" => rgb <= "111111";
					when "10111011011100010" => rgb <= "111111";
					when "10111011011100011" => rgb <= "101010";
					when "10111011011100100" => rgb <= "111111";
					when "10111011011100101" => rgb <= "111111";
					when "10111011011100110" => rgb <= "000000";
					when "10111011011100111" => rgb <= "000000";
					when "10111011011101000" => rgb <= "000000";
					when "10111011011101001" => rgb <= "000000";
					when "10111011011101010" => rgb <= "000000";
					when "10111011011101011" => rgb <= "000000";
					when "10111011011101100" => rgb <= "000000";
					when "10111011011101101" => rgb <= "010101";
					when "10111011011101110" => rgb <= "111111";
					when "10111011011101111" => rgb <= "101010";
					when "10111011011110000" => rgb <= "111111";
					when "10111011011110001" => rgb <= "111111";
					when "10111011011110010" => rgb <= "111111";
					when "10111011011110011" => rgb <= "101010";
					when "10111011011110100" => rgb <= "101010";
					when "10111011011110101" => rgb <= "000000";
					when "10111011011110110" => rgb <= "000000";
					when "10111011011110111" => rgb <= "000000";
					when "10111011011111000" => rgb <= "000000";
					when "10111011011111001" => rgb <= "000000";
					when "10111011011111010" => rgb <= "000000";
					when "10111011011111011" => rgb <= "000000";
					when "10111011011111100" => rgb <= "000000";
					when "10111011011111101" => rgb <= "000000";
					when "10111011011111110" => rgb <= "000000";
					when "10111011011111111" => rgb <= "000000";
					when "10111011100000000" => rgb <= "000000";
					when "10111011100000001" => rgb <= "000000";
					when "10111011100000010" => rgb <= "000000";
					when "10111011100000011" => rgb <= "000000";
					when "10111011100000100" => rgb <= "101010";
					when "10111011100000101" => rgb <= "111111";
					when "10111011100000110" => rgb <= "101010";
					when "10111011100000111" => rgb <= "101010";
					when "10111011100001000" => rgb <= "101010";
					when "10111011100001001" => rgb <= "111111";
					when "10111011100001010" => rgb <= "111111";
					when "10111011100001011" => rgb <= "111111";
					when "10111011100001100" => rgb <= "111111";
					when "10111011100001101" => rgb <= "111111";
					when "10111011100001110" => rgb <= "101010";
					when "10111011100001111" => rgb <= "111111";
					when "10111011100010000" => rgb <= "111111";
					when "10111011100010001" => rgb <= "111111";
					when "10111011100010010" => rgb <= "111111";
					when "10111011100010011" => rgb <= "111111";
					when "10111011100010100" => rgb <= "111111";
					when "10111011100010101" => rgb <= "111111";
					when "10111011100010110" => rgb <= "111111";
					when "10111011100010111" => rgb <= "111111";
					when "10111011100011000" => rgb <= "101010";
					when "10111011100011001" => rgb <= "111111";
					when "10111011100011010" => rgb <= "101010";
					when "10111011100011011" => rgb <= "000000";
					when "10111011100011100" => rgb <= "000000";
					when "10111011100011101" => rgb <= "000000";
					when "10111011100011110" => rgb <= "000000";
					when "10111011100011111" => rgb <= "000000";
					when "10111011100100000" => rgb <= "000000";
					when "10111011100100001" => rgb <= "000000";
					when "10111011100100010" => rgb <= "101010";
					when "10111011100100011" => rgb <= "101010";
					when "10111011100100100" => rgb <= "101010";
					when "10111011100100101" => rgb <= "111111";
					when "10111011100100110" => rgb <= "111111";
					when "10111011100100111" => rgb <= "111111";
					when "10111011100101000" => rgb <= "111111";
					when "10111011100101001" => rgb <= "111111";
					when "10111011100101010" => rgb <= "111111";
					when "10111011100101011" => rgb <= "111111";
					when "10111011100101100" => rgb <= "111111";
					when "10111011100101101" => rgb <= "111111";
					when "10111011100101110" => rgb <= "101010";
					when "10111011100101111" => rgb <= "101010";
					when "10111011100110000" => rgb <= "111111";
					when "10111011100110001" => rgb <= "010101";
					when "10111011100110010" => rgb <= "000000";
					when "10111011100110011" => rgb <= "000000";
					when "10111011100110100" => rgb <= "000000";
					when "10111011100110101" => rgb <= "000000";
					when "10111011100110110" => rgb <= "000000";
					when "10111011100110111" => rgb <= "000000";
					when "10111011100111000" => rgb <= "000000";
					when "10111011100111001" => rgb <= "000000";
					when "10111011100111010" => rgb <= "000000";
					when "10111011100111011" => rgb <= "000000";
					when "10111011100111100" => rgb <= "000000";
					when "10111011100111101" => rgb <= "000000";
					when "10111011100111110" => rgb <= "000000";
					when "10111011100111111" => rgb <= "000000";
					when "10111100000000000" => rgb <= "000000";
					when "10111100000000001" => rgb <= "000000";
					when "10111100000000010" => rgb <= "000000";
					when "10111100000000011" => rgb <= "000000";
					when "10111100000000100" => rgb <= "000000";
					when "10111100000000101" => rgb <= "000000";
					when "10111100000000110" => rgb <= "000000";
					when "10111100000000111" => rgb <= "000000";
					when "10111100000001000" => rgb <= "000000";
					when "10111100000001001" => rgb <= "000000";
					when "10111100000001010" => rgb <= "000000";
					when "10111100000001011" => rgb <= "000000";
					when "10111100000001100" => rgb <= "010101";
					when "10111100000001101" => rgb <= "101010";
					when "10111100000001110" => rgb <= "101010";
					when "10111100000001111" => rgb <= "101010";
					when "10111100000010000" => rgb <= "101010";
					when "10111100000010001" => rgb <= "111111";
					when "10111100000010010" => rgb <= "101010";
					when "10111100000010011" => rgb <= "101010";
					when "10111100000010100" => rgb <= "111111";
					when "10111100000010101" => rgb <= "111111";
					when "10111100000010110" => rgb <= "101010";
					when "10111100000010111" => rgb <= "111111";
					when "10111100000011000" => rgb <= "111111";
					when "10111100000011001" => rgb <= "111111";
					when "10111100000011010" => rgb <= "111111";
					when "10111100000011011" => rgb <= "111111";
					when "10111100000011100" => rgb <= "111111";
					when "10111100000011101" => rgb <= "111111";
					when "10111100000011110" => rgb <= "111111";
					when "10111100000011111" => rgb <= "111111";
					when "10111100000100000" => rgb <= "111111";
					when "10111100000100001" => rgb <= "101010";
					when "10111100000100010" => rgb <= "111111";
					when "10111100000100011" => rgb <= "101010";
					when "10111100000100100" => rgb <= "101010";
					when "10111100000100101" => rgb <= "111111";
					when "10111100000100110" => rgb <= "111111";
					when "10111100000100111" => rgb <= "111111";
					when "10111100000101000" => rgb <= "111111";
					when "10111100000101001" => rgb <= "101010";
					when "10111100000101010" => rgb <= "101010";
					when "10111100000101011" => rgb <= "000000";
					when "10111100000101100" => rgb <= "000000";
					when "10111100000101101" => rgb <= "000000";
					when "10111100000101110" => rgb <= "000000";
					when "10111100000101111" => rgb <= "000000";
					when "10111100000110000" => rgb <= "000000";
					when "10111100000110001" => rgb <= "000000";
					when "10111100000110010" => rgb <= "000000";
					when "10111100000110011" => rgb <= "000000";
					when "10111100000110100" => rgb <= "000000";
					when "10111100000110101" => rgb <= "000000";
					when "10111100000110110" => rgb <= "000000";
					when "10111100000110111" => rgb <= "000000";
					when "10111100000111000" => rgb <= "000000";
					when "10111100000111001" => rgb <= "010101";
					when "10111100000111010" => rgb <= "111111";
					when "10111100000111011" => rgb <= "101010";
					when "10111100000111100" => rgb <= "101010";
					when "10111100000111101" => rgb <= "111111";
					when "10111100000111110" => rgb <= "111111";
					when "10111100000111111" => rgb <= "111111";
					when "10111100001000000" => rgb <= "101010";
					when "10111100001000001" => rgb <= "000000";
					when "10111100001000010" => rgb <= "000000";
					when "10111100001000011" => rgb <= "000000";
					when "10111100001000100" => rgb <= "000000";
					when "10111100001000101" => rgb <= "000000";
					when "10111100001000110" => rgb <= "000000";
					when "10111100001000111" => rgb <= "000000";
					when "10111100001001000" => rgb <= "000000";
					when "10111100001001001" => rgb <= "000000";
					when "10111100001001010" => rgb <= "000000";
					when "10111100001001011" => rgb <= "000000";
					when "10111100001001100" => rgb <= "000000";
					when "10111100001001101" => rgb <= "000000";
					when "10111100001001110" => rgb <= "000000";
					when "10111100001001111" => rgb <= "000000";
					when "10111100001010000" => rgb <= "101010";
					when "10111100001010001" => rgb <= "101010";
					when "10111100001010010" => rgb <= "101010";
					when "10111100001010011" => rgb <= "101010";
					when "10111100001010100" => rgb <= "111111";
					when "10111100001010101" => rgb <= "111111";
					when "10111100001010110" => rgb <= "101010";
					when "10111100001010111" => rgb <= "111111";
					when "10111100001011000" => rgb <= "111111";
					when "10111100001011001" => rgb <= "111111";
					when "10111100001011010" => rgb <= "111111";
					when "10111100001011011" => rgb <= "101010";
					when "10111100001011100" => rgb <= "111111";
					when "10111100001011101" => rgb <= "101010";
					when "10111100001011110" => rgb <= "101010";
					when "10111100001011111" => rgb <= "000000";
					when "10111100001100000" => rgb <= "000000";
					when "10111100001100001" => rgb <= "000000";
					when "10111100001100010" => rgb <= "000000";
					when "10111100001100011" => rgb <= "000000";
					when "10111100001100100" => rgb <= "000000";
					when "10111100001100101" => rgb <= "000000";
					when "10111100001100110" => rgb <= "010101";
					when "10111100001100111" => rgb <= "111111";
					when "10111100001101000" => rgb <= "101010";
					when "10111100001101001" => rgb <= "111111";
					when "10111100001101010" => rgb <= "101010";
					when "10111100001101011" => rgb <= "111111";
					when "10111100001101100" => rgb <= "101010";
					when "10111100001101101" => rgb <= "101010";
					when "10111100001101110" => rgb <= "000000";
					when "10111100001101111" => rgb <= "000000";
					when "10111100001110000" => rgb <= "000000";
					when "10111100001110001" => rgb <= "000000";
					when "10111100001110010" => rgb <= "000000";
					when "10111100001110011" => rgb <= "000000";
					when "10111100001110100" => rgb <= "000000";
					when "10111100001110101" => rgb <= "000000";
					when "10111100001110110" => rgb <= "000000";
					when "10111100001110111" => rgb <= "000000";
					when "10111100001111000" => rgb <= "000000";
					when "10111100001111001" => rgb <= "000000";
					when "10111100001111010" => rgb <= "000000";
					when "10111100001111011" => rgb <= "000000";
					when "10111100001111100" => rgb <= "000000";
					when "10111100001111101" => rgb <= "101010";
					when "10111100001111110" => rgb <= "111111";
					when "10111100001111111" => rgb <= "111111";
					when "10111100010000000" => rgb <= "111111";
					when "10111100010000001" => rgb <= "111111";
					when "10111100010000010" => rgb <= "111111";
					when "10111100010000011" => rgb <= "111111";
					when "10111100010000100" => rgb <= "111111";
					when "10111100010000101" => rgb <= "111111";
					when "10111100010000110" => rgb <= "111111";
					when "10111100010000111" => rgb <= "111111";
					when "10111100010001000" => rgb <= "111111";
					when "10111100010001001" => rgb <= "111111";
					when "10111100010001010" => rgb <= "111111";
					when "10111100010001011" => rgb <= "101010";
					when "10111100010001100" => rgb <= "000000";
					when "10111100010001101" => rgb <= "000000";
					when "10111100010001110" => rgb <= "000000";
					when "10111100010001111" => rgb <= "000000";
					when "10111100010010000" => rgb <= "000000";
					when "10111100010010001" => rgb <= "000000";
					when "10111100010010010" => rgb <= "000000";
					when "10111100010010011" => rgb <= "000000";
					when "10111100010010100" => rgb <= "000000";
					when "10111100010010101" => rgb <= "000000";
					when "10111100010010110" => rgb <= "000000";
					when "10111100010010111" => rgb <= "000000";
					when "10111100010011000" => rgb <= "000000";
					when "10111100010011001" => rgb <= "000000";
					when "10111100010011010" => rgb <= "000000";
					when "10111100010011011" => rgb <= "000000";
					when "10111100010011100" => rgb <= "000000";
					when "10111100010011101" => rgb <= "000000";
					when "10111100010011110" => rgb <= "000000";
					when "10111100010011111" => rgb <= "000000";
					when "10111100010100000" => rgb <= "000000";
					when "10111100010100001" => rgb <= "000000";
					when "10111100010100010" => rgb <= "010101";
					when "10111100010100011" => rgb <= "111111";
					when "10111100010100100" => rgb <= "101010";
					when "10111100010100101" => rgb <= "111111";
					when "10111100010100110" => rgb <= "111111";
					when "10111100010100111" => rgb <= "111111";
					when "10111100010101000" => rgb <= "111111";
					when "10111100010101001" => rgb <= "111111";
					when "10111100010101010" => rgb <= "000000";
					when "10111100010101011" => rgb <= "000000";
					when "10111100010101100" => rgb <= "000000";
					when "10111100010101101" => rgb <= "000000";
					when "10111100010101110" => rgb <= "000000";
					when "10111100010101111" => rgb <= "000000";
					when "10111100010110000" => rgb <= "000000";
					when "10111100010110001" => rgb <= "010101";
					when "10111100010110010" => rgb <= "101010";
					when "10111100010110011" => rgb <= "101010";
					when "10111100010110100" => rgb <= "111111";
					when "10111100010110101" => rgb <= "111111";
					when "10111100010110110" => rgb <= "101010";
					when "10111100010110111" => rgb <= "111111";
					when "10111100010111000" => rgb <= "101010";
					when "10111100010111001" => rgb <= "000000";
					when "10111100010111010" => rgb <= "000000";
					when "10111100010111011" => rgb <= "000000";
					when "10111100010111100" => rgb <= "000000";
					when "10111100010111101" => rgb <= "000000";
					when "10111100010111110" => rgb <= "000000";
					when "10111100010111111" => rgb <= "000000";
					when "10111100011000000" => rgb <= "010101";
					when "10111100011000001" => rgb <= "101010";
					when "10111100011000010" => rgb <= "101010";
					when "10111100011000011" => rgb <= "111111";
					when "10111100011000100" => rgb <= "111111";
					when "10111100011000101" => rgb <= "111111";
					when "10111100011000110" => rgb <= "111111";
					when "10111100011000111" => rgb <= "111111";
					when "10111100011001000" => rgb <= "111111";
					when "10111100011001001" => rgb <= "111111";
					when "10111100011001010" => rgb <= "111111";
					when "10111100011001011" => rgb <= "101010";
					when "10111100011001100" => rgb <= "111111";
					when "10111100011001101" => rgb <= "101010";
					when "10111100011001110" => rgb <= "111111";
					when "10111100011001111" => rgb <= "101010";
					when "10111100011010000" => rgb <= "000000";
					when "10111100011010001" => rgb <= "000000";
					when "10111100011010010" => rgb <= "000000";
					when "10111100011010011" => rgb <= "000000";
					when "10111100011010100" => rgb <= "000000";
					when "10111100011010101" => rgb <= "000000";
					when "10111100011010110" => rgb <= "000000";
					when "10111100011010111" => rgb <= "101010";
					when "10111100011011000" => rgb <= "101010";
					when "10111100011011001" => rgb <= "101010";
					when "10111100011011010" => rgb <= "101010";
					when "10111100011011011" => rgb <= "111111";
					when "10111100011011100" => rgb <= "111111";
					when "10111100011011101" => rgb <= "111111";
					when "10111100011011110" => rgb <= "111111";
					when "10111100011011111" => rgb <= "111111";
					when "10111100011100000" => rgb <= "111111";
					when "10111100011100001" => rgb <= "111111";
					when "10111100011100010" => rgb <= "111111";
					when "10111100011100011" => rgb <= "101010";
					when "10111100011100100" => rgb <= "111111";
					when "10111100011100101" => rgb <= "111111";
					when "10111100011100110" => rgb <= "000000";
					when "10111100011100111" => rgb <= "000000";
					when "10111100011101000" => rgb <= "000000";
					when "10111100011101001" => rgb <= "000000";
					when "10111100011101010" => rgb <= "000000";
					when "10111100011101011" => rgb <= "000000";
					when "10111100011101100" => rgb <= "000000";
					when "10111100011101101" => rgb <= "010101";
					when "10111100011101110" => rgb <= "111111";
					when "10111100011101111" => rgb <= "101010";
					when "10111100011110000" => rgb <= "111111";
					when "10111100011110001" => rgb <= "111111";
					when "10111100011110010" => rgb <= "111111";
					when "10111100011110011" => rgb <= "101010";
					when "10111100011110100" => rgb <= "101010";
					when "10111100011110101" => rgb <= "000000";
					when "10111100011110110" => rgb <= "000000";
					when "10111100011110111" => rgb <= "000000";
					when "10111100011111000" => rgb <= "000000";
					when "10111100011111001" => rgb <= "000000";
					when "10111100011111010" => rgb <= "000000";
					when "10111100011111011" => rgb <= "000000";
					when "10111100011111100" => rgb <= "000000";
					when "10111100011111101" => rgb <= "000000";
					when "10111100011111110" => rgb <= "000000";
					when "10111100011111111" => rgb <= "000000";
					when "10111100100000000" => rgb <= "000000";
					when "10111100100000001" => rgb <= "000000";
					when "10111100100000010" => rgb <= "000000";
					when "10111100100000011" => rgb <= "000000";
					when "10111100100000100" => rgb <= "101010";
					when "10111100100000101" => rgb <= "101010";
					when "10111100100000110" => rgb <= "111111";
					when "10111100100000111" => rgb <= "101010";
					when "10111100100001000" => rgb <= "101010";
					when "10111100100001001" => rgb <= "101010";
					when "10111100100001010" => rgb <= "111111";
					when "10111100100001011" => rgb <= "111111";
					when "10111100100001100" => rgb <= "101010";
					when "10111100100001101" => rgb <= "111111";
					when "10111100100001110" => rgb <= "101010";
					when "10111100100001111" => rgb <= "111111";
					when "10111100100010000" => rgb <= "111111";
					when "10111100100010001" => rgb <= "111111";
					when "10111100100010010" => rgb <= "111111";
					when "10111100100010011" => rgb <= "111111";
					when "10111100100010100" => rgb <= "111111";
					when "10111100100010101" => rgb <= "111111";
					when "10111100100010110" => rgb <= "111111";
					when "10111100100010111" => rgb <= "111111";
					when "10111100100011000" => rgb <= "101010";
					when "10111100100011001" => rgb <= "111111";
					when "10111100100011010" => rgb <= "101010";
					when "10111100100011011" => rgb <= "000000";
					when "10111100100011100" => rgb <= "000000";
					when "10111100100011101" => rgb <= "000000";
					when "10111100100011110" => rgb <= "000000";
					when "10111100100011111" => rgb <= "000000";
					when "10111100100100000" => rgb <= "000000";
					when "10111100100100001" => rgb <= "000000";
					when "10111100100100010" => rgb <= "101010";
					when "10111100100100011" => rgb <= "101010";
					when "10111100100100100" => rgb <= "101010";
					when "10111100100100101" => rgb <= "111111";
					when "10111100100100110" => rgb <= "111111";
					when "10111100100100111" => rgb <= "111111";
					when "10111100100101000" => rgb <= "111111";
					when "10111100100101001" => rgb <= "111111";
					when "10111100100101010" => rgb <= "111111";
					when "10111100100101011" => rgb <= "111111";
					when "10111100100101100" => rgb <= "111111";
					when "10111100100101101" => rgb <= "111111";
					when "10111100100101110" => rgb <= "101010";
					when "10111100100101111" => rgb <= "101010";
					when "10111100100110000" => rgb <= "111111";
					when "10111100100110001" => rgb <= "010101";
					when "10111100100110010" => rgb <= "000000";
					when "10111100100110011" => rgb <= "000000";
					when "10111100100110100" => rgb <= "000000";
					when "10111100100110101" => rgb <= "000000";
					when "10111100100110110" => rgb <= "000000";
					when "10111100100110111" => rgb <= "000000";
					when "10111100100111000" => rgb <= "000000";
					when "10111100100111001" => rgb <= "000000";
					when "10111100100111010" => rgb <= "000000";
					when "10111100100111011" => rgb <= "000000";
					when "10111100100111100" => rgb <= "000000";
					when "10111100100111101" => rgb <= "000000";
					when "10111100100111110" => rgb <= "000000";
					when "10111100100111111" => rgb <= "000000";
					when "10111101000000000" => rgb <= "000000";
					when "10111101000000001" => rgb <= "000000";
					when "10111101000000010" => rgb <= "000000";
					when "10111101000000011" => rgb <= "000000";
					when "10111101000000100" => rgb <= "000000";
					when "10111101000000101" => rgb <= "000000";
					when "10111101000000110" => rgb <= "000000";
					when "10111101000000111" => rgb <= "000000";
					when "10111101000001000" => rgb <= "000000";
					when "10111101000001001" => rgb <= "000000";
					when "10111101000001010" => rgb <= "000000";
					when "10111101000001011" => rgb <= "000000";
					when "10111101000001100" => rgb <= "010101";
					when "10111101000001101" => rgb <= "111111";
					when "10111101000001110" => rgb <= "101010";
					when "10111101000001111" => rgb <= "111111";
					when "10111101000010000" => rgb <= "111111";
					when "10111101000010001" => rgb <= "101010";
					when "10111101000010010" => rgb <= "101010";
					when "10111101000010011" => rgb <= "111111";
					when "10111101000010100" => rgb <= "101010";
					when "10111101000010101" => rgb <= "101010";
					when "10111101000010110" => rgb <= "101010";
					when "10111101000010111" => rgb <= "101010";
					when "10111101000011000" => rgb <= "111111";
					when "10111101000011001" => rgb <= "111111";
					when "10111101000011010" => rgb <= "111111";
					when "10111101000011011" => rgb <= "111111";
					when "10111101000011100" => rgb <= "111111";
					when "10111101000011101" => rgb <= "111111";
					when "10111101000011110" => rgb <= "111111";
					when "10111101000011111" => rgb <= "111111";
					when "10111101000100000" => rgb <= "111111";
					when "10111101000100001" => rgb <= "101010";
					when "10111101000100010" => rgb <= "101010";
					when "10111101000100011" => rgb <= "111111";
					when "10111101000100100" => rgb <= "111111";
					when "10111101000100101" => rgb <= "101010";
					when "10111101000100110" => rgb <= "101010";
					when "10111101000100111" => rgb <= "111111";
					when "10111101000101000" => rgb <= "101010";
					when "10111101000101001" => rgb <= "111111";
					when "10111101000101010" => rgb <= "101010";
					when "10111101000101011" => rgb <= "000000";
					when "10111101000101100" => rgb <= "000000";
					when "10111101000101101" => rgb <= "000000";
					when "10111101000101110" => rgb <= "000000";
					when "10111101000101111" => rgb <= "000000";
					when "10111101000110000" => rgb <= "000000";
					when "10111101000110001" => rgb <= "000000";
					when "10111101000110010" => rgb <= "000000";
					when "10111101000110011" => rgb <= "000000";
					when "10111101000110100" => rgb <= "000000";
					when "10111101000110101" => rgb <= "000000";
					when "10111101000110110" => rgb <= "000000";
					when "10111101000110111" => rgb <= "000000";
					when "10111101000111000" => rgb <= "000000";
					when "10111101000111001" => rgb <= "010101";
					when "10111101000111010" => rgb <= "111111";
					when "10111101000111011" => rgb <= "101010";
					when "10111101000111100" => rgb <= "111111";
					when "10111101000111101" => rgb <= "111111";
					when "10111101000111110" => rgb <= "111111";
					when "10111101000111111" => rgb <= "111111";
					when "10111101001000000" => rgb <= "101010";
					when "10111101001000001" => rgb <= "000000";
					when "10111101001000010" => rgb <= "000000";
					when "10111101001000011" => rgb <= "000000";
					when "10111101001000100" => rgb <= "000000";
					when "10111101001000101" => rgb <= "000000";
					when "10111101001000110" => rgb <= "000000";
					when "10111101001000111" => rgb <= "000000";
					when "10111101001001000" => rgb <= "000000";
					when "10111101001001001" => rgb <= "000000";
					when "10111101001001010" => rgb <= "000000";
					when "10111101001001011" => rgb <= "000000";
					when "10111101001001100" => rgb <= "000000";
					when "10111101001001101" => rgb <= "000000";
					when "10111101001001110" => rgb <= "000000";
					when "10111101001001111" => rgb <= "000000";
					when "10111101001010000" => rgb <= "101010";
					when "10111101001010001" => rgb <= "101010";
					when "10111101001010010" => rgb <= "101010";
					when "10111101001010011" => rgb <= "101010";
					when "10111101001010100" => rgb <= "111111";
					when "10111101001010101" => rgb <= "111111";
					when "10111101001010110" => rgb <= "101010";
					when "10111101001010111" => rgb <= "111111";
					when "10111101001011000" => rgb <= "111111";
					when "10111101001011001" => rgb <= "111111";
					when "10111101001011010" => rgb <= "111111";
					when "10111101001011011" => rgb <= "101010";
					when "10111101001011100" => rgb <= "111111";
					when "10111101001011101" => rgb <= "101010";
					when "10111101001011110" => rgb <= "101010";
					when "10111101001011111" => rgb <= "000000";
					when "10111101001100000" => rgb <= "000000";
					when "10111101001100001" => rgb <= "000000";
					when "10111101001100010" => rgb <= "000000";
					when "10111101001100011" => rgb <= "000000";
					when "10111101001100100" => rgb <= "000000";
					when "10111101001100101" => rgb <= "000000";
					when "10111101001100110" => rgb <= "010101";
					when "10111101001100111" => rgb <= "111111";
					when "10111101001101000" => rgb <= "101010";
					when "10111101001101001" => rgb <= "111111";
					when "10111101001101010" => rgb <= "101010";
					when "10111101001101011" => rgb <= "111111";
					when "10111101001101100" => rgb <= "101010";
					when "10111101001101101" => rgb <= "101010";
					when "10111101001101110" => rgb <= "000000";
					when "10111101001101111" => rgb <= "000000";
					when "10111101001110000" => rgb <= "000000";
					when "10111101001110001" => rgb <= "000000";
					when "10111101001110010" => rgb <= "000000";
					when "10111101001110011" => rgb <= "000000";
					when "10111101001110100" => rgb <= "000000";
					when "10111101001110101" => rgb <= "000000";
					when "10111101001110110" => rgb <= "000000";
					when "10111101001110111" => rgb <= "000000";
					when "10111101001111000" => rgb <= "000000";
					when "10111101001111001" => rgb <= "000000";
					when "10111101001111010" => rgb <= "000000";
					when "10111101001111011" => rgb <= "000000";
					when "10111101001111100" => rgb <= "000000";
					when "10111101001111101" => rgb <= "101010";
					when "10111101001111110" => rgb <= "111111";
					when "10111101001111111" => rgb <= "111111";
					when "10111101010000000" => rgb <= "111111";
					when "10111101010000001" => rgb <= "111111";
					when "10111101010000010" => rgb <= "111111";
					when "10111101010000011" => rgb <= "111111";
					when "10111101010000100" => rgb <= "111111";
					when "10111101010000101" => rgb <= "111111";
					when "10111101010000110" => rgb <= "111111";
					when "10111101010000111" => rgb <= "111111";
					when "10111101010001000" => rgb <= "111111";
					when "10111101010001001" => rgb <= "111111";
					when "10111101010001010" => rgb <= "111111";
					when "10111101010001011" => rgb <= "101010";
					when "10111101010001100" => rgb <= "000000";
					when "10111101010001101" => rgb <= "000000";
					when "10111101010001110" => rgb <= "000000";
					when "10111101010001111" => rgb <= "000000";
					when "10111101010010000" => rgb <= "000000";
					when "10111101010010001" => rgb <= "000000";
					when "10111101010010010" => rgb <= "000000";
					when "10111101010010011" => rgb <= "000000";
					when "10111101010010100" => rgb <= "000000";
					when "10111101010010101" => rgb <= "000000";
					when "10111101010010110" => rgb <= "000000";
					when "10111101010010111" => rgb <= "000000";
					when "10111101010011000" => rgb <= "000000";
					when "10111101010011001" => rgb <= "000000";
					when "10111101010011010" => rgb <= "000000";
					when "10111101010011011" => rgb <= "000000";
					when "10111101010011100" => rgb <= "000000";
					when "10111101010011101" => rgb <= "000000";
					when "10111101010011110" => rgb <= "000000";
					when "10111101010011111" => rgb <= "000000";
					when "10111101010100000" => rgb <= "000000";
					when "10111101010100001" => rgb <= "000000";
					when "10111101010100010" => rgb <= "010101";
					when "10111101010100011" => rgb <= "111111";
					when "10111101010100100" => rgb <= "101010";
					when "10111101010100101" => rgb <= "111111";
					when "10111101010100110" => rgb <= "111111";
					when "10111101010100111" => rgb <= "111111";
					when "10111101010101000" => rgb <= "111111";
					when "10111101010101001" => rgb <= "111111";
					when "10111101010101010" => rgb <= "000000";
					when "10111101010101011" => rgb <= "000000";
					when "10111101010101100" => rgb <= "000000";
					when "10111101010101101" => rgb <= "000000";
					when "10111101010101110" => rgb <= "000000";
					when "10111101010101111" => rgb <= "000000";
					when "10111101010110000" => rgb <= "000000";
					when "10111101010110001" => rgb <= "010101";
					when "10111101010110010" => rgb <= "101010";
					when "10111101010110011" => rgb <= "101010";
					when "10111101010110100" => rgb <= "111111";
					when "10111101010110101" => rgb <= "111111";
					when "10111101010110110" => rgb <= "101010";
					when "10111101010110111" => rgb <= "111111";
					when "10111101010111000" => rgb <= "101010";
					when "10111101010111001" => rgb <= "000000";
					when "10111101010111010" => rgb <= "000000";
					when "10111101010111011" => rgb <= "000000";
					when "10111101010111100" => rgb <= "000000";
					when "10111101010111101" => rgb <= "000000";
					when "10111101010111110" => rgb <= "000000";
					when "10111101010111111" => rgb <= "000000";
					when "10111101011000000" => rgb <= "010101";
					when "10111101011000001" => rgb <= "101010";
					when "10111101011000010" => rgb <= "101010";
					when "10111101011000011" => rgb <= "111111";
					when "10111101011000100" => rgb <= "111111";
					when "10111101011000101" => rgb <= "111111";
					when "10111101011000110" => rgb <= "111111";
					when "10111101011000111" => rgb <= "111111";
					when "10111101011001000" => rgb <= "111111";
					when "10111101011001001" => rgb <= "111111";
					when "10111101011001010" => rgb <= "111111";
					when "10111101011001011" => rgb <= "101010";
					when "10111101011001100" => rgb <= "111111";
					when "10111101011001101" => rgb <= "101010";
					when "10111101011001110" => rgb <= "111111";
					when "10111101011001111" => rgb <= "101010";
					when "10111101011010000" => rgb <= "000000";
					when "10111101011010001" => rgb <= "000000";
					when "10111101011010010" => rgb <= "000000";
					when "10111101011010011" => rgb <= "000000";
					when "10111101011010100" => rgb <= "000000";
					when "10111101011010101" => rgb <= "000000";
					when "10111101011010110" => rgb <= "000000";
					when "10111101011010111" => rgb <= "101010";
					when "10111101011011000" => rgb <= "101010";
					when "10111101011011001" => rgb <= "101010";
					when "10111101011011010" => rgb <= "101010";
					when "10111101011011011" => rgb <= "111111";
					when "10111101011011100" => rgb <= "111111";
					when "10111101011011101" => rgb <= "111111";
					when "10111101011011110" => rgb <= "111111";
					when "10111101011011111" => rgb <= "111111";
					when "10111101011100000" => rgb <= "111111";
					when "10111101011100001" => rgb <= "111111";
					when "10111101011100010" => rgb <= "111111";
					when "10111101011100011" => rgb <= "101010";
					when "10111101011100100" => rgb <= "111111";
					when "10111101011100101" => rgb <= "111111";
					when "10111101011100110" => rgb <= "000000";
					when "10111101011100111" => rgb <= "000000";
					when "10111101011101000" => rgb <= "000000";
					when "10111101011101001" => rgb <= "000000";
					when "10111101011101010" => rgb <= "000000";
					when "10111101011101011" => rgb <= "000000";
					when "10111101011101100" => rgb <= "000000";
					when "10111101011101101" => rgb <= "010101";
					when "10111101011101110" => rgb <= "111111";
					when "10111101011101111" => rgb <= "101010";
					when "10111101011110000" => rgb <= "111111";
					when "10111101011110001" => rgb <= "111111";
					when "10111101011110010" => rgb <= "111111";
					when "10111101011110011" => rgb <= "101010";
					when "10111101011110100" => rgb <= "101010";
					when "10111101011110101" => rgb <= "000000";
					when "10111101011110110" => rgb <= "000000";
					when "10111101011110111" => rgb <= "000000";
					when "10111101011111000" => rgb <= "000000";
					when "10111101011111001" => rgb <= "000000";
					when "10111101011111010" => rgb <= "000000";
					when "10111101011111011" => rgb <= "000000";
					when "10111101011111100" => rgb <= "000000";
					when "10111101011111101" => rgb <= "000000";
					when "10111101011111110" => rgb <= "000000";
					when "10111101011111111" => rgb <= "000000";
					when "10111101100000000" => rgb <= "000000";
					when "10111101100000001" => rgb <= "000000";
					when "10111101100000010" => rgb <= "000000";
					when "10111101100000011" => rgb <= "000000";
					when "10111101100000100" => rgb <= "101010";
					when "10111101100000101" => rgb <= "111111";
					when "10111101100000110" => rgb <= "111111";
					when "10111101100000111" => rgb <= "111111";
					when "10111101100001000" => rgb <= "111111";
					when "10111101100001001" => rgb <= "111111";
					when "10111101100001010" => rgb <= "111111";
					when "10111101100001011" => rgb <= "101010";
					when "10111101100001100" => rgb <= "101010";
					when "10111101100001101" => rgb <= "111111";
					when "10111101100001110" => rgb <= "111111";
					when "10111101100001111" => rgb <= "111111";
					when "10111101100010000" => rgb <= "111111";
					when "10111101100010001" => rgb <= "111111";
					when "10111101100010010" => rgb <= "111111";
					when "10111101100010011" => rgb <= "111111";
					when "10111101100010100" => rgb <= "111111";
					when "10111101100010101" => rgb <= "111111";
					when "10111101100010110" => rgb <= "111111";
					when "10111101100010111" => rgb <= "111111";
					when "10111101100011000" => rgb <= "101010";
					when "10111101100011001" => rgb <= "111111";
					when "10111101100011010" => rgb <= "101010";
					when "10111101100011011" => rgb <= "000000";
					when "10111101100011100" => rgb <= "000000";
					when "10111101100011101" => rgb <= "000000";
					when "10111101100011110" => rgb <= "000000";
					when "10111101100011111" => rgb <= "000000";
					when "10111101100100000" => rgb <= "000000";
					when "10111101100100001" => rgb <= "000000";
					when "10111101100100010" => rgb <= "101010";
					when "10111101100100011" => rgb <= "101010";
					when "10111101100100100" => rgb <= "101010";
					when "10111101100100101" => rgb <= "111111";
					when "10111101100100110" => rgb <= "111111";
					when "10111101100100111" => rgb <= "111111";
					when "10111101100101000" => rgb <= "111111";
					when "10111101100101001" => rgb <= "111111";
					when "10111101100101010" => rgb <= "111111";
					when "10111101100101011" => rgb <= "111111";
					when "10111101100101100" => rgb <= "111111";
					when "10111101100101101" => rgb <= "111111";
					when "10111101100101110" => rgb <= "101010";
					when "10111101100101111" => rgb <= "101010";
					when "10111101100110000" => rgb <= "111111";
					when "10111101100110001" => rgb <= "010101";
					when "10111101100110010" => rgb <= "000000";
					when "10111101100110011" => rgb <= "000000";
					when "10111101100110100" => rgb <= "000000";
					when "10111101100110101" => rgb <= "000000";
					when "10111101100110110" => rgb <= "000000";
					when "10111101100110111" => rgb <= "000000";
					when "10111101100111000" => rgb <= "000000";
					when "10111101100111001" => rgb <= "000000";
					when "10111101100111010" => rgb <= "000000";
					when "10111101100111011" => rgb <= "000000";
					when "10111101100111100" => rgb <= "000000";
					when "10111101100111101" => rgb <= "000000";
					when "10111101100111110" => rgb <= "000000";
					when "10111101100111111" => rgb <= "000000";
					when "10111110000000000" => rgb <= "000000";
					when "10111110000000001" => rgb <= "000000";
					when "10111110000000010" => rgb <= "000000";
					when "10111110000000011" => rgb <= "000000";
					when "10111110000000100" => rgb <= "000000";
					when "10111110000000101" => rgb <= "000000";
					when "10111110000000110" => rgb <= "000000";
					when "10111110000000111" => rgb <= "000000";
					when "10111110000001000" => rgb <= "000000";
					when "10111110000001001" => rgb <= "000000";
					when "10111110000001010" => rgb <= "000000";
					when "10111110000001011" => rgb <= "000000";
					when "10111110000001100" => rgb <= "010101";
					when "10111110000001101" => rgb <= "101010";
					when "10111110000001110" => rgb <= "101010";
					when "10111110000001111" => rgb <= "101010";
					when "10111110000010000" => rgb <= "101010";
					when "10111110000010001" => rgb <= "101010";
					when "10111110000010010" => rgb <= "101010";
					when "10111110000010011" => rgb <= "101010";
					when "10111110000010100" => rgb <= "101010";
					when "10111110000010101" => rgb <= "101010";
					when "10111110000010110" => rgb <= "111111";
					when "10111110000010111" => rgb <= "111111";
					when "10111110000011000" => rgb <= "101010";
					when "10111110000011001" => rgb <= "101010";
					when "10111110000011010" => rgb <= "111111";
					when "10111110000011011" => rgb <= "111111";
					when "10111110000011100" => rgb <= "111111";
					when "10111110000011101" => rgb <= "111111";
					when "10111110000011110" => rgb <= "111111";
					when "10111110000011111" => rgb <= "111111";
					when "10111110000100000" => rgb <= "101010";
					when "10111110000100001" => rgb <= "101010";
					when "10111110000100010" => rgb <= "111111";
					when "10111110000100011" => rgb <= "101010";
					when "10111110000100100" => rgb <= "101010";
					when "10111110000100101" => rgb <= "101010";
					when "10111110000100110" => rgb <= "101010";
					when "10111110000100111" => rgb <= "101010";
					when "10111110000101000" => rgb <= "101010";
					when "10111110000101001" => rgb <= "101010";
					when "10111110000101010" => rgb <= "010101";
					when "10111110000101011" => rgb <= "000000";
					when "10111110000101100" => rgb <= "000000";
					when "10111110000101101" => rgb <= "000000";
					when "10111110000101110" => rgb <= "000000";
					when "10111110000101111" => rgb <= "000000";
					when "10111110000110000" => rgb <= "000000";
					when "10111110000110001" => rgb <= "000000";
					when "10111110000110010" => rgb <= "000000";
					when "10111110000110011" => rgb <= "000000";
					when "10111110000110100" => rgb <= "000000";
					when "10111110000110101" => rgb <= "000000";
					when "10111110000110110" => rgb <= "000000";
					when "10111110000110111" => rgb <= "000000";
					when "10111110000111000" => rgb <= "000000";
					when "10111110000111001" => rgb <= "010101";
					when "10111110000111010" => rgb <= "111111";
					when "10111110000111011" => rgb <= "101010";
					when "10111110000111100" => rgb <= "111111";
					when "10111110000111101" => rgb <= "111111";
					when "10111110000111110" => rgb <= "111111";
					when "10111110000111111" => rgb <= "111111";
					when "10111110001000000" => rgb <= "101010";
					when "10111110001000001" => rgb <= "000000";
					when "10111110001000010" => rgb <= "000000";
					when "10111110001000011" => rgb <= "000000";
					when "10111110001000100" => rgb <= "000000";
					when "10111110001000101" => rgb <= "000000";
					when "10111110001000110" => rgb <= "000000";
					when "10111110001000111" => rgb <= "000000";
					when "10111110001001000" => rgb <= "000000";
					when "10111110001001001" => rgb <= "000000";
					when "10111110001001010" => rgb <= "000000";
					when "10111110001001011" => rgb <= "000000";
					when "10111110001001100" => rgb <= "000000";
					when "10111110001001101" => rgb <= "000000";
					when "10111110001001110" => rgb <= "000000";
					when "10111110001001111" => rgb <= "000000";
					when "10111110001010000" => rgb <= "101010";
					when "10111110001010001" => rgb <= "101010";
					when "10111110001010010" => rgb <= "101010";
					when "10111110001010011" => rgb <= "101010";
					when "10111110001010100" => rgb <= "111111";
					when "10111110001010101" => rgb <= "111111";
					when "10111110001010110" => rgb <= "101010";
					when "10111110001010111" => rgb <= "111111";
					when "10111110001011000" => rgb <= "111111";
					when "10111110001011001" => rgb <= "111111";
					when "10111110001011010" => rgb <= "111111";
					when "10111110001011011" => rgb <= "101010";
					when "10111110001011100" => rgb <= "111111";
					when "10111110001011101" => rgb <= "101010";
					when "10111110001011110" => rgb <= "101010";
					when "10111110001011111" => rgb <= "000000";
					when "10111110001100000" => rgb <= "000000";
					when "10111110001100001" => rgb <= "000000";
					when "10111110001100010" => rgb <= "000000";
					when "10111110001100011" => rgb <= "000000";
					when "10111110001100100" => rgb <= "000000";
					when "10111110001100101" => rgb <= "000000";
					when "10111110001100110" => rgb <= "010101";
					when "10111110001100111" => rgb <= "111111";
					when "10111110001101000" => rgb <= "101010";
					when "10111110001101001" => rgb <= "111111";
					when "10111110001101010" => rgb <= "101010";
					when "10111110001101011" => rgb <= "111111";
					when "10111110001101100" => rgb <= "101010";
					when "10111110001101101" => rgb <= "101010";
					when "10111110001101110" => rgb <= "000000";
					when "10111110001101111" => rgb <= "000000";
					when "10111110001110000" => rgb <= "000000";
					when "10111110001110001" => rgb <= "000000";
					when "10111110001110010" => rgb <= "000000";
					when "10111110001110011" => rgb <= "000000";
					when "10111110001110100" => rgb <= "000000";
					when "10111110001110101" => rgb <= "000000";
					when "10111110001110110" => rgb <= "000000";
					when "10111110001110111" => rgb <= "000000";
					when "10111110001111000" => rgb <= "000000";
					when "10111110001111001" => rgb <= "000000";
					when "10111110001111010" => rgb <= "000000";
					when "10111110001111011" => rgb <= "000000";
					when "10111110001111100" => rgb <= "000000";
					when "10111110001111101" => rgb <= "101010";
					when "10111110001111110" => rgb <= "111111";
					when "10111110001111111" => rgb <= "111111";
					when "10111110010000000" => rgb <= "111111";
					when "10111110010000001" => rgb <= "111111";
					when "10111110010000010" => rgb <= "111111";
					when "10111110010000011" => rgb <= "111111";
					when "10111110010000100" => rgb <= "111111";
					when "10111110010000101" => rgb <= "111111";
					when "10111110010000110" => rgb <= "111111";
					when "10111110010000111" => rgb <= "111111";
					when "10111110010001000" => rgb <= "111111";
					when "10111110010001001" => rgb <= "111111";
					when "10111110010001010" => rgb <= "111111";
					when "10111110010001011" => rgb <= "101010";
					when "10111110010001100" => rgb <= "000000";
					when "10111110010001101" => rgb <= "000000";
					when "10111110010001110" => rgb <= "000000";
					when "10111110010001111" => rgb <= "000000";
					when "10111110010010000" => rgb <= "000000";
					when "10111110010010001" => rgb <= "000000";
					when "10111110010010010" => rgb <= "000000";
					when "10111110010010011" => rgb <= "000000";
					when "10111110010010100" => rgb <= "000000";
					when "10111110010010101" => rgb <= "000000";
					when "10111110010010110" => rgb <= "000000";
					when "10111110010010111" => rgb <= "000000";
					when "10111110010011000" => rgb <= "000000";
					when "10111110010011001" => rgb <= "000000";
					when "10111110010011010" => rgb <= "000000";
					when "10111110010011011" => rgb <= "000000";
					when "10111110010011100" => rgb <= "000000";
					when "10111110010011101" => rgb <= "000000";
					when "10111110010011110" => rgb <= "000000";
					when "10111110010011111" => rgb <= "000000";
					when "10111110010100000" => rgb <= "000000";
					when "10111110010100001" => rgb <= "000000";
					when "10111110010100010" => rgb <= "010101";
					when "10111110010100011" => rgb <= "111111";
					when "10111110010100100" => rgb <= "101010";
					when "10111110010100101" => rgb <= "111111";
					when "10111110010100110" => rgb <= "111111";
					when "10111110010100111" => rgb <= "111111";
					when "10111110010101000" => rgb <= "111111";
					when "10111110010101001" => rgb <= "111111";
					when "10111110010101010" => rgb <= "000000";
					when "10111110010101011" => rgb <= "000000";
					when "10111110010101100" => rgb <= "000000";
					when "10111110010101101" => rgb <= "000000";
					when "10111110010101110" => rgb <= "000000";
					when "10111110010101111" => rgb <= "000000";
					when "10111110010110000" => rgb <= "000000";
					when "10111110010110001" => rgb <= "010101";
					when "10111110010110010" => rgb <= "101010";
					when "10111110010110011" => rgb <= "101010";
					when "10111110010110100" => rgb <= "111111";
					when "10111110010110101" => rgb <= "111111";
					when "10111110010110110" => rgb <= "111111";
					when "10111110010110111" => rgb <= "111111";
					when "10111110010111000" => rgb <= "101010";
					when "10111110010111001" => rgb <= "000000";
					when "10111110010111010" => rgb <= "000000";
					when "10111110010111011" => rgb <= "000000";
					when "10111110010111100" => rgb <= "000000";
					when "10111110010111101" => rgb <= "000000";
					when "10111110010111110" => rgb <= "000000";
					when "10111110010111111" => rgb <= "000000";
					when "10111110011000000" => rgb <= "010101";
					when "10111110011000001" => rgb <= "111111";
					when "10111110011000010" => rgb <= "101010";
					when "10111110011000011" => rgb <= "111111";
					when "10111110011000100" => rgb <= "101010";
					when "10111110011000101" => rgb <= "111111";
					when "10111110011000110" => rgb <= "111111";
					when "10111110011000111" => rgb <= "111111";
					when "10111110011001000" => rgb <= "111111";
					when "10111110011001001" => rgb <= "111111";
					when "10111110011001010" => rgb <= "111111";
					when "10111110011001011" => rgb <= "101010";
					when "10111110011001100" => rgb <= "111111";
					when "10111110011001101" => rgb <= "101010";
					when "10111110011001110" => rgb <= "111111";
					when "10111110011001111" => rgb <= "101010";
					when "10111110011010000" => rgb <= "000000";
					when "10111110011010001" => rgb <= "000000";
					when "10111110011010010" => rgb <= "000000";
					when "10111110011010011" => rgb <= "000000";
					when "10111110011010100" => rgb <= "000000";
					when "10111110011010101" => rgb <= "000000";
					when "10111110011010110" => rgb <= "000000";
					when "10111110011010111" => rgb <= "101010";
					when "10111110011011000" => rgb <= "101010";
					when "10111110011011001" => rgb <= "101010";
					when "10111110011011010" => rgb <= "101010";
					when "10111110011011011" => rgb <= "111111";
					when "10111110011011100" => rgb <= "111111";
					when "10111110011011101" => rgb <= "111111";
					when "10111110011011110" => rgb <= "111111";
					when "10111110011011111" => rgb <= "111111";
					when "10111110011100000" => rgb <= "111111";
					when "10111110011100001" => rgb <= "111111";
					when "10111110011100010" => rgb <= "111111";
					when "10111110011100011" => rgb <= "101010";
					when "10111110011100100" => rgb <= "111111";
					when "10111110011100101" => rgb <= "111111";
					when "10111110011100110" => rgb <= "000000";
					when "10111110011100111" => rgb <= "000000";
					when "10111110011101000" => rgb <= "000000";
					when "10111110011101001" => rgb <= "000000";
					when "10111110011101010" => rgb <= "000000";
					when "10111110011101011" => rgb <= "000000";
					when "10111110011101100" => rgb <= "000000";
					when "10111110011101101" => rgb <= "010101";
					when "10111110011101110" => rgb <= "111111";
					when "10111110011101111" => rgb <= "101010";
					when "10111110011110000" => rgb <= "111111";
					when "10111110011110001" => rgb <= "111111";
					when "10111110011110010" => rgb <= "111111";
					when "10111110011110011" => rgb <= "101010";
					when "10111110011110100" => rgb <= "101010";
					when "10111110011110101" => rgb <= "000000";
					when "10111110011110110" => rgb <= "000000";
					when "10111110011110111" => rgb <= "000000";
					when "10111110011111000" => rgb <= "000000";
					when "10111110011111001" => rgb <= "000000";
					when "10111110011111010" => rgb <= "000000";
					when "10111110011111011" => rgb <= "000000";
					when "10111110011111100" => rgb <= "000000";
					when "10111110011111101" => rgb <= "000000";
					when "10111110011111110" => rgb <= "000000";
					when "10111110011111111" => rgb <= "000000";
					when "10111110100000000" => rgb <= "000000";
					when "10111110100000001" => rgb <= "000000";
					when "10111110100000010" => rgb <= "000000";
					when "10111110100000011" => rgb <= "000000";
					when "10111110100000100" => rgb <= "101010";
					when "10111110100000101" => rgb <= "101010";
					when "10111110100000110" => rgb <= "101010";
					when "10111110100000111" => rgb <= "101010";
					when "10111110100001000" => rgb <= "101010";
					when "10111110100001001" => rgb <= "101010";
					when "10111110100001010" => rgb <= "101010";
					when "10111110100001011" => rgb <= "101010";
					when "10111110100001100" => rgb <= "111111";
					when "10111110100001101" => rgb <= "101010";
					when "10111110100001110" => rgb <= "101010";
					when "10111110100001111" => rgb <= "101010";
					when "10111110100010000" => rgb <= "111111";
					when "10111110100010001" => rgb <= "111111";
					when "10111110100010010" => rgb <= "111111";
					when "10111110100010011" => rgb <= "111111";
					when "10111110100010100" => rgb <= "111111";
					when "10111110100010101" => rgb <= "111111";
					when "10111110100010110" => rgb <= "111111";
					when "10111110100010111" => rgb <= "111111";
					when "10111110100011000" => rgb <= "101010";
					when "10111110100011001" => rgb <= "111111";
					when "10111110100011010" => rgb <= "101010";
					when "10111110100011011" => rgb <= "000000";
					when "10111110100011100" => rgb <= "000000";
					when "10111110100011101" => rgb <= "000000";
					when "10111110100011110" => rgb <= "000000";
					when "10111110100011111" => rgb <= "000000";
					when "10111110100100000" => rgb <= "000000";
					when "10111110100100001" => rgb <= "000000";
					when "10111110100100010" => rgb <= "101010";
					when "10111110100100011" => rgb <= "101010";
					when "10111110100100100" => rgb <= "101010";
					when "10111110100100101" => rgb <= "111111";
					when "10111110100100110" => rgb <= "111111";
					when "10111110100100111" => rgb <= "111111";
					when "10111110100101000" => rgb <= "111111";
					when "10111110100101001" => rgb <= "111111";
					when "10111110100101010" => rgb <= "111111";
					when "10111110100101011" => rgb <= "111111";
					when "10111110100101100" => rgb <= "111111";
					when "10111110100101101" => rgb <= "111111";
					when "10111110100101110" => rgb <= "101010";
					when "10111110100101111" => rgb <= "101010";
					when "10111110100110000" => rgb <= "111111";
					when "10111110100110001" => rgb <= "010101";
					when "10111110100110010" => rgb <= "000000";
					when "10111110100110011" => rgb <= "000000";
					when "10111110100110100" => rgb <= "000000";
					when "10111110100110101" => rgb <= "000000";
					when "10111110100110110" => rgb <= "000000";
					when "10111110100110111" => rgb <= "000000";
					when "10111110100111000" => rgb <= "000000";
					when "10111110100111001" => rgb <= "000000";
					when "10111110100111010" => rgb <= "000000";
					when "10111110100111011" => rgb <= "000000";
					when "10111110100111100" => rgb <= "000000";
					when "10111110100111101" => rgb <= "000000";
					when "10111110100111110" => rgb <= "000000";
					when "10111110100111111" => rgb <= "000000";
					when "10111111000000000" => rgb <= "000000";
					when "10111111000000001" => rgb <= "000000";
					when "10111111000000010" => rgb <= "000000";
					when "10111111000000011" => rgb <= "000000";
					when "10111111000000100" => rgb <= "000000";
					when "10111111000000101" => rgb <= "000000";
					when "10111111000000110" => rgb <= "000000";
					when "10111111000000111" => rgb <= "000000";
					when "10111111000001000" => rgb <= "000000";
					when "10111111000001001" => rgb <= "000000";
					when "10111111000001010" => rgb <= "000000";
					when "10111111000001011" => rgb <= "000000";
					when "10111111000001100" => rgb <= "000000";
					when "10111111000001101" => rgb <= "000000";
					when "10111111000001110" => rgb <= "000000";
					when "10111111000001111" => rgb <= "000000";
					when "10111111000010000" => rgb <= "000000";
					when "10111111000010001" => rgb <= "000000";
					when "10111111000010010" => rgb <= "000000";
					when "10111111000010011" => rgb <= "000000";
					when "10111111000010100" => rgb <= "101010";
					when "10111111000010101" => rgb <= "111111";
					when "10111111000010110" => rgb <= "111111";
					when "10111111000010111" => rgb <= "101010";
					when "10111111000011000" => rgb <= "111111";
					when "10111111000011001" => rgb <= "111111";
					when "10111111000011010" => rgb <= "111111";
					when "10111111000011011" => rgb <= "111111";
					when "10111111000011100" => rgb <= "111111";
					when "10111111000011101" => rgb <= "111111";
					when "10111111000011110" => rgb <= "111111";
					when "10111111000011111" => rgb <= "111111";
					when "10111111000100000" => rgb <= "111111";
					when "10111111000100001" => rgb <= "101010";
					when "10111111000100010" => rgb <= "101010";
					when "10111111000100011" => rgb <= "000000";
					when "10111111000100100" => rgb <= "000000";
					when "10111111000100101" => rgb <= "000000";
					when "10111111000100110" => rgb <= "000000";
					when "10111111000100111" => rgb <= "000000";
					when "10111111000101000" => rgb <= "000000";
					when "10111111000101001" => rgb <= "000000";
					when "10111111000101010" => rgb <= "000000";
					when "10111111000101011" => rgb <= "000000";
					when "10111111000101100" => rgb <= "000000";
					when "10111111000101101" => rgb <= "000000";
					when "10111111000101110" => rgb <= "000000";
					when "10111111000101111" => rgb <= "000000";
					when "10111111000110000" => rgb <= "000000";
					when "10111111000110001" => rgb <= "000000";
					when "10111111000110010" => rgb <= "000000";
					when "10111111000110011" => rgb <= "000000";
					when "10111111000110100" => rgb <= "000000";
					when "10111111000110101" => rgb <= "000000";
					when "10111111000110110" => rgb <= "000000";
					when "10111111000110111" => rgb <= "000000";
					when "10111111000111000" => rgb <= "000000";
					when "10111111000111001" => rgb <= "010101";
					when "10111111000111010" => rgb <= "101010";
					when "10111111000111011" => rgb <= "101010";
					when "10111111000111100" => rgb <= "111111";
					when "10111111000111101" => rgb <= "111111";
					when "10111111000111110" => rgb <= "101010";
					when "10111111000111111" => rgb <= "111111";
					when "10111111001000000" => rgb <= "101010";
					when "10111111001000001" => rgb <= "000000";
					when "10111111001000010" => rgb <= "000000";
					when "10111111001000011" => rgb <= "000000";
					when "10111111001000100" => rgb <= "000000";
					when "10111111001000101" => rgb <= "000000";
					when "10111111001000110" => rgb <= "000000";
					when "10111111001000111" => rgb <= "000000";
					when "10111111001001000" => rgb <= "000000";
					when "10111111001001001" => rgb <= "000000";
					when "10111111001001010" => rgb <= "000000";
					when "10111111001001011" => rgb <= "000000";
					when "10111111001001100" => rgb <= "000000";
					when "10111111001001101" => rgb <= "000000";
					when "10111111001001110" => rgb <= "000000";
					when "10111111001001111" => rgb <= "000000";
					when "10111111001010000" => rgb <= "101010";
					when "10111111001010001" => rgb <= "101010";
					when "10111111001010010" => rgb <= "101010";
					when "10111111001010011" => rgb <= "101010";
					when "10111111001010100" => rgb <= "111111";
					when "10111111001010101" => rgb <= "111111";
					when "10111111001010110" => rgb <= "101010";
					when "10111111001010111" => rgb <= "111111";
					when "10111111001011000" => rgb <= "111111";
					when "10111111001011001" => rgb <= "111111";
					when "10111111001011010" => rgb <= "111111";
					when "10111111001011011" => rgb <= "101010";
					when "10111111001011100" => rgb <= "111111";
					when "10111111001011101" => rgb <= "101010";
					when "10111111001011110" => rgb <= "101010";
					when "10111111001011111" => rgb <= "000000";
					when "10111111001100000" => rgb <= "000000";
					when "10111111001100001" => rgb <= "000000";
					when "10111111001100010" => rgb <= "000000";
					when "10111111001100011" => rgb <= "000000";
					when "10111111001100100" => rgb <= "000000";
					when "10111111001100101" => rgb <= "000000";
					when "10111111001100110" => rgb <= "010101";
					when "10111111001100111" => rgb <= "111111";
					when "10111111001101000" => rgb <= "101010";
					when "10111111001101001" => rgb <= "111111";
					when "10111111001101010" => rgb <= "101010";
					when "10111111001101011" => rgb <= "111111";
					when "10111111001101100" => rgb <= "101010";
					when "10111111001101101" => rgb <= "101010";
					when "10111111001101110" => rgb <= "000000";
					when "10111111001101111" => rgb <= "000000";
					when "10111111001110000" => rgb <= "000000";
					when "10111111001110001" => rgb <= "000000";
					when "10111111001110010" => rgb <= "000000";
					when "10111111001110011" => rgb <= "000000";
					when "10111111001110100" => rgb <= "000000";
					when "10111111001110101" => rgb <= "000000";
					when "10111111001110110" => rgb <= "000000";
					when "10111111001110111" => rgb <= "000000";
					when "10111111001111000" => rgb <= "000000";
					when "10111111001111001" => rgb <= "000000";
					when "10111111001111010" => rgb <= "000000";
					when "10111111001111011" => rgb <= "000000";
					when "10111111001111100" => rgb <= "000000";
					when "10111111001111101" => rgb <= "101010";
					when "10111111001111110" => rgb <= "111111";
					when "10111111001111111" => rgb <= "111111";
					when "10111111010000000" => rgb <= "111111";
					when "10111111010000001" => rgb <= "111111";
					when "10111111010000010" => rgb <= "111111";
					when "10111111010000011" => rgb <= "111111";
					when "10111111010000100" => rgb <= "111111";
					when "10111111010000101" => rgb <= "111111";
					when "10111111010000110" => rgb <= "111111";
					when "10111111010000111" => rgb <= "111111";
					when "10111111010001000" => rgb <= "111111";
					when "10111111010001001" => rgb <= "111111";
					when "10111111010001010" => rgb <= "111111";
					when "10111111010001011" => rgb <= "101010";
					when "10111111010001100" => rgb <= "000000";
					when "10111111010001101" => rgb <= "000000";
					when "10111111010001110" => rgb <= "000000";
					when "10111111010001111" => rgb <= "000000";
					when "10111111010010000" => rgb <= "000000";
					when "10111111010010001" => rgb <= "000000";
					when "10111111010010010" => rgb <= "000000";
					when "10111111010010011" => rgb <= "000000";
					when "10111111010010100" => rgb <= "000000";
					when "10111111010010101" => rgb <= "000000";
					when "10111111010010110" => rgb <= "000000";
					when "10111111010010111" => rgb <= "000000";
					when "10111111010011000" => rgb <= "000000";
					when "10111111010011001" => rgb <= "000000";
					when "10111111010011010" => rgb <= "000000";
					when "10111111010011011" => rgb <= "000000";
					when "10111111010011100" => rgb <= "000000";
					when "10111111010011101" => rgb <= "000000";
					when "10111111010011110" => rgb <= "000000";
					when "10111111010011111" => rgb <= "000000";
					when "10111111010100000" => rgb <= "000000";
					when "10111111010100001" => rgb <= "000000";
					when "10111111010100010" => rgb <= "010101";
					when "10111111010100011" => rgb <= "111111";
					when "10111111010100100" => rgb <= "101010";
					when "10111111010100101" => rgb <= "111111";
					when "10111111010100110" => rgb <= "111111";
					when "10111111010100111" => rgb <= "111111";
					when "10111111010101000" => rgb <= "111111";
					when "10111111010101001" => rgb <= "111111";
					when "10111111010101010" => rgb <= "000000";
					when "10111111010101011" => rgb <= "000000";
					when "10111111010101100" => rgb <= "000000";
					when "10111111010101101" => rgb <= "000000";
					when "10111111010101110" => rgb <= "000000";
					when "10111111010101111" => rgb <= "000000";
					when "10111111010110000" => rgb <= "000000";
					when "10111111010110001" => rgb <= "010101";
					when "10111111010110010" => rgb <= "101010";
					when "10111111010110011" => rgb <= "101010";
					when "10111111010110100" => rgb <= "111111";
					when "10111111010110101" => rgb <= "111111";
					when "10111111010110110" => rgb <= "101010";
					when "10111111010110111" => rgb <= "111111";
					when "10111111010111000" => rgb <= "101010";
					when "10111111010111001" => rgb <= "000000";
					when "10111111010111010" => rgb <= "000000";
					when "10111111010111011" => rgb <= "000000";
					when "10111111010111100" => rgb <= "000000";
					when "10111111010111101" => rgb <= "000000";
					when "10111111010111110" => rgb <= "000000";
					when "10111111010111111" => rgb <= "000000";
					when "10111111011000000" => rgb <= "010101";
					when "10111111011000001" => rgb <= "111111";
					when "10111111011000010" => rgb <= "101010";
					when "10111111011000011" => rgb <= "111111";
					when "10111111011000100" => rgb <= "101010";
					when "10111111011000101" => rgb <= "111111";
					when "10111111011000110" => rgb <= "111111";
					when "10111111011000111" => rgb <= "111111";
					when "10111111011001000" => rgb <= "111111";
					when "10111111011001001" => rgb <= "111111";
					when "10111111011001010" => rgb <= "111111";
					when "10111111011001011" => rgb <= "101010";
					when "10111111011001100" => rgb <= "111111";
					when "10111111011001101" => rgb <= "101010";
					when "10111111011001110" => rgb <= "111111";
					when "10111111011001111" => rgb <= "101010";
					when "10111111011010000" => rgb <= "000000";
					when "10111111011010001" => rgb <= "000000";
					when "10111111011010010" => rgb <= "000000";
					when "10111111011010011" => rgb <= "000000";
					when "10111111011010100" => rgb <= "000000";
					when "10111111011010101" => rgb <= "000000";
					when "10111111011010110" => rgb <= "000000";
					when "10111111011010111" => rgb <= "101010";
					when "10111111011011000" => rgb <= "101010";
					when "10111111011011001" => rgb <= "101010";
					when "10111111011011010" => rgb <= "101010";
					when "10111111011011011" => rgb <= "111111";
					when "10111111011011100" => rgb <= "111111";
					when "10111111011011101" => rgb <= "111111";
					when "10111111011011110" => rgb <= "111111";
					when "10111111011011111" => rgb <= "111111";
					when "10111111011100000" => rgb <= "111111";
					when "10111111011100001" => rgb <= "111111";
					when "10111111011100010" => rgb <= "111111";
					when "10111111011100011" => rgb <= "101010";
					when "10111111011100100" => rgb <= "111111";
					when "10111111011100101" => rgb <= "111111";
					when "10111111011100110" => rgb <= "000000";
					when "10111111011100111" => rgb <= "000000";
					when "10111111011101000" => rgb <= "000000";
					when "10111111011101001" => rgb <= "000000";
					when "10111111011101010" => rgb <= "000000";
					when "10111111011101011" => rgb <= "000000";
					when "10111111011101100" => rgb <= "000000";
					when "10111111011101101" => rgb <= "010101";
					when "10111111011101110" => rgb <= "111111";
					when "10111111011101111" => rgb <= "101010";
					when "10111111011110000" => rgb <= "111111";
					when "10111111011110001" => rgb <= "111111";
					when "10111111011110010" => rgb <= "111111";
					when "10111111011110011" => rgb <= "101010";
					when "10111111011110100" => rgb <= "101010";
					when "10111111011110101" => rgb <= "000000";
					when "10111111011110110" => rgb <= "000000";
					when "10111111011110111" => rgb <= "000000";
					when "10111111011111000" => rgb <= "000000";
					when "10111111011111001" => rgb <= "000000";
					when "10111111011111010" => rgb <= "000000";
					when "10111111011111011" => rgb <= "000000";
					when "10111111011111100" => rgb <= "000000";
					when "10111111011111101" => rgb <= "000000";
					when "10111111011111110" => rgb <= "000000";
					when "10111111011111111" => rgb <= "000000";
					when "10111111100000000" => rgb <= "000000";
					when "10111111100000001" => rgb <= "000000";
					when "10111111100000010" => rgb <= "000000";
					when "10111111100000011" => rgb <= "000000";
					when "10111111100000100" => rgb <= "000000";
					when "10111111100000101" => rgb <= "000000";
					when "10111111100000110" => rgb <= "000000";
					when "10111111100000111" => rgb <= "000000";
					when "10111111100001000" => rgb <= "000000";
					when "10111111100001001" => rgb <= "000000";
					when "10111111100001010" => rgb <= "000000";
					when "10111111100001011" => rgb <= "010101";
					when "10111111100001100" => rgb <= "101010";
					when "10111111100001101" => rgb <= "101010";
					when "10111111100001110" => rgb <= "101010";
					when "10111111100001111" => rgb <= "111111";
					when "10111111100010000" => rgb <= "111111";
					when "10111111100010001" => rgb <= "111111";
					when "10111111100010010" => rgb <= "111111";
					when "10111111100010011" => rgb <= "111111";
					when "10111111100010100" => rgb <= "111111";
					when "10111111100010101" => rgb <= "111111";
					when "10111111100010110" => rgb <= "111111";
					when "10111111100010111" => rgb <= "111111";
					when "10111111100011000" => rgb <= "101010";
					when "10111111100011001" => rgb <= "111111";
					when "10111111100011010" => rgb <= "101010";
					when "10111111100011011" => rgb <= "000000";
					when "10111111100011100" => rgb <= "000000";
					when "10111111100011101" => rgb <= "000000";
					when "10111111100011110" => rgb <= "000000";
					when "10111111100011111" => rgb <= "000000";
					when "10111111100100000" => rgb <= "000000";
					when "10111111100100001" => rgb <= "000000";
					when "10111111100100010" => rgb <= "101010";
					when "10111111100100011" => rgb <= "101010";
					when "10111111100100100" => rgb <= "101010";
					when "10111111100100101" => rgb <= "111111";
					when "10111111100100110" => rgb <= "111111";
					when "10111111100100111" => rgb <= "111111";
					when "10111111100101000" => rgb <= "111111";
					when "10111111100101001" => rgb <= "111111";
					when "10111111100101010" => rgb <= "111111";
					when "10111111100101011" => rgb <= "111111";
					when "10111111100101100" => rgb <= "111111";
					when "10111111100101101" => rgb <= "111111";
					when "10111111100101110" => rgb <= "101010";
					when "10111111100101111" => rgb <= "101010";
					when "10111111100110000" => rgb <= "111111";
					when "10111111100110001" => rgb <= "010101";
					when "10111111100110010" => rgb <= "000000";
					when "10111111100110011" => rgb <= "000000";
					when "10111111100110100" => rgb <= "000000";
					when "10111111100110101" => rgb <= "000000";
					when "10111111100110110" => rgb <= "000000";
					when "10111111100110111" => rgb <= "000000";
					when "10111111100111000" => rgb <= "000000";
					when "10111111100111001" => rgb <= "000000";
					when "10111111100111010" => rgb <= "000000";
					when "10111111100111011" => rgb <= "000000";
					when "10111111100111100" => rgb <= "000000";
					when "10111111100111101" => rgb <= "000000";
					when "10111111100111110" => rgb <= "000000";
					when "10111111100111111" => rgb <= "000000";
					when "11000000000000000" => rgb <= "000000";
					when "11000000000000001" => rgb <= "000000";
					when "11000000000000010" => rgb <= "000000";
					when "11000000000000011" => rgb <= "000000";
					when "11000000000000100" => rgb <= "000000";
					when "11000000000000101" => rgb <= "000000";
					when "11000000000000110" => rgb <= "000000";
					when "11000000000000111" => rgb <= "000000";
					when "11000000000001000" => rgb <= "000000";
					when "11000000000001001" => rgb <= "000000";
					when "11000000000001010" => rgb <= "000000";
					when "11000000000001011" => rgb <= "000000";
					when "11000000000001100" => rgb <= "000000";
					when "11000000000001101" => rgb <= "000000";
					when "11000000000001110" => rgb <= "000000";
					when "11000000000001111" => rgb <= "000000";
					when "11000000000010000" => rgb <= "000000";
					when "11000000000010001" => rgb <= "000000";
					when "11000000000010010" => rgb <= "000000";
					when "11000000000010011" => rgb <= "000000";
					when "11000000000010100" => rgb <= "101010";
					when "11000000000010101" => rgb <= "111111";
					when "11000000000010110" => rgb <= "101010";
					when "11000000000010111" => rgb <= "111111";
					when "11000000000011000" => rgb <= "111111";
					when "11000000000011001" => rgb <= "111111";
					when "11000000000011010" => rgb <= "111111";
					when "11000000000011011" => rgb <= "111111";
					when "11000000000011100" => rgb <= "111111";
					when "11000000000011101" => rgb <= "111111";
					when "11000000000011110" => rgb <= "111111";
					when "11000000000011111" => rgb <= "111111";
					when "11000000000100000" => rgb <= "111111";
					when "11000000000100001" => rgb <= "101010";
					when "11000000000100010" => rgb <= "101010";
					when "11000000000100011" => rgb <= "000000";
					when "11000000000100100" => rgb <= "000000";
					when "11000000000100101" => rgb <= "000000";
					when "11000000000100110" => rgb <= "000000";
					when "11000000000100111" => rgb <= "000000";
					when "11000000000101000" => rgb <= "000000";
					when "11000000000101001" => rgb <= "000000";
					when "11000000000101010" => rgb <= "000000";
					when "11000000000101011" => rgb <= "000000";
					when "11000000000101100" => rgb <= "000000";
					when "11000000000101101" => rgb <= "000000";
					when "11000000000101110" => rgb <= "000000";
					when "11000000000101111" => rgb <= "000000";
					when "11000000000110000" => rgb <= "000000";
					when "11000000000110001" => rgb <= "000000";
					when "11000000000110010" => rgb <= "000000";
					when "11000000000110011" => rgb <= "000000";
					when "11000000000110100" => rgb <= "000000";
					when "11000000000110101" => rgb <= "000000";
					when "11000000000110110" => rgb <= "000000";
					when "11000000000110111" => rgb <= "000000";
					when "11000000000111000" => rgb <= "000000";
					when "11000000000111001" => rgb <= "010101";
					when "11000000000111010" => rgb <= "101010";
					when "11000000000111011" => rgb <= "101010";
					when "11000000000111100" => rgb <= "101010";
					when "11000000000111101" => rgb <= "111111";
					when "11000000000111110" => rgb <= "111111";
					when "11000000000111111" => rgb <= "111111";
					when "11000000001000000" => rgb <= "101010";
					when "11000000001000001" => rgb <= "000000";
					when "11000000001000010" => rgb <= "000000";
					when "11000000001000011" => rgb <= "000000";
					when "11000000001000100" => rgb <= "000000";
					when "11000000001000101" => rgb <= "000000";
					when "11000000001000110" => rgb <= "000000";
					when "11000000001000111" => rgb <= "000000";
					when "11000000001001000" => rgb <= "000000";
					when "11000000001001001" => rgb <= "000000";
					when "11000000001001010" => rgb <= "000000";
					when "11000000001001011" => rgb <= "000000";
					when "11000000001001100" => rgb <= "000000";
					when "11000000001001101" => rgb <= "000000";
					when "11000000001001110" => rgb <= "000000";
					when "11000000001001111" => rgb <= "000000";
					when "11000000001010000" => rgb <= "101010";
					when "11000000001010001" => rgb <= "101010";
					when "11000000001010010" => rgb <= "101010";
					when "11000000001010011" => rgb <= "101010";
					when "11000000001010100" => rgb <= "111111";
					when "11000000001010101" => rgb <= "111111";
					when "11000000001010110" => rgb <= "101010";
					when "11000000001010111" => rgb <= "111111";
					when "11000000001011000" => rgb <= "111111";
					when "11000000001011001" => rgb <= "111111";
					when "11000000001011010" => rgb <= "111111";
					when "11000000001011011" => rgb <= "101010";
					when "11000000001011100" => rgb <= "111111";
					when "11000000001011101" => rgb <= "101010";
					when "11000000001011110" => rgb <= "101010";
					when "11000000001011111" => rgb <= "000000";
					when "11000000001100000" => rgb <= "000000";
					when "11000000001100001" => rgb <= "000000";
					when "11000000001100010" => rgb <= "000000";
					when "11000000001100011" => rgb <= "000000";
					when "11000000001100100" => rgb <= "000000";
					when "11000000001100101" => rgb <= "000000";
					when "11000000001100110" => rgb <= "010101";
					when "11000000001100111" => rgb <= "111111";
					when "11000000001101000" => rgb <= "101010";
					when "11000000001101001" => rgb <= "111111";
					when "11000000001101010" => rgb <= "101010";
					when "11000000001101011" => rgb <= "111111";
					when "11000000001101100" => rgb <= "101010";
					when "11000000001101101" => rgb <= "101010";
					when "11000000001101110" => rgb <= "000000";
					when "11000000001101111" => rgb <= "000000";
					when "11000000001110000" => rgb <= "000000";
					when "11000000001110001" => rgb <= "000000";
					when "11000000001110010" => rgb <= "000000";
					when "11000000001110011" => rgb <= "000000";
					when "11000000001110100" => rgb <= "000000";
					when "11000000001110101" => rgb <= "000000";
					when "11000000001110110" => rgb <= "000000";
					when "11000000001110111" => rgb <= "000000";
					when "11000000001111000" => rgb <= "000000";
					when "11000000001111001" => rgb <= "000000";
					when "11000000001111010" => rgb <= "000000";
					when "11000000001111011" => rgb <= "000000";
					when "11000000001111100" => rgb <= "000000";
					when "11000000001111101" => rgb <= "101010";
					when "11000000001111110" => rgb <= "111111";
					when "11000000001111111" => rgb <= "111111";
					when "11000000010000000" => rgb <= "111111";
					when "11000000010000001" => rgb <= "111111";
					when "11000000010000010" => rgb <= "111111";
					when "11000000010000011" => rgb <= "111111";
					when "11000000010000100" => rgb <= "111111";
					when "11000000010000101" => rgb <= "111111";
					when "11000000010000110" => rgb <= "111111";
					when "11000000010000111" => rgb <= "111111";
					when "11000000010001000" => rgb <= "111111";
					when "11000000010001001" => rgb <= "111111";
					when "11000000010001010" => rgb <= "111111";
					when "11000000010001011" => rgb <= "101010";
					when "11000000010001100" => rgb <= "000000";
					when "11000000010001101" => rgb <= "000000";
					when "11000000010001110" => rgb <= "000000";
					when "11000000010001111" => rgb <= "000000";
					when "11000000010010000" => rgb <= "000000";
					when "11000000010010001" => rgb <= "000000";
					when "11000000010010010" => rgb <= "000000";
					when "11000000010010011" => rgb <= "000000";
					when "11000000010010100" => rgb <= "000000";
					when "11000000010010101" => rgb <= "000000";
					when "11000000010010110" => rgb <= "000000";
					when "11000000010010111" => rgb <= "000000";
					when "11000000010011000" => rgb <= "000000";
					when "11000000010011001" => rgb <= "000000";
					when "11000000010011010" => rgb <= "000000";
					when "11000000010011011" => rgb <= "000000";
					when "11000000010011100" => rgb <= "000000";
					when "11000000010011101" => rgb <= "000000";
					when "11000000010011110" => rgb <= "000000";
					when "11000000010011111" => rgb <= "000000";
					when "11000000010100000" => rgb <= "000000";
					when "11000000010100001" => rgb <= "000000";
					when "11000000010100010" => rgb <= "010101";
					when "11000000010100011" => rgb <= "111111";
					when "11000000010100100" => rgb <= "101010";
					when "11000000010100101" => rgb <= "111111";
					when "11000000010100110" => rgb <= "111111";
					when "11000000010100111" => rgb <= "111111";
					when "11000000010101000" => rgb <= "111111";
					when "11000000010101001" => rgb <= "111111";
					when "11000000010101010" => rgb <= "000000";
					when "11000000010101011" => rgb <= "000000";
					when "11000000010101100" => rgb <= "000000";
					when "11000000010101101" => rgb <= "000000";
					when "11000000010101110" => rgb <= "000000";
					when "11000000010101111" => rgb <= "000000";
					when "11000000010110000" => rgb <= "000000";
					when "11000000010110001" => rgb <= "010101";
					when "11000000010110010" => rgb <= "101010";
					when "11000000010110011" => rgb <= "101010";
					when "11000000010110100" => rgb <= "111111";
					when "11000000010110101" => rgb <= "111111";
					when "11000000010110110" => rgb <= "101010";
					when "11000000010110111" => rgb <= "111111";
					when "11000000010111000" => rgb <= "101010";
					when "11000000010111001" => rgb <= "000000";
					when "11000000010111010" => rgb <= "000000";
					when "11000000010111011" => rgb <= "000000";
					when "11000000010111100" => rgb <= "000000";
					when "11000000010111101" => rgb <= "000000";
					when "11000000010111110" => rgb <= "000000";
					when "11000000010111111" => rgb <= "000000";
					when "11000000011000000" => rgb <= "010101";
					when "11000000011000001" => rgb <= "111111";
					when "11000000011000010" => rgb <= "101010";
					when "11000000011000011" => rgb <= "111111";
					when "11000000011000100" => rgb <= "101010";
					when "11000000011000101" => rgb <= "111111";
					when "11000000011000110" => rgb <= "111111";
					when "11000000011000111" => rgb <= "111111";
					when "11000000011001000" => rgb <= "111111";
					when "11000000011001001" => rgb <= "111111";
					when "11000000011001010" => rgb <= "111111";
					when "11000000011001011" => rgb <= "101010";
					when "11000000011001100" => rgb <= "111111";
					when "11000000011001101" => rgb <= "101010";
					when "11000000011001110" => rgb <= "111111";
					when "11000000011001111" => rgb <= "101010";
					when "11000000011010000" => rgb <= "000000";
					when "11000000011010001" => rgb <= "000000";
					when "11000000011010010" => rgb <= "000000";
					when "11000000011010011" => rgb <= "000000";
					when "11000000011010100" => rgb <= "000000";
					when "11000000011010101" => rgb <= "000000";
					when "11000000011010110" => rgb <= "000000";
					when "11000000011010111" => rgb <= "101010";
					when "11000000011011000" => rgb <= "101010";
					when "11000000011011001" => rgb <= "101010";
					when "11000000011011010" => rgb <= "101010";
					when "11000000011011011" => rgb <= "111111";
					when "11000000011011100" => rgb <= "111111";
					when "11000000011011101" => rgb <= "111111";
					when "11000000011011110" => rgb <= "111111";
					when "11000000011011111" => rgb <= "111111";
					when "11000000011100000" => rgb <= "111111";
					when "11000000011100001" => rgb <= "111111";
					when "11000000011100010" => rgb <= "111111";
					when "11000000011100011" => rgb <= "101010";
					when "11000000011100100" => rgb <= "111111";
					when "11000000011100101" => rgb <= "111111";
					when "11000000011100110" => rgb <= "000000";
					when "11000000011100111" => rgb <= "000000";
					when "11000000011101000" => rgb <= "000000";
					when "11000000011101001" => rgb <= "000000";
					when "11000000011101010" => rgb <= "000000";
					when "11000000011101011" => rgb <= "000000";
					when "11000000011101100" => rgb <= "000000";
					when "11000000011101101" => rgb <= "010101";
					when "11000000011101110" => rgb <= "111111";
					when "11000000011101111" => rgb <= "101010";
					when "11000000011110000" => rgb <= "111111";
					when "11000000011110001" => rgb <= "111111";
					when "11000000011110010" => rgb <= "111111";
					when "11000000011110011" => rgb <= "101010";
					when "11000000011110100" => rgb <= "101010";
					when "11000000011110101" => rgb <= "000000";
					when "11000000011110110" => rgb <= "000000";
					when "11000000011110111" => rgb <= "000000";
					when "11000000011111000" => rgb <= "000000";
					when "11000000011111001" => rgb <= "000000";
					when "11000000011111010" => rgb <= "000000";
					when "11000000011111011" => rgb <= "000000";
					when "11000000011111100" => rgb <= "000000";
					when "11000000011111101" => rgb <= "000000";
					when "11000000011111110" => rgb <= "000000";
					when "11000000011111111" => rgb <= "000000";
					when "11000000100000000" => rgb <= "000000";
					when "11000000100000001" => rgb <= "000000";
					when "11000000100000010" => rgb <= "000000";
					when "11000000100000011" => rgb <= "000000";
					when "11000000100000100" => rgb <= "000000";
					when "11000000100000101" => rgb <= "000000";
					when "11000000100000110" => rgb <= "000000";
					when "11000000100000111" => rgb <= "000000";
					when "11000000100001000" => rgb <= "000000";
					when "11000000100001001" => rgb <= "000000";
					when "11000000100001010" => rgb <= "000000";
					when "11000000100001011" => rgb <= "010101";
					when "11000000100001100" => rgb <= "111111";
					when "11000000100001101" => rgb <= "101010";
					when "11000000100001110" => rgb <= "111111";
					when "11000000100001111" => rgb <= "111111";
					when "11000000100010000" => rgb <= "111111";
					when "11000000100010001" => rgb <= "111111";
					when "11000000100010010" => rgb <= "111111";
					when "11000000100010011" => rgb <= "111111";
					when "11000000100010100" => rgb <= "111111";
					when "11000000100010101" => rgb <= "111111";
					when "11000000100010110" => rgb <= "111111";
					when "11000000100010111" => rgb <= "111111";
					when "11000000100011000" => rgb <= "101010";
					when "11000000100011001" => rgb <= "101010";
					when "11000000100011010" => rgb <= "101010";
					when "11000000100011011" => rgb <= "000000";
					when "11000000100011100" => rgb <= "000000";
					when "11000000100011101" => rgb <= "000000";
					when "11000000100011110" => rgb <= "000000";
					when "11000000100011111" => rgb <= "000000";
					when "11000000100100000" => rgb <= "000000";
					when "11000000100100001" => rgb <= "000000";
					when "11000000100100010" => rgb <= "101010";
					when "11000000100100011" => rgb <= "111111";
					when "11000000100100100" => rgb <= "111111";
					when "11000000100100101" => rgb <= "101010";
					when "11000000100100110" => rgb <= "111111";
					when "11000000100100111" => rgb <= "111111";
					when "11000000100101000" => rgb <= "101010";
					when "11000000100101001" => rgb <= "111111";
					when "11000000100101010" => rgb <= "111111";
					when "11000000100101011" => rgb <= "111111";
					when "11000000100101100" => rgb <= "111111";
					when "11000000100101101" => rgb <= "111111";
					when "11000000100101110" => rgb <= "111111";
					when "11000000100101111" => rgb <= "101010";
					when "11000000100110000" => rgb <= "111111";
					when "11000000100110001" => rgb <= "010101";
					when "11000000100110010" => rgb <= "000000";
					when "11000000100110011" => rgb <= "000000";
					when "11000000100110100" => rgb <= "000000";
					when "11000000100110101" => rgb <= "000000";
					when "11000000100110110" => rgb <= "000000";
					when "11000000100110111" => rgb <= "000000";
					when "11000000100111000" => rgb <= "000000";
					when "11000000100111001" => rgb <= "000000";
					when "11000000100111010" => rgb <= "000000";
					when "11000000100111011" => rgb <= "000000";
					when "11000000100111100" => rgb <= "000000";
					when "11000000100111101" => rgb <= "000000";
					when "11000000100111110" => rgb <= "000000";
					when "11000000100111111" => rgb <= "000000";
					when "11000001000000000" => rgb <= "000000";
					when "11000001000000001" => rgb <= "000000";
					when "11000001000000010" => rgb <= "000000";
					when "11000001000000011" => rgb <= "000000";
					when "11000001000000100" => rgb <= "000000";
					when "11000001000000101" => rgb <= "000000";
					when "11000001000000110" => rgb <= "000000";
					when "11000001000000111" => rgb <= "000000";
					when "11000001000001000" => rgb <= "000000";
					when "11000001000001001" => rgb <= "000000";
					when "11000001000001010" => rgb <= "000000";
					when "11000001000001011" => rgb <= "000000";
					when "11000001000001100" => rgb <= "000000";
					when "11000001000001101" => rgb <= "000000";
					when "11000001000001110" => rgb <= "000000";
					when "11000001000001111" => rgb <= "000000";
					when "11000001000010000" => rgb <= "000000";
					when "11000001000010001" => rgb <= "000000";
					when "11000001000010010" => rgb <= "000000";
					when "11000001000010011" => rgb <= "000000";
					when "11000001000010100" => rgb <= "101010";
					when "11000001000010101" => rgb <= "111111";
					when "11000001000010110" => rgb <= "101010";
					when "11000001000010111" => rgb <= "111111";
					when "11000001000011000" => rgb <= "111111";
					when "11000001000011001" => rgb <= "111111";
					when "11000001000011010" => rgb <= "111111";
					when "11000001000011011" => rgb <= "111111";
					when "11000001000011100" => rgb <= "111111";
					when "11000001000011101" => rgb <= "111111";
					when "11000001000011110" => rgb <= "111111";
					when "11000001000011111" => rgb <= "111111";
					when "11000001000100000" => rgb <= "111111";
					when "11000001000100001" => rgb <= "111111";
					when "11000001000100010" => rgb <= "111111";
					when "11000001000100011" => rgb <= "000000";
					when "11000001000100100" => rgb <= "000000";
					when "11000001000100101" => rgb <= "000000";
					when "11000001000100110" => rgb <= "000000";
					when "11000001000100111" => rgb <= "000000";
					when "11000001000101000" => rgb <= "000000";
					when "11000001000101001" => rgb <= "000000";
					when "11000001000101010" => rgb <= "000000";
					when "11000001000101011" => rgb <= "000000";
					when "11000001000101100" => rgb <= "000000";
					when "11000001000101101" => rgb <= "000000";
					when "11000001000101110" => rgb <= "000000";
					when "11000001000101111" => rgb <= "000000";
					when "11000001000110000" => rgb <= "000000";
					when "11000001000110001" => rgb <= "000000";
					when "11000001000110010" => rgb <= "000000";
					when "11000001000110011" => rgb <= "000000";
					when "11000001000110100" => rgb <= "000000";
					when "11000001000110101" => rgb <= "000000";
					when "11000001000110110" => rgb <= "000000";
					when "11000001000110111" => rgb <= "000000";
					when "11000001000111000" => rgb <= "000000";
					when "11000001000111001" => rgb <= "010101";
					when "11000001000111010" => rgb <= "101010";
					when "11000001000111011" => rgb <= "101010";
					when "11000001000111100" => rgb <= "101010";
					when "11000001000111101" => rgb <= "111111";
					when "11000001000111110" => rgb <= "111111";
					when "11000001000111111" => rgb <= "111111";
					when "11000001001000000" => rgb <= "101010";
					when "11000001001000001" => rgb <= "000000";
					when "11000001001000010" => rgb <= "000000";
					when "11000001001000011" => rgb <= "000000";
					when "11000001001000100" => rgb <= "000000";
					when "11000001001000101" => rgb <= "000000";
					when "11000001001000110" => rgb <= "000000";
					when "11000001001000111" => rgb <= "000000";
					when "11000001001001000" => rgb <= "000000";
					when "11000001001001001" => rgb <= "000000";
					when "11000001001001010" => rgb <= "000000";
					when "11000001001001011" => rgb <= "000000";
					when "11000001001001100" => rgb <= "000000";
					when "11000001001001101" => rgb <= "000000";
					when "11000001001001110" => rgb <= "000000";
					when "11000001001001111" => rgb <= "000000";
					when "11000001001010000" => rgb <= "101010";
					when "11000001001010001" => rgb <= "101010";
					when "11000001001010010" => rgb <= "101010";
					when "11000001001010011" => rgb <= "101010";
					when "11000001001010100" => rgb <= "111111";
					when "11000001001010101" => rgb <= "111111";
					when "11000001001010110" => rgb <= "101010";
					when "11000001001010111" => rgb <= "111111";
					when "11000001001011000" => rgb <= "111111";
					when "11000001001011001" => rgb <= "111111";
					when "11000001001011010" => rgb <= "111111";
					when "11000001001011011" => rgb <= "101010";
					when "11000001001011100" => rgb <= "111111";
					when "11000001001011101" => rgb <= "101010";
					when "11000001001011110" => rgb <= "101010";
					when "11000001001011111" => rgb <= "000000";
					when "11000001001100000" => rgb <= "000000";
					when "11000001001100001" => rgb <= "000000";
					when "11000001001100010" => rgb <= "000000";
					when "11000001001100011" => rgb <= "000000";
					when "11000001001100100" => rgb <= "000000";
					when "11000001001100101" => rgb <= "000000";
					when "11000001001100110" => rgb <= "010101";
					when "11000001001100111" => rgb <= "111111";
					when "11000001001101000" => rgb <= "101010";
					when "11000001001101001" => rgb <= "111111";
					when "11000001001101010" => rgb <= "101010";
					when "11000001001101011" => rgb <= "111111";
					when "11000001001101100" => rgb <= "101010";
					when "11000001001101101" => rgb <= "101010";
					when "11000001001101110" => rgb <= "000000";
					when "11000001001101111" => rgb <= "000000";
					when "11000001001110000" => rgb <= "000000";
					when "11000001001110001" => rgb <= "000000";
					when "11000001001110010" => rgb <= "000000";
					when "11000001001110011" => rgb <= "000000";
					when "11000001001110100" => rgb <= "000000";
					when "11000001001110101" => rgb <= "000000";
					when "11000001001110110" => rgb <= "000000";
					when "11000001001110111" => rgb <= "000000";
					when "11000001001111000" => rgb <= "000000";
					when "11000001001111001" => rgb <= "000000";
					when "11000001001111010" => rgb <= "000000";
					when "11000001001111011" => rgb <= "000000";
					when "11000001001111100" => rgb <= "000000";
					when "11000001001111101" => rgb <= "101010";
					when "11000001001111110" => rgb <= "111111";
					when "11000001001111111" => rgb <= "111111";
					when "11000001010000000" => rgb <= "111111";
					when "11000001010000001" => rgb <= "111111";
					when "11000001010000010" => rgb <= "111111";
					when "11000001010000011" => rgb <= "111111";
					when "11000001010000100" => rgb <= "111111";
					when "11000001010000101" => rgb <= "111111";
					when "11000001010000110" => rgb <= "111111";
					when "11000001010000111" => rgb <= "111111";
					when "11000001010001000" => rgb <= "111111";
					when "11000001010001001" => rgb <= "111111";
					when "11000001010001010" => rgb <= "111111";
					when "11000001010001011" => rgb <= "101010";
					when "11000001010001100" => rgb <= "000000";
					when "11000001010001101" => rgb <= "000000";
					when "11000001010001110" => rgb <= "000000";
					when "11000001010001111" => rgb <= "000000";
					when "11000001010010000" => rgb <= "000000";
					when "11000001010010001" => rgb <= "000000";
					when "11000001010010010" => rgb <= "000000";
					when "11000001010010011" => rgb <= "000000";
					when "11000001010010100" => rgb <= "000000";
					when "11000001010010101" => rgb <= "000000";
					when "11000001010010110" => rgb <= "000000";
					when "11000001010010111" => rgb <= "000000";
					when "11000001010011000" => rgb <= "000000";
					when "11000001010011001" => rgb <= "000000";
					when "11000001010011010" => rgb <= "000000";
					when "11000001010011011" => rgb <= "000000";
					when "11000001010011100" => rgb <= "000000";
					when "11000001010011101" => rgb <= "000000";
					when "11000001010011110" => rgb <= "000000";
					when "11000001010011111" => rgb <= "000000";
					when "11000001010100000" => rgb <= "000000";
					when "11000001010100001" => rgb <= "000000";
					when "11000001010100010" => rgb <= "010101";
					when "11000001010100011" => rgb <= "111111";
					when "11000001010100100" => rgb <= "101010";
					when "11000001010100101" => rgb <= "111111";
					when "11000001010100110" => rgb <= "111111";
					when "11000001010100111" => rgb <= "111111";
					when "11000001010101000" => rgb <= "111111";
					when "11000001010101001" => rgb <= "111111";
					when "11000001010101010" => rgb <= "000000";
					when "11000001010101011" => rgb <= "000000";
					when "11000001010101100" => rgb <= "000000";
					when "11000001010101101" => rgb <= "000000";
					when "11000001010101110" => rgb <= "000000";
					when "11000001010101111" => rgb <= "000000";
					when "11000001010110000" => rgb <= "000000";
					when "11000001010110001" => rgb <= "010101";
					when "11000001010110010" => rgb <= "101010";
					when "11000001010110011" => rgb <= "101010";
					when "11000001010110100" => rgb <= "111111";
					when "11000001010110101" => rgb <= "111111";
					when "11000001010110110" => rgb <= "101010";
					when "11000001010110111" => rgb <= "111111";
					when "11000001010111000" => rgb <= "101010";
					when "11000001010111001" => rgb <= "000000";
					when "11000001010111010" => rgb <= "000000";
					when "11000001010111011" => rgb <= "000000";
					when "11000001010111100" => rgb <= "000000";
					when "11000001010111101" => rgb <= "000000";
					when "11000001010111110" => rgb <= "000000";
					when "11000001010111111" => rgb <= "000000";
					when "11000001011000000" => rgb <= "010101";
					when "11000001011000001" => rgb <= "111111";
					when "11000001011000010" => rgb <= "101010";
					when "11000001011000011" => rgb <= "111111";
					when "11000001011000100" => rgb <= "101010";
					when "11000001011000101" => rgb <= "111111";
					when "11000001011000110" => rgb <= "111111";
					when "11000001011000111" => rgb <= "111111";
					when "11000001011001000" => rgb <= "111111";
					when "11000001011001001" => rgb <= "111111";
					when "11000001011001010" => rgb <= "111111";
					when "11000001011001011" => rgb <= "101010";
					when "11000001011001100" => rgb <= "111111";
					when "11000001011001101" => rgb <= "101010";
					when "11000001011001110" => rgb <= "111111";
					when "11000001011001111" => rgb <= "101010";
					when "11000001011010000" => rgb <= "000000";
					when "11000001011010001" => rgb <= "000000";
					when "11000001011010010" => rgb <= "000000";
					when "11000001011010011" => rgb <= "000000";
					when "11000001011010100" => rgb <= "000000";
					when "11000001011010101" => rgb <= "000000";
					when "11000001011010110" => rgb <= "000000";
					when "11000001011010111" => rgb <= "101010";
					when "11000001011011000" => rgb <= "101010";
					when "11000001011011001" => rgb <= "101010";
					when "11000001011011010" => rgb <= "101010";
					when "11000001011011011" => rgb <= "111111";
					when "11000001011011100" => rgb <= "111111";
					when "11000001011011101" => rgb <= "111111";
					when "11000001011011110" => rgb <= "111111";
					when "11000001011011111" => rgb <= "111111";
					when "11000001011100000" => rgb <= "111111";
					when "11000001011100001" => rgb <= "111111";
					when "11000001011100010" => rgb <= "111111";
					when "11000001011100011" => rgb <= "101010";
					when "11000001011100100" => rgb <= "111111";
					when "11000001011100101" => rgb <= "111111";
					when "11000001011100110" => rgb <= "000000";
					when "11000001011100111" => rgb <= "000000";
					when "11000001011101000" => rgb <= "000000";
					when "11000001011101001" => rgb <= "000000";
					when "11000001011101010" => rgb <= "000000";
					when "11000001011101011" => rgb <= "000000";
					when "11000001011101100" => rgb <= "000000";
					when "11000001011101101" => rgb <= "010101";
					when "11000001011101110" => rgb <= "111111";
					when "11000001011101111" => rgb <= "101010";
					when "11000001011110000" => rgb <= "111111";
					when "11000001011110001" => rgb <= "111111";
					when "11000001011110010" => rgb <= "111111";
					when "11000001011110011" => rgb <= "101010";
					when "11000001011110100" => rgb <= "101010";
					when "11000001011110101" => rgb <= "000000";
					when "11000001011110110" => rgb <= "000000";
					when "11000001011110111" => rgb <= "000000";
					when "11000001011111000" => rgb <= "000000";
					when "11000001011111001" => rgb <= "000000";
					when "11000001011111010" => rgb <= "000000";
					when "11000001011111011" => rgb <= "000000";
					when "11000001011111100" => rgb <= "000000";
					when "11000001011111101" => rgb <= "000000";
					when "11000001011111110" => rgb <= "000000";
					when "11000001011111111" => rgb <= "000000";
					when "11000001100000000" => rgb <= "000000";
					when "11000001100000001" => rgb <= "000000";
					when "11000001100000010" => rgb <= "000000";
					when "11000001100000011" => rgb <= "000000";
					when "11000001100000100" => rgb <= "000000";
					when "11000001100000101" => rgb <= "000000";
					when "11000001100000110" => rgb <= "000000";
					when "11000001100000111" => rgb <= "000000";
					when "11000001100001000" => rgb <= "000000";
					when "11000001100001001" => rgb <= "000000";
					when "11000001100001010" => rgb <= "000000";
					when "11000001100001011" => rgb <= "010101";
					when "11000001100001100" => rgb <= "111111";
					when "11000001100001101" => rgb <= "101010";
					when "11000001100001110" => rgb <= "111111";
					when "11000001100001111" => rgb <= "111111";
					when "11000001100010000" => rgb <= "111111";
					when "11000001100010001" => rgb <= "111111";
					when "11000001100010010" => rgb <= "111111";
					when "11000001100010011" => rgb <= "111111";
					when "11000001100010100" => rgb <= "111111";
					when "11000001100010101" => rgb <= "111111";
					when "11000001100010110" => rgb <= "111111";
					when "11000001100010111" => rgb <= "111111";
					when "11000001100011000" => rgb <= "101010";
					when "11000001100011001" => rgb <= "101010";
					when "11000001100011010" => rgb <= "101010";
					when "11000001100011011" => rgb <= "000000";
					when "11000001100011100" => rgb <= "000000";
					when "11000001100011101" => rgb <= "000000";
					when "11000001100011110" => rgb <= "000000";
					when "11000001100011111" => rgb <= "000000";
					when "11000001100100000" => rgb <= "000000";
					when "11000001100100001" => rgb <= "000000";
					when "11000001100100010" => rgb <= "101010";
					when "11000001100100011" => rgb <= "111111";
					when "11000001100100100" => rgb <= "101010";
					when "11000001100100101" => rgb <= "111111";
					when "11000001100100110" => rgb <= "101010";
					when "11000001100100111" => rgb <= "111111";
					when "11000001100101000" => rgb <= "111111";
					when "11000001100101001" => rgb <= "111111";
					when "11000001100101010" => rgb <= "111111";
					when "11000001100101011" => rgb <= "111111";
					when "11000001100101100" => rgb <= "111111";
					when "11000001100101101" => rgb <= "111111";
					when "11000001100101110" => rgb <= "101010";
					when "11000001100101111" => rgb <= "101010";
					when "11000001100110000" => rgb <= "111111";
					when "11000001100110001" => rgb <= "010101";
					when "11000001100110010" => rgb <= "000000";
					when "11000001100110011" => rgb <= "000000";
					when "11000001100110100" => rgb <= "000000";
					when "11000001100110101" => rgb <= "000000";
					when "11000001100110110" => rgb <= "000000";
					when "11000001100110111" => rgb <= "000000";
					when "11000001100111000" => rgb <= "000000";
					when "11000001100111001" => rgb <= "000000";
					when "11000001100111010" => rgb <= "000000";
					when "11000001100111011" => rgb <= "000000";
					when "11000001100111100" => rgb <= "000000";
					when "11000001100111101" => rgb <= "000000";
					when "11000001100111110" => rgb <= "000000";
					when "11000001100111111" => rgb <= "000000";
					when "11000010000000000" => rgb <= "000000";
					when "11000010000000001" => rgb <= "000000";
					when "11000010000000010" => rgb <= "000000";
					when "11000010000000011" => rgb <= "000000";
					when "11000010000000100" => rgb <= "000000";
					when "11000010000000101" => rgb <= "000000";
					when "11000010000000110" => rgb <= "000000";
					when "11000010000000111" => rgb <= "000000";
					when "11000010000001000" => rgb <= "000000";
					when "11000010000001001" => rgb <= "000000";
					when "11000010000001010" => rgb <= "000000";
					when "11000010000001011" => rgb <= "000000";
					when "11000010000001100" => rgb <= "000000";
					when "11000010000001101" => rgb <= "000000";
					when "11000010000001110" => rgb <= "000000";
					when "11000010000001111" => rgb <= "000000";
					when "11000010000010000" => rgb <= "000000";
					when "11000010000010001" => rgb <= "000000";
					when "11000010000010010" => rgb <= "000000";
					when "11000010000010011" => rgb <= "000000";
					when "11000010000010100" => rgb <= "101010";
					when "11000010000010101" => rgb <= "111111";
					when "11000010000010110" => rgb <= "101010";
					when "11000010000010111" => rgb <= "111111";
					when "11000010000011000" => rgb <= "111111";
					when "11000010000011001" => rgb <= "111111";
					when "11000010000011010" => rgb <= "111111";
					when "11000010000011011" => rgb <= "111111";
					when "11000010000011100" => rgb <= "111111";
					when "11000010000011101" => rgb <= "111111";
					when "11000010000011110" => rgb <= "111111";
					when "11000010000011111" => rgb <= "111111";
					when "11000010000100000" => rgb <= "111111";
					when "11000010000100001" => rgb <= "101010";
					when "11000010000100010" => rgb <= "111111";
					when "11000010000100011" => rgb <= "000000";
					when "11000010000100100" => rgb <= "000000";
					when "11000010000100101" => rgb <= "000000";
					when "11000010000100110" => rgb <= "000000";
					when "11000010000100111" => rgb <= "000000";
					when "11000010000101000" => rgb <= "000000";
					when "11000010000101001" => rgb <= "000000";
					when "11000010000101010" => rgb <= "000000";
					when "11000010000101011" => rgb <= "000000";
					when "11000010000101100" => rgb <= "000000";
					when "11000010000101101" => rgb <= "000000";
					when "11000010000101110" => rgb <= "000000";
					when "11000010000101111" => rgb <= "000000";
					when "11000010000110000" => rgb <= "000000";
					when "11000010000110001" => rgb <= "000000";
					when "11000010000110010" => rgb <= "000000";
					when "11000010000110011" => rgb <= "000000";
					when "11000010000110100" => rgb <= "000000";
					when "11000010000110101" => rgb <= "000000";
					when "11000010000110110" => rgb <= "000000";
					when "11000010000110111" => rgb <= "000000";
					when "11000010000111000" => rgb <= "000000";
					when "11000010000111001" => rgb <= "010101";
					when "11000010000111010" => rgb <= "101010";
					when "11000010000111011" => rgb <= "101010";
					when "11000010000111100" => rgb <= "101010";
					when "11000010000111101" => rgb <= "111111";
					when "11000010000111110" => rgb <= "111111";
					when "11000010000111111" => rgb <= "111111";
					when "11000010001000000" => rgb <= "101010";
					when "11000010001000001" => rgb <= "000000";
					when "11000010001000010" => rgb <= "000000";
					when "11000010001000011" => rgb <= "000000";
					when "11000010001000100" => rgb <= "000000";
					when "11000010001000101" => rgb <= "000000";
					when "11000010001000110" => rgb <= "000000";
					when "11000010001000111" => rgb <= "000000";
					when "11000010001001000" => rgb <= "000000";
					when "11000010001001001" => rgb <= "000000";
					when "11000010001001010" => rgb <= "000000";
					when "11000010001001011" => rgb <= "000000";
					when "11000010001001100" => rgb <= "000000";
					when "11000010001001101" => rgb <= "000000";
					when "11000010001001110" => rgb <= "000000";
					when "11000010001001111" => rgb <= "000000";
					when "11000010001010000" => rgb <= "101010";
					when "11000010001010001" => rgb <= "101010";
					when "11000010001010010" => rgb <= "101010";
					when "11000010001010011" => rgb <= "101010";
					when "11000010001010100" => rgb <= "111111";
					when "11000010001010101" => rgb <= "111111";
					when "11000010001010110" => rgb <= "101010";
					when "11000010001010111" => rgb <= "111111";
					when "11000010001011000" => rgb <= "111111";
					when "11000010001011001" => rgb <= "111111";
					when "11000010001011010" => rgb <= "111111";
					when "11000010001011011" => rgb <= "101010";
					when "11000010001011100" => rgb <= "111111";
					when "11000010001011101" => rgb <= "101010";
					when "11000010001011110" => rgb <= "101010";
					when "11000010001011111" => rgb <= "000000";
					when "11000010001100000" => rgb <= "000000";
					when "11000010001100001" => rgb <= "000000";
					when "11000010001100010" => rgb <= "000000";
					when "11000010001100011" => rgb <= "000000";
					when "11000010001100100" => rgb <= "000000";
					when "11000010001100101" => rgb <= "000000";
					when "11000010001100110" => rgb <= "010101";
					when "11000010001100111" => rgb <= "111111";
					when "11000010001101000" => rgb <= "101010";
					when "11000010001101001" => rgb <= "111111";
					when "11000010001101010" => rgb <= "101010";
					when "11000010001101011" => rgb <= "111111";
					when "11000010001101100" => rgb <= "101010";
					when "11000010001101101" => rgb <= "101010";
					when "11000010001101110" => rgb <= "000000";
					when "11000010001101111" => rgb <= "000000";
					when "11000010001110000" => rgb <= "000000";
					when "11000010001110001" => rgb <= "000000";
					when "11000010001110010" => rgb <= "000000";
					when "11000010001110011" => rgb <= "000000";
					when "11000010001110100" => rgb <= "000000";
					when "11000010001110101" => rgb <= "000000";
					when "11000010001110110" => rgb <= "000000";
					when "11000010001110111" => rgb <= "000000";
					when "11000010001111000" => rgb <= "000000";
					when "11000010001111001" => rgb <= "000000";
					when "11000010001111010" => rgb <= "000000";
					when "11000010001111011" => rgb <= "000000";
					when "11000010001111100" => rgb <= "000000";
					when "11000010001111101" => rgb <= "101010";
					when "11000010001111110" => rgb <= "111111";
					when "11000010001111111" => rgb <= "111111";
					when "11000010010000000" => rgb <= "111111";
					when "11000010010000001" => rgb <= "111111";
					when "11000010010000010" => rgb <= "111111";
					when "11000010010000011" => rgb <= "111111";
					when "11000010010000100" => rgb <= "111111";
					when "11000010010000101" => rgb <= "111111";
					when "11000010010000110" => rgb <= "111111";
					when "11000010010000111" => rgb <= "111111";
					when "11000010010001000" => rgb <= "111111";
					when "11000010010001001" => rgb <= "111111";
					when "11000010010001010" => rgb <= "111111";
					when "11000010010001011" => rgb <= "101010";
					when "11000010010001100" => rgb <= "000000";
					when "11000010010001101" => rgb <= "000000";
					when "11000010010001110" => rgb <= "000000";
					when "11000010010001111" => rgb <= "000000";
					when "11000010010010000" => rgb <= "000000";
					when "11000010010010001" => rgb <= "000000";
					when "11000010010010010" => rgb <= "000000";
					when "11000010010010011" => rgb <= "000000";
					when "11000010010010100" => rgb <= "000000";
					when "11000010010010101" => rgb <= "000000";
					when "11000010010010110" => rgb <= "000000";
					when "11000010010010111" => rgb <= "000000";
					when "11000010010011000" => rgb <= "000000";
					when "11000010010011001" => rgb <= "000000";
					when "11000010010011010" => rgb <= "000000";
					when "11000010010011011" => rgb <= "000000";
					when "11000010010011100" => rgb <= "000000";
					when "11000010010011101" => rgb <= "000000";
					when "11000010010011110" => rgb <= "000000";
					when "11000010010011111" => rgb <= "000000";
					when "11000010010100000" => rgb <= "000000";
					when "11000010010100001" => rgb <= "000000";
					when "11000010010100010" => rgb <= "010101";
					when "11000010010100011" => rgb <= "111111";
					when "11000010010100100" => rgb <= "101010";
					when "11000010010100101" => rgb <= "111111";
					when "11000010010100110" => rgb <= "111111";
					when "11000010010100111" => rgb <= "111111";
					when "11000010010101000" => rgb <= "111111";
					when "11000010010101001" => rgb <= "111111";
					when "11000010010101010" => rgb <= "000000";
					when "11000010010101011" => rgb <= "000000";
					when "11000010010101100" => rgb <= "000000";
					when "11000010010101101" => rgb <= "000000";
					when "11000010010101110" => rgb <= "000000";
					when "11000010010101111" => rgb <= "000000";
					when "11000010010110000" => rgb <= "000000";
					when "11000010010110001" => rgb <= "010101";
					when "11000010010110010" => rgb <= "101010";
					when "11000010010110011" => rgb <= "101010";
					when "11000010010110100" => rgb <= "111111";
					when "11000010010110101" => rgb <= "111111";
					when "11000010010110110" => rgb <= "101010";
					when "11000010010110111" => rgb <= "111111";
					when "11000010010111000" => rgb <= "101010";
					when "11000010010111001" => rgb <= "000000";
					when "11000010010111010" => rgb <= "000000";
					when "11000010010111011" => rgb <= "000000";
					when "11000010010111100" => rgb <= "000000";
					when "11000010010111101" => rgb <= "000000";
					when "11000010010111110" => rgb <= "000000";
					when "11000010010111111" => rgb <= "000000";
					when "11000010011000000" => rgb <= "010101";
					when "11000010011000001" => rgb <= "111111";
					when "11000010011000010" => rgb <= "101010";
					when "11000010011000011" => rgb <= "111111";
					when "11000010011000100" => rgb <= "101010";
					when "11000010011000101" => rgb <= "111111";
					when "11000010011000110" => rgb <= "111111";
					when "11000010011000111" => rgb <= "111111";
					when "11000010011001000" => rgb <= "111111";
					when "11000010011001001" => rgb <= "111111";
					when "11000010011001010" => rgb <= "111111";
					when "11000010011001011" => rgb <= "101010";
					when "11000010011001100" => rgb <= "111111";
					when "11000010011001101" => rgb <= "101010";
					when "11000010011001110" => rgb <= "111111";
					when "11000010011001111" => rgb <= "101010";
					when "11000010011010000" => rgb <= "000000";
					when "11000010011010001" => rgb <= "000000";
					when "11000010011010010" => rgb <= "000000";
					when "11000010011010011" => rgb <= "000000";
					when "11000010011010100" => rgb <= "000000";
					when "11000010011010101" => rgb <= "000000";
					when "11000010011010110" => rgb <= "000000";
					when "11000010011010111" => rgb <= "101010";
					when "11000010011011000" => rgb <= "101010";
					when "11000010011011001" => rgb <= "101010";
					when "11000010011011010" => rgb <= "101010";
					when "11000010011011011" => rgb <= "111111";
					when "11000010011011100" => rgb <= "111111";
					when "11000010011011101" => rgb <= "111111";
					when "11000010011011110" => rgb <= "111111";
					when "11000010011011111" => rgb <= "111111";
					when "11000010011100000" => rgb <= "111111";
					when "11000010011100001" => rgb <= "111111";
					when "11000010011100010" => rgb <= "111111";
					when "11000010011100011" => rgb <= "101010";
					when "11000010011100100" => rgb <= "111111";
					when "11000010011100101" => rgb <= "111111";
					when "11000010011100110" => rgb <= "000000";
					when "11000010011100111" => rgb <= "000000";
					when "11000010011101000" => rgb <= "000000";
					when "11000010011101001" => rgb <= "000000";
					when "11000010011101010" => rgb <= "000000";
					when "11000010011101011" => rgb <= "000000";
					when "11000010011101100" => rgb <= "000000";
					when "11000010011101101" => rgb <= "010101";
					when "11000010011101110" => rgb <= "111111";
					when "11000010011101111" => rgb <= "101010";
					when "11000010011110000" => rgb <= "111111";
					when "11000010011110001" => rgb <= "111111";
					when "11000010011110010" => rgb <= "111111";
					when "11000010011110011" => rgb <= "101010";
					when "11000010011110100" => rgb <= "101010";
					when "11000010011110101" => rgb <= "000000";
					when "11000010011110110" => rgb <= "000000";
					when "11000010011110111" => rgb <= "000000";
					when "11000010011111000" => rgb <= "000000";
					when "11000010011111001" => rgb <= "000000";
					when "11000010011111010" => rgb <= "000000";
					when "11000010011111011" => rgb <= "000000";
					when "11000010011111100" => rgb <= "000000";
					when "11000010011111101" => rgb <= "000000";
					when "11000010011111110" => rgb <= "000000";
					when "11000010011111111" => rgb <= "000000";
					when "11000010100000000" => rgb <= "000000";
					when "11000010100000001" => rgb <= "000000";
					when "11000010100000010" => rgb <= "000000";
					when "11000010100000011" => rgb <= "000000";
					when "11000010100000100" => rgb <= "000000";
					when "11000010100000101" => rgb <= "000000";
					when "11000010100000110" => rgb <= "000000";
					when "11000010100000111" => rgb <= "000000";
					when "11000010100001000" => rgb <= "000000";
					when "11000010100001001" => rgb <= "000000";
					when "11000010100001010" => rgb <= "000000";
					when "11000010100001011" => rgb <= "010101";
					when "11000010100001100" => rgb <= "111111";
					when "11000010100001101" => rgb <= "101010";
					when "11000010100001110" => rgb <= "111111";
					when "11000010100001111" => rgb <= "111111";
					when "11000010100010000" => rgb <= "111111";
					when "11000010100010001" => rgb <= "111111";
					when "11000010100010010" => rgb <= "111111";
					when "11000010100010011" => rgb <= "111111";
					when "11000010100010100" => rgb <= "111111";
					when "11000010100010101" => rgb <= "111111";
					when "11000010100010110" => rgb <= "111111";
					when "11000010100010111" => rgb <= "111111";
					when "11000010100011000" => rgb <= "101010";
					when "11000010100011001" => rgb <= "101010";
					when "11000010100011010" => rgb <= "101010";
					when "11000010100011011" => rgb <= "000000";
					when "11000010100011100" => rgb <= "000000";
					when "11000010100011101" => rgb <= "000000";
					when "11000010100011110" => rgb <= "000000";
					when "11000010100011111" => rgb <= "000000";
					when "11000010100100000" => rgb <= "000000";
					when "11000010100100001" => rgb <= "000000";
					when "11000010100100010" => rgb <= "101010";
					when "11000010100100011" => rgb <= "101010";
					when "11000010100100100" => rgb <= "101010";
					when "11000010100100101" => rgb <= "111111";
					when "11000010100100110" => rgb <= "101010";
					when "11000010100100111" => rgb <= "111111";
					when "11000010100101000" => rgb <= "111111";
					when "11000010100101001" => rgb <= "111111";
					when "11000010100101010" => rgb <= "111111";
					when "11000010100101011" => rgb <= "111111";
					when "11000010100101100" => rgb <= "111111";
					when "11000010100101101" => rgb <= "111111";
					when "11000010100101110" => rgb <= "111111";
					when "11000010100101111" => rgb <= "101010";
					when "11000010100110000" => rgb <= "111111";
					when "11000010100110001" => rgb <= "010101";
					when "11000010100110010" => rgb <= "000000";
					when "11000010100110011" => rgb <= "000000";
					when "11000010100110100" => rgb <= "000000";
					when "11000010100110101" => rgb <= "000000";
					when "11000010100110110" => rgb <= "000000";
					when "11000010100110111" => rgb <= "000000";
					when "11000010100111000" => rgb <= "000000";
					when "11000010100111001" => rgb <= "000000";
					when "11000010100111010" => rgb <= "000000";
					when "11000010100111011" => rgb <= "000000";
					when "11000010100111100" => rgb <= "000000";
					when "11000010100111101" => rgb <= "000000";
					when "11000010100111110" => rgb <= "000000";
					when "11000010100111111" => rgb <= "000000";
					when "11000011000000000" => rgb <= "000000";
					when "11000011000000001" => rgb <= "000000";
					when "11000011000000010" => rgb <= "000000";
					when "11000011000000011" => rgb <= "000000";
					when "11000011000000100" => rgb <= "000000";
					when "11000011000000101" => rgb <= "000000";
					when "11000011000000110" => rgb <= "000000";
					when "11000011000000111" => rgb <= "000000";
					when "11000011000001000" => rgb <= "000000";
					when "11000011000001001" => rgb <= "000000";
					when "11000011000001010" => rgb <= "000000";
					when "11000011000001011" => rgb <= "000000";
					when "11000011000001100" => rgb <= "000000";
					when "11000011000001101" => rgb <= "000000";
					when "11000011000001110" => rgb <= "000000";
					when "11000011000001111" => rgb <= "000000";
					when "11000011000010000" => rgb <= "000000";
					when "11000011000010001" => rgb <= "000000";
					when "11000011000010010" => rgb <= "000000";
					when "11000011000010011" => rgb <= "000000";
					when "11000011000010100" => rgb <= "101010";
					when "11000011000010101" => rgb <= "111111";
					when "11000011000010110" => rgb <= "101010";
					when "11000011000010111" => rgb <= "111111";
					when "11000011000011000" => rgb <= "111111";
					when "11000011000011001" => rgb <= "111111";
					when "11000011000011010" => rgb <= "111111";
					when "11000011000011011" => rgb <= "111111";
					when "11000011000011100" => rgb <= "111111";
					when "11000011000011101" => rgb <= "111111";
					when "11000011000011110" => rgb <= "111111";
					when "11000011000011111" => rgb <= "111111";
					when "11000011000100000" => rgb <= "111111";
					when "11000011000100001" => rgb <= "101010";
					when "11000011000100010" => rgb <= "101010";
					when "11000011000100011" => rgb <= "000000";
					when "11000011000100100" => rgb <= "000000";
					when "11000011000100101" => rgb <= "000000";
					when "11000011000100110" => rgb <= "000000";
					when "11000011000100111" => rgb <= "000000";
					when "11000011000101000" => rgb <= "000000";
					when "11000011000101001" => rgb <= "000000";
					when "11000011000101010" => rgb <= "000000";
					when "11000011000101011" => rgb <= "000000";
					when "11000011000101100" => rgb <= "000000";
					when "11000011000101101" => rgb <= "000000";
					when "11000011000101110" => rgb <= "000000";
					when "11000011000101111" => rgb <= "000000";
					when "11000011000110000" => rgb <= "000000";
					when "11000011000110001" => rgb <= "000000";
					when "11000011000110010" => rgb <= "000000";
					when "11000011000110011" => rgb <= "000000";
					when "11000011000110100" => rgb <= "000000";
					when "11000011000110101" => rgb <= "000000";
					when "11000011000110110" => rgb <= "000000";
					when "11000011000110111" => rgb <= "000000";
					when "11000011000111000" => rgb <= "000000";
					when "11000011000111001" => rgb <= "010101";
					when "11000011000111010" => rgb <= "101010";
					when "11000011000111011" => rgb <= "101010";
					when "11000011000111100" => rgb <= "101010";
					when "11000011000111101" => rgb <= "111111";
					when "11000011000111110" => rgb <= "111111";
					when "11000011000111111" => rgb <= "111111";
					when "11000011001000000" => rgb <= "101010";
					when "11000011001000001" => rgb <= "000000";
					when "11000011001000010" => rgb <= "000000";
					when "11000011001000011" => rgb <= "000000";
					when "11000011001000100" => rgb <= "000000";
					when "11000011001000101" => rgb <= "000000";
					when "11000011001000110" => rgb <= "000000";
					when "11000011001000111" => rgb <= "000000";
					when "11000011001001000" => rgb <= "000000";
					when "11000011001001001" => rgb <= "000000";
					when "11000011001001010" => rgb <= "000000";
					when "11000011001001011" => rgb <= "000000";
					when "11000011001001100" => rgb <= "000000";
					when "11000011001001101" => rgb <= "000000";
					when "11000011001001110" => rgb <= "000000";
					when "11000011001001111" => rgb <= "000000";
					when "11000011001010000" => rgb <= "101010";
					when "11000011001010001" => rgb <= "101010";
					when "11000011001010010" => rgb <= "101010";
					when "11000011001010011" => rgb <= "101010";
					when "11000011001010100" => rgb <= "111111";
					when "11000011001010101" => rgb <= "111111";
					when "11000011001010110" => rgb <= "101010";
					when "11000011001010111" => rgb <= "111111";
					when "11000011001011000" => rgb <= "111111";
					when "11000011001011001" => rgb <= "111111";
					when "11000011001011010" => rgb <= "111111";
					when "11000011001011011" => rgb <= "101010";
					when "11000011001011100" => rgb <= "111111";
					when "11000011001011101" => rgb <= "101010";
					when "11000011001011110" => rgb <= "101010";
					when "11000011001011111" => rgb <= "000000";
					when "11000011001100000" => rgb <= "000000";
					when "11000011001100001" => rgb <= "000000";
					when "11000011001100010" => rgb <= "000000";
					when "11000011001100011" => rgb <= "000000";
					when "11000011001100100" => rgb <= "000000";
					when "11000011001100101" => rgb <= "000000";
					when "11000011001100110" => rgb <= "010101";
					when "11000011001100111" => rgb <= "111111";
					when "11000011001101000" => rgb <= "101010";
					when "11000011001101001" => rgb <= "111111";
					when "11000011001101010" => rgb <= "101010";
					when "11000011001101011" => rgb <= "111111";
					when "11000011001101100" => rgb <= "101010";
					when "11000011001101101" => rgb <= "101010";
					when "11000011001101110" => rgb <= "000000";
					when "11000011001101111" => rgb <= "000000";
					when "11000011001110000" => rgb <= "000000";
					when "11000011001110001" => rgb <= "000000";
					when "11000011001110010" => rgb <= "000000";
					when "11000011001110011" => rgb <= "000000";
					when "11000011001110100" => rgb <= "000000";
					when "11000011001110101" => rgb <= "000000";
					when "11000011001110110" => rgb <= "000000";
					when "11000011001110111" => rgb <= "000000";
					when "11000011001111000" => rgb <= "000000";
					when "11000011001111001" => rgb <= "000000";
					when "11000011001111010" => rgb <= "000000";
					when "11000011001111011" => rgb <= "000000";
					when "11000011001111100" => rgb <= "000000";
					when "11000011001111101" => rgb <= "101010";
					when "11000011001111110" => rgb <= "111111";
					when "11000011001111111" => rgb <= "111111";
					when "11000011010000000" => rgb <= "111111";
					when "11000011010000001" => rgb <= "111111";
					when "11000011010000010" => rgb <= "111111";
					when "11000011010000011" => rgb <= "111111";
					when "11000011010000100" => rgb <= "111111";
					when "11000011010000101" => rgb <= "111111";
					when "11000011010000110" => rgb <= "111111";
					when "11000011010000111" => rgb <= "111111";
					when "11000011010001000" => rgb <= "111111";
					when "11000011010001001" => rgb <= "111111";
					when "11000011010001010" => rgb <= "111111";
					when "11000011010001011" => rgb <= "101010";
					when "11000011010001100" => rgb <= "000000";
					when "11000011010001101" => rgb <= "000000";
					when "11000011010001110" => rgb <= "000000";
					when "11000011010001111" => rgb <= "000000";
					when "11000011010010000" => rgb <= "000000";
					when "11000011010010001" => rgb <= "000000";
					when "11000011010010010" => rgb <= "000000";
					when "11000011010010011" => rgb <= "000000";
					when "11000011010010100" => rgb <= "000000";
					when "11000011010010101" => rgb <= "000000";
					when "11000011010010110" => rgb <= "000000";
					when "11000011010010111" => rgb <= "000000";
					when "11000011010011000" => rgb <= "000000";
					when "11000011010011001" => rgb <= "000000";
					when "11000011010011010" => rgb <= "000000";
					when "11000011010011011" => rgb <= "000000";
					when "11000011010011100" => rgb <= "000000";
					when "11000011010011101" => rgb <= "000000";
					when "11000011010011110" => rgb <= "000000";
					when "11000011010011111" => rgb <= "000000";
					when "11000011010100000" => rgb <= "000000";
					when "11000011010100001" => rgb <= "000000";
					when "11000011010100010" => rgb <= "010101";
					when "11000011010100011" => rgb <= "111111";
					when "11000011010100100" => rgb <= "101010";
					when "11000011010100101" => rgb <= "111111";
					when "11000011010100110" => rgb <= "111111";
					when "11000011010100111" => rgb <= "111111";
					when "11000011010101000" => rgb <= "111111";
					when "11000011010101001" => rgb <= "111111";
					when "11000011010101010" => rgb <= "000000";
					when "11000011010101011" => rgb <= "000000";
					when "11000011010101100" => rgb <= "000000";
					when "11000011010101101" => rgb <= "000000";
					when "11000011010101110" => rgb <= "000000";
					when "11000011010101111" => rgb <= "000000";
					when "11000011010110000" => rgb <= "000000";
					when "11000011010110001" => rgb <= "010101";
					when "11000011010110010" => rgb <= "101010";
					when "11000011010110011" => rgb <= "101010";
					when "11000011010110100" => rgb <= "111111";
					when "11000011010110101" => rgb <= "111111";
					when "11000011010110110" => rgb <= "101010";
					when "11000011010110111" => rgb <= "111111";
					when "11000011010111000" => rgb <= "101010";
					when "11000011010111001" => rgb <= "000000";
					when "11000011010111010" => rgb <= "000000";
					when "11000011010111011" => rgb <= "000000";
					when "11000011010111100" => rgb <= "000000";
					when "11000011010111101" => rgb <= "000000";
					when "11000011010111110" => rgb <= "000000";
					when "11000011010111111" => rgb <= "000000";
					when "11000011011000000" => rgb <= "010101";
					when "11000011011000001" => rgb <= "111111";
					when "11000011011000010" => rgb <= "101010";
					when "11000011011000011" => rgb <= "111111";
					when "11000011011000100" => rgb <= "101010";
					when "11000011011000101" => rgb <= "111111";
					when "11000011011000110" => rgb <= "111111";
					when "11000011011000111" => rgb <= "111111";
					when "11000011011001000" => rgb <= "111111";
					when "11000011011001001" => rgb <= "111111";
					when "11000011011001010" => rgb <= "111111";
					when "11000011011001011" => rgb <= "101010";
					when "11000011011001100" => rgb <= "111111";
					when "11000011011001101" => rgb <= "101010";
					when "11000011011001110" => rgb <= "111111";
					when "11000011011001111" => rgb <= "101010";
					when "11000011011010000" => rgb <= "000000";
					when "11000011011010001" => rgb <= "000000";
					when "11000011011010010" => rgb <= "000000";
					when "11000011011010011" => rgb <= "000000";
					when "11000011011010100" => rgb <= "000000";
					when "11000011011010101" => rgb <= "000000";
					when "11000011011010110" => rgb <= "000000";
					when "11000011011010111" => rgb <= "101010";
					when "11000011011011000" => rgb <= "101010";
					when "11000011011011001" => rgb <= "101010";
					when "11000011011011010" => rgb <= "101010";
					when "11000011011011011" => rgb <= "111111";
					when "11000011011011100" => rgb <= "111111";
					when "11000011011011101" => rgb <= "111111";
					when "11000011011011110" => rgb <= "111111";
					when "11000011011011111" => rgb <= "111111";
					when "11000011011100000" => rgb <= "111111";
					when "11000011011100001" => rgb <= "111111";
					when "11000011011100010" => rgb <= "111111";
					when "11000011011100011" => rgb <= "101010";
					when "11000011011100100" => rgb <= "111111";
					when "11000011011100101" => rgb <= "111111";
					when "11000011011100110" => rgb <= "000000";
					when "11000011011100111" => rgb <= "000000";
					when "11000011011101000" => rgb <= "000000";
					when "11000011011101001" => rgb <= "000000";
					when "11000011011101010" => rgb <= "000000";
					when "11000011011101011" => rgb <= "000000";
					when "11000011011101100" => rgb <= "000000";
					when "11000011011101101" => rgb <= "010101";
					when "11000011011101110" => rgb <= "111111";
					when "11000011011101111" => rgb <= "101010";
					when "11000011011110000" => rgb <= "111111";
					when "11000011011110001" => rgb <= "111111";
					when "11000011011110010" => rgb <= "111111";
					when "11000011011110011" => rgb <= "101010";
					when "11000011011110100" => rgb <= "101010";
					when "11000011011110101" => rgb <= "000000";
					when "11000011011110110" => rgb <= "000000";
					when "11000011011110111" => rgb <= "000000";
					when "11000011011111000" => rgb <= "000000";
					when "11000011011111001" => rgb <= "000000";
					when "11000011011111010" => rgb <= "000000";
					when "11000011011111011" => rgb <= "000000";
					when "11000011011111100" => rgb <= "000000";
					when "11000011011111101" => rgb <= "000000";
					when "11000011011111110" => rgb <= "000000";
					when "11000011011111111" => rgb <= "000000";
					when "11000011100000000" => rgb <= "000000";
					when "11000011100000001" => rgb <= "000000";
					when "11000011100000010" => rgb <= "000000";
					when "11000011100000011" => rgb <= "000000";
					when "11000011100000100" => rgb <= "000000";
					when "11000011100000101" => rgb <= "000000";
					when "11000011100000110" => rgb <= "000000";
					when "11000011100000111" => rgb <= "000000";
					when "11000011100001000" => rgb <= "000000";
					when "11000011100001001" => rgb <= "000000";
					when "11000011100001010" => rgb <= "000000";
					when "11000011100001011" => rgb <= "010101";
					when "11000011100001100" => rgb <= "111111";
					when "11000011100001101" => rgb <= "101010";
					when "11000011100001110" => rgb <= "111111";
					when "11000011100001111" => rgb <= "111111";
					when "11000011100010000" => rgb <= "111111";
					when "11000011100010001" => rgb <= "111111";
					when "11000011100010010" => rgb <= "111111";
					when "11000011100010011" => rgb <= "111111";
					when "11000011100010100" => rgb <= "111111";
					when "11000011100010101" => rgb <= "111111";
					when "11000011100010110" => rgb <= "111111";
					when "11000011100010111" => rgb <= "111111";
					when "11000011100011000" => rgb <= "101010";
					when "11000011100011001" => rgb <= "101010";
					when "11000011100011010" => rgb <= "101010";
					when "11000011100011011" => rgb <= "000000";
					when "11000011100011100" => rgb <= "000000";
					when "11000011100011101" => rgb <= "000000";
					when "11000011100011110" => rgb <= "000000";
					when "11000011100011111" => rgb <= "000000";
					when "11000011100100000" => rgb <= "000000";
					when "11000011100100001" => rgb <= "000000";
					when "11000011100100010" => rgb <= "101010";
					when "11000011100100011" => rgb <= "101010";
					when "11000011100100100" => rgb <= "101010";
					when "11000011100100101" => rgb <= "101010";
					when "11000011100100110" => rgb <= "111111";
					when "11000011100100111" => rgb <= "111111";
					when "11000011100101000" => rgb <= "111111";
					when "11000011100101001" => rgb <= "101010";
					when "11000011100101010" => rgb <= "101010";
					when "11000011100101011" => rgb <= "101010";
					when "11000011100101100" => rgb <= "101010";
					when "11000011100101101" => rgb <= "111111";
					when "11000011100101110" => rgb <= "101010";
					when "11000011100101111" => rgb <= "101010";
					when "11000011100110000" => rgb <= "101010";
					when "11000011100110001" => rgb <= "010101";
					when "11000011100110010" => rgb <= "000000";
					when "11000011100110011" => rgb <= "000000";
					when "11000011100110100" => rgb <= "000000";
					when "11000011100110101" => rgb <= "000000";
					when "11000011100110110" => rgb <= "000000";
					when "11000011100110111" => rgb <= "000000";
					when "11000011100111000" => rgb <= "000000";
					when "11000011100111001" => rgb <= "000000";
					when "11000011100111010" => rgb <= "000000";
					when "11000011100111011" => rgb <= "000000";
					when "11000011100111100" => rgb <= "000000";
					when "11000011100111101" => rgb <= "000000";
					when "11000011100111110" => rgb <= "000000";
					when "11000011100111111" => rgb <= "000000";
					when "11000100000000000" => rgb <= "000000";
					when "11000100000000001" => rgb <= "000000";
					when "11000100000000010" => rgb <= "000000";
					when "11000100000000011" => rgb <= "000000";
					when "11000100000000100" => rgb <= "000000";
					when "11000100000000101" => rgb <= "000000";
					when "11000100000000110" => rgb <= "000000";
					when "11000100000000111" => rgb <= "000000";
					when "11000100000001000" => rgb <= "000000";
					when "11000100000001001" => rgb <= "000000";
					when "11000100000001010" => rgb <= "000000";
					when "11000100000001011" => rgb <= "000000";
					when "11000100000001100" => rgb <= "000000";
					when "11000100000001101" => rgb <= "000000";
					when "11000100000001110" => rgb <= "000000";
					when "11000100000001111" => rgb <= "000000";
					when "11000100000010000" => rgb <= "000000";
					when "11000100000010001" => rgb <= "000000";
					when "11000100000010010" => rgb <= "000000";
					when "11000100000010011" => rgb <= "000000";
					when "11000100000010100" => rgb <= "101010";
					when "11000100000010101" => rgb <= "111111";
					when "11000100000010110" => rgb <= "101010";
					when "11000100000010111" => rgb <= "111111";
					when "11000100000011000" => rgb <= "111111";
					when "11000100000011001" => rgb <= "111111";
					when "11000100000011010" => rgb <= "111111";
					when "11000100000011011" => rgb <= "111111";
					when "11000100000011100" => rgb <= "111111";
					when "11000100000011101" => rgb <= "111111";
					when "11000100000011110" => rgb <= "111111";
					when "11000100000011111" => rgb <= "111111";
					when "11000100000100000" => rgb <= "111111";
					when "11000100000100001" => rgb <= "111111";
					when "11000100000100010" => rgb <= "111111";
					when "11000100000100011" => rgb <= "000000";
					when "11000100000100100" => rgb <= "000000";
					when "11000100000100101" => rgb <= "000000";
					when "11000100000100110" => rgb <= "000000";
					when "11000100000100111" => rgb <= "000000";
					when "11000100000101000" => rgb <= "000000";
					when "11000100000101001" => rgb <= "000000";
					when "11000100000101010" => rgb <= "000000";
					when "11000100000101011" => rgb <= "000000";
					when "11000100000101100" => rgb <= "000000";
					when "11000100000101101" => rgb <= "000000";
					when "11000100000101110" => rgb <= "000000";
					when "11000100000101111" => rgb <= "000000";
					when "11000100000110000" => rgb <= "000000";
					when "11000100000110001" => rgb <= "000000";
					when "11000100000110010" => rgb <= "000000";
					when "11000100000110011" => rgb <= "000000";
					when "11000100000110100" => rgb <= "000000";
					when "11000100000110101" => rgb <= "000000";
					when "11000100000110110" => rgb <= "000000";
					when "11000100000110111" => rgb <= "000000";
					when "11000100000111000" => rgb <= "000000";
					when "11000100000111001" => rgb <= "010101";
					when "11000100000111010" => rgb <= "101010";
					when "11000100000111011" => rgb <= "101010";
					when "11000100000111100" => rgb <= "101010";
					when "11000100000111101" => rgb <= "111111";
					when "11000100000111110" => rgb <= "111111";
					when "11000100000111111" => rgb <= "111111";
					when "11000100001000000" => rgb <= "101010";
					when "11000100001000001" => rgb <= "000000";
					when "11000100001000010" => rgb <= "000000";
					when "11000100001000011" => rgb <= "000000";
					when "11000100001000100" => rgb <= "000000";
					when "11000100001000101" => rgb <= "000000";
					when "11000100001000110" => rgb <= "000000";
					when "11000100001000111" => rgb <= "000000";
					when "11000100001001000" => rgb <= "000000";
					when "11000100001001001" => rgb <= "000000";
					when "11000100001001010" => rgb <= "000000";
					when "11000100001001011" => rgb <= "000000";
					when "11000100001001100" => rgb <= "000000";
					when "11000100001001101" => rgb <= "000000";
					when "11000100001001110" => rgb <= "000000";
					when "11000100001001111" => rgb <= "000000";
					when "11000100001010000" => rgb <= "101010";
					when "11000100001010001" => rgb <= "101010";
					when "11000100001010010" => rgb <= "101010";
					when "11000100001010011" => rgb <= "101010";
					when "11000100001010100" => rgb <= "111111";
					when "11000100001010101" => rgb <= "111111";
					when "11000100001010110" => rgb <= "101010";
					when "11000100001010111" => rgb <= "111111";
					when "11000100001011000" => rgb <= "111111";
					when "11000100001011001" => rgb <= "111111";
					when "11000100001011010" => rgb <= "111111";
					when "11000100001011011" => rgb <= "101010";
					when "11000100001011100" => rgb <= "111111";
					when "11000100001011101" => rgb <= "101010";
					when "11000100001011110" => rgb <= "101010";
					when "11000100001011111" => rgb <= "000000";
					when "11000100001100000" => rgb <= "000000";
					when "11000100001100001" => rgb <= "000000";
					when "11000100001100010" => rgb <= "000000";
					when "11000100001100011" => rgb <= "000000";
					when "11000100001100100" => rgb <= "000000";
					when "11000100001100101" => rgb <= "000000";
					when "11000100001100110" => rgb <= "010101";
					when "11000100001100111" => rgb <= "111111";
					when "11000100001101000" => rgb <= "101010";
					when "11000100001101001" => rgb <= "111111";
					when "11000100001101010" => rgb <= "101010";
					when "11000100001101011" => rgb <= "111111";
					when "11000100001101100" => rgb <= "101010";
					when "11000100001101101" => rgb <= "101010";
					when "11000100001101110" => rgb <= "000000";
					when "11000100001101111" => rgb <= "000000";
					when "11000100001110000" => rgb <= "000000";
					when "11000100001110001" => rgb <= "000000";
					when "11000100001110010" => rgb <= "000000";
					when "11000100001110011" => rgb <= "000000";
					when "11000100001110100" => rgb <= "000000";
					when "11000100001110101" => rgb <= "000000";
					when "11000100001110110" => rgb <= "000000";
					when "11000100001110111" => rgb <= "000000";
					when "11000100001111000" => rgb <= "000000";
					when "11000100001111001" => rgb <= "000000";
					when "11000100001111010" => rgb <= "000000";
					when "11000100001111011" => rgb <= "000000";
					when "11000100001111100" => rgb <= "000000";
					when "11000100001111101" => rgb <= "101010";
					when "11000100001111110" => rgb <= "111111";
					when "11000100001111111" => rgb <= "111111";
					when "11000100010000000" => rgb <= "111111";
					when "11000100010000001" => rgb <= "111111";
					when "11000100010000010" => rgb <= "111111";
					when "11000100010000011" => rgb <= "111111";
					when "11000100010000100" => rgb <= "111111";
					when "11000100010000101" => rgb <= "111111";
					when "11000100010000110" => rgb <= "111111";
					when "11000100010000111" => rgb <= "111111";
					when "11000100010001000" => rgb <= "111111";
					when "11000100010001001" => rgb <= "111111";
					when "11000100010001010" => rgb <= "111111";
					when "11000100010001011" => rgb <= "101010";
					when "11000100010001100" => rgb <= "000000";
					when "11000100010001101" => rgb <= "000000";
					when "11000100010001110" => rgb <= "000000";
					when "11000100010001111" => rgb <= "000000";
					when "11000100010010000" => rgb <= "000000";
					when "11000100010010001" => rgb <= "000000";
					when "11000100010010010" => rgb <= "000000";
					when "11000100010010011" => rgb <= "000000";
					when "11000100010010100" => rgb <= "000000";
					when "11000100010010101" => rgb <= "000000";
					when "11000100010010110" => rgb <= "000000";
					when "11000100010010111" => rgb <= "000000";
					when "11000100010011000" => rgb <= "000000";
					when "11000100010011001" => rgb <= "000000";
					when "11000100010011010" => rgb <= "000000";
					when "11000100010011011" => rgb <= "000000";
					when "11000100010011100" => rgb <= "000000";
					when "11000100010011101" => rgb <= "000000";
					when "11000100010011110" => rgb <= "000000";
					when "11000100010011111" => rgb <= "000000";
					when "11000100010100000" => rgb <= "000000";
					when "11000100010100001" => rgb <= "000000";
					when "11000100010100010" => rgb <= "010101";
					when "11000100010100011" => rgb <= "111111";
					when "11000100010100100" => rgb <= "101010";
					when "11000100010100101" => rgb <= "111111";
					when "11000100010100110" => rgb <= "111111";
					when "11000100010100111" => rgb <= "111111";
					when "11000100010101000" => rgb <= "111111";
					when "11000100010101001" => rgb <= "111111";
					when "11000100010101010" => rgb <= "000000";
					when "11000100010101011" => rgb <= "000000";
					when "11000100010101100" => rgb <= "000000";
					when "11000100010101101" => rgb <= "000000";
					when "11000100010101110" => rgb <= "000000";
					when "11000100010101111" => rgb <= "000000";
					when "11000100010110000" => rgb <= "000000";
					when "11000100010110001" => rgb <= "010101";
					when "11000100010110010" => rgb <= "101010";
					when "11000100010110011" => rgb <= "101010";
					when "11000100010110100" => rgb <= "111111";
					when "11000100010110101" => rgb <= "111111";
					when "11000100010110110" => rgb <= "101010";
					when "11000100010110111" => rgb <= "111111";
					when "11000100010111000" => rgb <= "101010";
					when "11000100010111001" => rgb <= "000000";
					when "11000100010111010" => rgb <= "000000";
					when "11000100010111011" => rgb <= "000000";
					when "11000100010111100" => rgb <= "000000";
					when "11000100010111101" => rgb <= "000000";
					when "11000100010111110" => rgb <= "000000";
					when "11000100010111111" => rgb <= "000000";
					when "11000100011000000" => rgb <= "010101";
					when "11000100011000001" => rgb <= "111111";
					when "11000100011000010" => rgb <= "101010";
					when "11000100011000011" => rgb <= "111111";
					when "11000100011000100" => rgb <= "101010";
					when "11000100011000101" => rgb <= "111111";
					when "11000100011000110" => rgb <= "111111";
					when "11000100011000111" => rgb <= "111111";
					when "11000100011001000" => rgb <= "111111";
					when "11000100011001001" => rgb <= "111111";
					when "11000100011001010" => rgb <= "111111";
					when "11000100011001011" => rgb <= "101010";
					when "11000100011001100" => rgb <= "111111";
					when "11000100011001101" => rgb <= "101010";
					when "11000100011001110" => rgb <= "111111";
					when "11000100011001111" => rgb <= "101010";
					when "11000100011010000" => rgb <= "000000";
					when "11000100011010001" => rgb <= "000000";
					when "11000100011010010" => rgb <= "000000";
					when "11000100011010011" => rgb <= "000000";
					when "11000100011010100" => rgb <= "000000";
					when "11000100011010101" => rgb <= "000000";
					when "11000100011010110" => rgb <= "000000";
					when "11000100011010111" => rgb <= "101010";
					when "11000100011011000" => rgb <= "101010";
					when "11000100011011001" => rgb <= "101010";
					when "11000100011011010" => rgb <= "101010";
					when "11000100011011011" => rgb <= "111111";
					when "11000100011011100" => rgb <= "111111";
					when "11000100011011101" => rgb <= "111111";
					when "11000100011011110" => rgb <= "111111";
					when "11000100011011111" => rgb <= "111111";
					when "11000100011100000" => rgb <= "111111";
					when "11000100011100001" => rgb <= "111111";
					when "11000100011100010" => rgb <= "111111";
					when "11000100011100011" => rgb <= "101010";
					when "11000100011100100" => rgb <= "111111";
					when "11000100011100101" => rgb <= "111111";
					when "11000100011100110" => rgb <= "000000";
					when "11000100011100111" => rgb <= "000000";
					when "11000100011101000" => rgb <= "000000";
					when "11000100011101001" => rgb <= "000000";
					when "11000100011101010" => rgb <= "000000";
					when "11000100011101011" => rgb <= "000000";
					when "11000100011101100" => rgb <= "000000";
					when "11000100011101101" => rgb <= "010101";
					when "11000100011101110" => rgb <= "111111";
					when "11000100011101111" => rgb <= "101010";
					when "11000100011110000" => rgb <= "111111";
					when "11000100011110001" => rgb <= "111111";
					when "11000100011110010" => rgb <= "111111";
					when "11000100011110011" => rgb <= "101010";
					when "11000100011110100" => rgb <= "101010";
					when "11000100011110101" => rgb <= "000000";
					when "11000100011110110" => rgb <= "000000";
					when "11000100011110111" => rgb <= "000000";
					when "11000100011111000" => rgb <= "000000";
					when "11000100011111001" => rgb <= "000000";
					when "11000100011111010" => rgb <= "000000";
					when "11000100011111011" => rgb <= "000000";
					when "11000100011111100" => rgb <= "000000";
					when "11000100011111101" => rgb <= "000000";
					when "11000100011111110" => rgb <= "000000";
					when "11000100011111111" => rgb <= "000000";
					when "11000100100000000" => rgb <= "000000";
					when "11000100100000001" => rgb <= "000000";
					when "11000100100000010" => rgb <= "000000";
					when "11000100100000011" => rgb <= "000000";
					when "11000100100000100" => rgb <= "000000";
					when "11000100100000101" => rgb <= "000000";
					when "11000100100000110" => rgb <= "000000";
					when "11000100100000111" => rgb <= "000000";
					when "11000100100001000" => rgb <= "000000";
					when "11000100100001001" => rgb <= "000000";
					when "11000100100001010" => rgb <= "000000";
					when "11000100100001011" => rgb <= "010101";
					when "11000100100001100" => rgb <= "111111";
					when "11000100100001101" => rgb <= "101010";
					when "11000100100001110" => rgb <= "111111";
					when "11000100100001111" => rgb <= "111111";
					when "11000100100010000" => rgb <= "111111";
					when "11000100100010001" => rgb <= "111111";
					when "11000100100010010" => rgb <= "111111";
					when "11000100100010011" => rgb <= "111111";
					when "11000100100010100" => rgb <= "111111";
					when "11000100100010101" => rgb <= "111111";
					when "11000100100010110" => rgb <= "111111";
					when "11000100100010111" => rgb <= "111111";
					when "11000100100011000" => rgb <= "101010";
					when "11000100100011001" => rgb <= "101010";
					when "11000100100011010" => rgb <= "101010";
					when "11000100100011011" => rgb <= "000000";
					when "11000100100011100" => rgb <= "000000";
					when "11000100100011101" => rgb <= "000000";
					when "11000100100011110" => rgb <= "000000";
					when "11000100100011111" => rgb <= "000000";
					when "11000100100100000" => rgb <= "000000";
					when "11000100100100001" => rgb <= "000000";
					when "11000100100100010" => rgb <= "101010";
					when "11000100100100011" => rgb <= "111111";
					when "11000100100100100" => rgb <= "101010";
					when "11000100100100101" => rgb <= "101010";
					when "11000100100100110" => rgb <= "111111";
					when "11000100100100111" => rgb <= "101010";
					when "11000100100101000" => rgb <= "101010";
					when "11000100100101001" => rgb <= "101010";
					when "11000100100101010" => rgb <= "101010";
					when "11000100100101011" => rgb <= "101010";
					when "11000100100101100" => rgb <= "101010";
					when "11000100100101101" => rgb <= "101010";
					when "11000100100101110" => rgb <= "101010";
					when "11000100100101111" => rgb <= "101010";
					when "11000100100110000" => rgb <= "111111";
					when "11000100100110001" => rgb <= "010101";
					when "11000100100110010" => rgb <= "000000";
					when "11000100100110011" => rgb <= "000000";
					when "11000100100110100" => rgb <= "000000";
					when "11000100100110101" => rgb <= "000000";
					when "11000100100110110" => rgb <= "000000";
					when "11000100100110111" => rgb <= "000000";
					when "11000100100111000" => rgb <= "000000";
					when "11000100100111001" => rgb <= "000000";
					when "11000100100111010" => rgb <= "000000";
					when "11000100100111011" => rgb <= "000000";
					when "11000100100111100" => rgb <= "000000";
					when "11000100100111101" => rgb <= "000000";
					when "11000100100111110" => rgb <= "000000";
					when "11000100100111111" => rgb <= "000000";
					when "11000101000000000" => rgb <= "000000";
					when "11000101000000001" => rgb <= "000000";
					when "11000101000000010" => rgb <= "000000";
					when "11000101000000011" => rgb <= "000000";
					when "11000101000000100" => rgb <= "000000";
					when "11000101000000101" => rgb <= "000000";
					when "11000101000000110" => rgb <= "000000";
					when "11000101000000111" => rgb <= "000000";
					when "11000101000001000" => rgb <= "000000";
					when "11000101000001001" => rgb <= "000000";
					when "11000101000001010" => rgb <= "000000";
					when "11000101000001011" => rgb <= "000000";
					when "11000101000001100" => rgb <= "000000";
					when "11000101000001101" => rgb <= "000000";
					when "11000101000001110" => rgb <= "000000";
					when "11000101000001111" => rgb <= "000000";
					when "11000101000010000" => rgb <= "000000";
					when "11000101000010001" => rgb <= "000000";
					when "11000101000010010" => rgb <= "000000";
					when "11000101000010011" => rgb <= "000000";
					when "11000101000010100" => rgb <= "101010";
					when "11000101000010101" => rgb <= "111111";
					when "11000101000010110" => rgb <= "101010";
					when "11000101000010111" => rgb <= "111111";
					when "11000101000011000" => rgb <= "111111";
					when "11000101000011001" => rgb <= "111111";
					when "11000101000011010" => rgb <= "111111";
					when "11000101000011011" => rgb <= "111111";
					when "11000101000011100" => rgb <= "111111";
					when "11000101000011101" => rgb <= "111111";
					when "11000101000011110" => rgb <= "111111";
					when "11000101000011111" => rgb <= "111111";
					when "11000101000100000" => rgb <= "111111";
					when "11000101000100001" => rgb <= "101010";
					when "11000101000100010" => rgb <= "111111";
					when "11000101000100011" => rgb <= "000000";
					when "11000101000100100" => rgb <= "000000";
					when "11000101000100101" => rgb <= "000000";
					when "11000101000100110" => rgb <= "000000";
					when "11000101000100111" => rgb <= "000000";
					when "11000101000101000" => rgb <= "000000";
					when "11000101000101001" => rgb <= "000000";
					when "11000101000101010" => rgb <= "000000";
					when "11000101000101011" => rgb <= "000000";
					when "11000101000101100" => rgb <= "000000";
					when "11000101000101101" => rgb <= "000000";
					when "11000101000101110" => rgb <= "000000";
					when "11000101000101111" => rgb <= "000000";
					when "11000101000110000" => rgb <= "000000";
					when "11000101000110001" => rgb <= "000000";
					when "11000101000110010" => rgb <= "000000";
					when "11000101000110011" => rgb <= "000000";
					when "11000101000110100" => rgb <= "000000";
					when "11000101000110101" => rgb <= "000000";
					when "11000101000110110" => rgb <= "000000";
					when "11000101000110111" => rgb <= "000000";
					when "11000101000111000" => rgb <= "000000";
					when "11000101000111001" => rgb <= "010101";
					when "11000101000111010" => rgb <= "101010";
					when "11000101000111011" => rgb <= "101010";
					when "11000101000111100" => rgb <= "101010";
					when "11000101000111101" => rgb <= "111111";
					when "11000101000111110" => rgb <= "111111";
					when "11000101000111111" => rgb <= "111111";
					when "11000101001000000" => rgb <= "101010";
					when "11000101001000001" => rgb <= "000000";
					when "11000101001000010" => rgb <= "000000";
					when "11000101001000011" => rgb <= "000000";
					when "11000101001000100" => rgb <= "000000";
					when "11000101001000101" => rgb <= "000000";
					when "11000101001000110" => rgb <= "000000";
					when "11000101001000111" => rgb <= "000000";
					when "11000101001001000" => rgb <= "000000";
					when "11000101001001001" => rgb <= "000000";
					when "11000101001001010" => rgb <= "000000";
					when "11000101001001011" => rgb <= "000000";
					when "11000101001001100" => rgb <= "000000";
					when "11000101001001101" => rgb <= "000000";
					when "11000101001001110" => rgb <= "000000";
					when "11000101001001111" => rgb <= "000000";
					when "11000101001010000" => rgb <= "101010";
					when "11000101001010001" => rgb <= "101010";
					when "11000101001010010" => rgb <= "101010";
					when "11000101001010011" => rgb <= "101010";
					when "11000101001010100" => rgb <= "111111";
					when "11000101001010101" => rgb <= "111111";
					when "11000101001010110" => rgb <= "101010";
					when "11000101001010111" => rgb <= "111111";
					when "11000101001011000" => rgb <= "111111";
					when "11000101001011001" => rgb <= "111111";
					when "11000101001011010" => rgb <= "111111";
					when "11000101001011011" => rgb <= "101010";
					when "11000101001011100" => rgb <= "111111";
					when "11000101001011101" => rgb <= "101010";
					when "11000101001011110" => rgb <= "101010";
					when "11000101001011111" => rgb <= "000000";
					when "11000101001100000" => rgb <= "000000";
					when "11000101001100001" => rgb <= "000000";
					when "11000101001100010" => rgb <= "000000";
					when "11000101001100011" => rgb <= "000000";
					when "11000101001100100" => rgb <= "000000";
					when "11000101001100101" => rgb <= "000000";
					when "11000101001100110" => rgb <= "010101";
					when "11000101001100111" => rgb <= "111111";
					when "11000101001101000" => rgb <= "101010";
					when "11000101001101001" => rgb <= "111111";
					when "11000101001101010" => rgb <= "101010";
					when "11000101001101011" => rgb <= "111111";
					when "11000101001101100" => rgb <= "101010";
					when "11000101001101101" => rgb <= "101010";
					when "11000101001101110" => rgb <= "000000";
					when "11000101001101111" => rgb <= "000000";
					when "11000101001110000" => rgb <= "000000";
					when "11000101001110001" => rgb <= "000000";
					when "11000101001110010" => rgb <= "000000";
					when "11000101001110011" => rgb <= "000000";
					when "11000101001110100" => rgb <= "000000";
					when "11000101001110101" => rgb <= "000000";
					when "11000101001110110" => rgb <= "000000";
					when "11000101001110111" => rgb <= "000000";
					when "11000101001111000" => rgb <= "000000";
					when "11000101001111001" => rgb <= "000000";
					when "11000101001111010" => rgb <= "000000";
					when "11000101001111011" => rgb <= "000000";
					when "11000101001111100" => rgb <= "000000";
					when "11000101001111101" => rgb <= "101010";
					when "11000101001111110" => rgb <= "111111";
					when "11000101001111111" => rgb <= "111111";
					when "11000101010000000" => rgb <= "111111";
					when "11000101010000001" => rgb <= "111111";
					when "11000101010000010" => rgb <= "111111";
					when "11000101010000011" => rgb <= "111111";
					when "11000101010000100" => rgb <= "111111";
					when "11000101010000101" => rgb <= "111111";
					when "11000101010000110" => rgb <= "111111";
					when "11000101010000111" => rgb <= "111111";
					when "11000101010001000" => rgb <= "111111";
					when "11000101010001001" => rgb <= "111111";
					when "11000101010001010" => rgb <= "111111";
					when "11000101010001011" => rgb <= "101010";
					when "11000101010001100" => rgb <= "000000";
					when "11000101010001101" => rgb <= "000000";
					when "11000101010001110" => rgb <= "000000";
					when "11000101010001111" => rgb <= "000000";
					when "11000101010010000" => rgb <= "000000";
					when "11000101010010001" => rgb <= "000000";
					when "11000101010010010" => rgb <= "000000";
					when "11000101010010011" => rgb <= "000000";
					when "11000101010010100" => rgb <= "000000";
					when "11000101010010101" => rgb <= "000000";
					when "11000101010010110" => rgb <= "000000";
					when "11000101010010111" => rgb <= "000000";
					when "11000101010011000" => rgb <= "000000";
					when "11000101010011001" => rgb <= "000000";
					when "11000101010011010" => rgb <= "000000";
					when "11000101010011011" => rgb <= "000000";
					when "11000101010011100" => rgb <= "000000";
					when "11000101010011101" => rgb <= "000000";
					when "11000101010011110" => rgb <= "000000";
					when "11000101010011111" => rgb <= "000000";
					when "11000101010100000" => rgb <= "000000";
					when "11000101010100001" => rgb <= "000000";
					when "11000101010100010" => rgb <= "010101";
					when "11000101010100011" => rgb <= "111111";
					when "11000101010100100" => rgb <= "101010";
					when "11000101010100101" => rgb <= "111111";
					when "11000101010100110" => rgb <= "111111";
					when "11000101010100111" => rgb <= "111111";
					when "11000101010101000" => rgb <= "111111";
					when "11000101010101001" => rgb <= "111111";
					when "11000101010101010" => rgb <= "000000";
					when "11000101010101011" => rgb <= "000000";
					when "11000101010101100" => rgb <= "000000";
					when "11000101010101101" => rgb <= "000000";
					when "11000101010101110" => rgb <= "000000";
					when "11000101010101111" => rgb <= "000000";
					when "11000101010110000" => rgb <= "000000";
					when "11000101010110001" => rgb <= "010101";
					when "11000101010110010" => rgb <= "101010";
					when "11000101010110011" => rgb <= "101010";
					when "11000101010110100" => rgb <= "111111";
					when "11000101010110101" => rgb <= "111111";
					when "11000101010110110" => rgb <= "101010";
					when "11000101010110111" => rgb <= "111111";
					when "11000101010111000" => rgb <= "101010";
					when "11000101010111001" => rgb <= "000000";
					when "11000101010111010" => rgb <= "000000";
					when "11000101010111011" => rgb <= "000000";
					when "11000101010111100" => rgb <= "000000";
					when "11000101010111101" => rgb <= "000000";
					when "11000101010111110" => rgb <= "000000";
					when "11000101010111111" => rgb <= "000000";
					when "11000101011000000" => rgb <= "010101";
					when "11000101011000001" => rgb <= "111111";
					when "11000101011000010" => rgb <= "101010";
					when "11000101011000011" => rgb <= "111111";
					when "11000101011000100" => rgb <= "101010";
					when "11000101011000101" => rgb <= "111111";
					when "11000101011000110" => rgb <= "111111";
					when "11000101011000111" => rgb <= "111111";
					when "11000101011001000" => rgb <= "111111";
					when "11000101011001001" => rgb <= "111111";
					when "11000101011001010" => rgb <= "111111";
					when "11000101011001011" => rgb <= "101010";
					when "11000101011001100" => rgb <= "111111";
					when "11000101011001101" => rgb <= "101010";
					when "11000101011001110" => rgb <= "111111";
					when "11000101011001111" => rgb <= "101010";
					when "11000101011010000" => rgb <= "000000";
					when "11000101011010001" => rgb <= "000000";
					when "11000101011010010" => rgb <= "000000";
					when "11000101011010011" => rgb <= "000000";
					when "11000101011010100" => rgb <= "000000";
					when "11000101011010101" => rgb <= "000000";
					when "11000101011010110" => rgb <= "000000";
					when "11000101011010111" => rgb <= "101010";
					when "11000101011011000" => rgb <= "101010";
					when "11000101011011001" => rgb <= "101010";
					when "11000101011011010" => rgb <= "101010";
					when "11000101011011011" => rgb <= "111111";
					when "11000101011011100" => rgb <= "111111";
					when "11000101011011101" => rgb <= "111111";
					when "11000101011011110" => rgb <= "111111";
					when "11000101011011111" => rgb <= "111111";
					when "11000101011100000" => rgb <= "111111";
					when "11000101011100001" => rgb <= "111111";
					when "11000101011100010" => rgb <= "111111";
					when "11000101011100011" => rgb <= "101010";
					when "11000101011100100" => rgb <= "111111";
					when "11000101011100101" => rgb <= "111111";
					when "11000101011100110" => rgb <= "000000";
					when "11000101011100111" => rgb <= "000000";
					when "11000101011101000" => rgb <= "000000";
					when "11000101011101001" => rgb <= "000000";
					when "11000101011101010" => rgb <= "000000";
					when "11000101011101011" => rgb <= "000000";
					when "11000101011101100" => rgb <= "000000";
					when "11000101011101101" => rgb <= "010101";
					when "11000101011101110" => rgb <= "111111";
					when "11000101011101111" => rgb <= "101010";
					when "11000101011110000" => rgb <= "111111";
					when "11000101011110001" => rgb <= "111111";
					when "11000101011110010" => rgb <= "111111";
					when "11000101011110011" => rgb <= "101010";
					when "11000101011110100" => rgb <= "101010";
					when "11000101011110101" => rgb <= "000000";
					when "11000101011110110" => rgb <= "000000";
					when "11000101011110111" => rgb <= "000000";
					when "11000101011111000" => rgb <= "000000";
					when "11000101011111001" => rgb <= "000000";
					when "11000101011111010" => rgb <= "000000";
					when "11000101011111011" => rgb <= "000000";
					when "11000101011111100" => rgb <= "000000";
					when "11000101011111101" => rgb <= "000000";
					when "11000101011111110" => rgb <= "000000";
					when "11000101011111111" => rgb <= "000000";
					when "11000101100000000" => rgb <= "000000";
					when "11000101100000001" => rgb <= "000000";
					when "11000101100000010" => rgb <= "000000";
					when "11000101100000011" => rgb <= "000000";
					when "11000101100000100" => rgb <= "000000";
					when "11000101100000101" => rgb <= "000000";
					when "11000101100000110" => rgb <= "000000";
					when "11000101100000111" => rgb <= "000000";
					when "11000101100001000" => rgb <= "000000";
					when "11000101100001001" => rgb <= "000000";
					when "11000101100001010" => rgb <= "000000";
					when "11000101100001011" => rgb <= "010101";
					when "11000101100001100" => rgb <= "111111";
					when "11000101100001101" => rgb <= "101010";
					when "11000101100001110" => rgb <= "111111";
					when "11000101100001111" => rgb <= "111111";
					when "11000101100010000" => rgb <= "111111";
					when "11000101100010001" => rgb <= "111111";
					when "11000101100010010" => rgb <= "111111";
					when "11000101100010011" => rgb <= "111111";
					when "11000101100010100" => rgb <= "111111";
					when "11000101100010101" => rgb <= "111111";
					when "11000101100010110" => rgb <= "111111";
					when "11000101100010111" => rgb <= "111111";
					when "11000101100011000" => rgb <= "101010";
					when "11000101100011001" => rgb <= "101010";
					when "11000101100011010" => rgb <= "101010";
					when "11000101100011011" => rgb <= "000000";
					when "11000101100011100" => rgb <= "000000";
					when "11000101100011101" => rgb <= "000000";
					when "11000101100011110" => rgb <= "000000";
					when "11000101100011111" => rgb <= "000000";
					when "11000101100100000" => rgb <= "000000";
					when "11000101100100001" => rgb <= "000000";
					when "11000101100100010" => rgb <= "101010";
					when "11000101100100011" => rgb <= "101010";
					when "11000101100100100" => rgb <= "101010";
					when "11000101100100101" => rgb <= "111111";
					when "11000101100100110" => rgb <= "101010";
					when "11000101100100111" => rgb <= "111111";
					when "11000101100101000" => rgb <= "101010";
					when "11000101100101001" => rgb <= "101010";
					when "11000101100101010" => rgb <= "101010";
					when "11000101100101011" => rgb <= "101010";
					when "11000101100101100" => rgb <= "111111";
					when "11000101100101101" => rgb <= "111111";
					when "11000101100101110" => rgb <= "101010";
					when "11000101100101111" => rgb <= "101010";
					when "11000101100110000" => rgb <= "101010";
					when "11000101100110001" => rgb <= "010101";
					when "11000101100110010" => rgb <= "000000";
					when "11000101100110011" => rgb <= "000000";
					when "11000101100110100" => rgb <= "000000";
					when "11000101100110101" => rgb <= "000000";
					when "11000101100110110" => rgb <= "000000";
					when "11000101100110111" => rgb <= "000000";
					when "11000101100111000" => rgb <= "000000";
					when "11000101100111001" => rgb <= "000000";
					when "11000101100111010" => rgb <= "000000";
					when "11000101100111011" => rgb <= "000000";
					when "11000101100111100" => rgb <= "000000";
					when "11000101100111101" => rgb <= "000000";
					when "11000101100111110" => rgb <= "000000";
					when "11000101100111111" => rgb <= "000000";
					when "11000110000000000" => rgb <= "000000";
					when "11000110000000001" => rgb <= "000000";
					when "11000110000000010" => rgb <= "000000";
					when "11000110000000011" => rgb <= "000000";
					when "11000110000000100" => rgb <= "000000";
					when "11000110000000101" => rgb <= "000000";
					when "11000110000000110" => rgb <= "000000";
					when "11000110000000111" => rgb <= "000000";
					when "11000110000001000" => rgb <= "000000";
					when "11000110000001001" => rgb <= "000000";
					when "11000110000001010" => rgb <= "000000";
					when "11000110000001011" => rgb <= "000000";
					when "11000110000001100" => rgb <= "000000";
					when "11000110000001101" => rgb <= "000000";
					when "11000110000001110" => rgb <= "000000";
					when "11000110000001111" => rgb <= "000000";
					when "11000110000010000" => rgb <= "000000";
					when "11000110000010001" => rgb <= "000000";
					when "11000110000010010" => rgb <= "000000";
					when "11000110000010011" => rgb <= "000000";
					when "11000110000010100" => rgb <= "101010";
					when "11000110000010101" => rgb <= "111111";
					when "11000110000010110" => rgb <= "101010";
					when "11000110000010111" => rgb <= "111111";
					when "11000110000011000" => rgb <= "111111";
					when "11000110000011001" => rgb <= "111111";
					when "11000110000011010" => rgb <= "111111";
					when "11000110000011011" => rgb <= "111111";
					when "11000110000011100" => rgb <= "111111";
					when "11000110000011101" => rgb <= "111111";
					when "11000110000011110" => rgb <= "111111";
					when "11000110000011111" => rgb <= "111111";
					when "11000110000100000" => rgb <= "111111";
					when "11000110000100001" => rgb <= "101010";
					when "11000110000100010" => rgb <= "101010";
					when "11000110000100011" => rgb <= "000000";
					when "11000110000100100" => rgb <= "000000";
					when "11000110000100101" => rgb <= "000000";
					when "11000110000100110" => rgb <= "000000";
					when "11000110000100111" => rgb <= "000000";
					when "11000110000101000" => rgb <= "000000";
					when "11000110000101001" => rgb <= "000000";
					when "11000110000101010" => rgb <= "000000";
					when "11000110000101011" => rgb <= "000000";
					when "11000110000101100" => rgb <= "000000";
					when "11000110000101101" => rgb <= "000000";
					when "11000110000101110" => rgb <= "000000";
					when "11000110000101111" => rgb <= "000000";
					when "11000110000110000" => rgb <= "000000";
					when "11000110000110001" => rgb <= "000000";
					when "11000110000110010" => rgb <= "000000";
					when "11000110000110011" => rgb <= "000000";
					when "11000110000110100" => rgb <= "000000";
					when "11000110000110101" => rgb <= "000000";
					when "11000110000110110" => rgb <= "000000";
					when "11000110000110111" => rgb <= "000000";
					when "11000110000111000" => rgb <= "000000";
					when "11000110000111001" => rgb <= "010101";
					when "11000110000111010" => rgb <= "101010";
					when "11000110000111011" => rgb <= "101010";
					when "11000110000111100" => rgb <= "101010";
					when "11000110000111101" => rgb <= "111111";
					when "11000110000111110" => rgb <= "111111";
					when "11000110000111111" => rgb <= "111111";
					when "11000110001000000" => rgb <= "101010";
					when "11000110001000001" => rgb <= "000000";
					when "11000110001000010" => rgb <= "000000";
					when "11000110001000011" => rgb <= "000000";
					when "11000110001000100" => rgb <= "000000";
					when "11000110001000101" => rgb <= "000000";
					when "11000110001000110" => rgb <= "000000";
					when "11000110001000111" => rgb <= "000000";
					when "11000110001001000" => rgb <= "000000";
					when "11000110001001001" => rgb <= "000000";
					when "11000110001001010" => rgb <= "000000";
					when "11000110001001011" => rgb <= "000000";
					when "11000110001001100" => rgb <= "000000";
					when "11000110001001101" => rgb <= "000000";
					when "11000110001001110" => rgb <= "000000";
					when "11000110001001111" => rgb <= "000000";
					when "11000110001010000" => rgb <= "101010";
					when "11000110001010001" => rgb <= "101010";
					when "11000110001010010" => rgb <= "101010";
					when "11000110001010011" => rgb <= "101010";
					when "11000110001010100" => rgb <= "111111";
					when "11000110001010101" => rgb <= "111111";
					when "11000110001010110" => rgb <= "101010";
					when "11000110001010111" => rgb <= "111111";
					when "11000110001011000" => rgb <= "111111";
					when "11000110001011001" => rgb <= "111111";
					when "11000110001011010" => rgb <= "111111";
					when "11000110001011011" => rgb <= "101010";
					when "11000110001011100" => rgb <= "111111";
					when "11000110001011101" => rgb <= "101010";
					when "11000110001011110" => rgb <= "101010";
					when "11000110001011111" => rgb <= "000000";
					when "11000110001100000" => rgb <= "000000";
					when "11000110001100001" => rgb <= "000000";
					when "11000110001100010" => rgb <= "000000";
					when "11000110001100011" => rgb <= "000000";
					when "11000110001100100" => rgb <= "000000";
					when "11000110001100101" => rgb <= "000000";
					when "11000110001100110" => rgb <= "010101";
					when "11000110001100111" => rgb <= "111111";
					when "11000110001101000" => rgb <= "101010";
					when "11000110001101001" => rgb <= "111111";
					when "11000110001101010" => rgb <= "101010";
					when "11000110001101011" => rgb <= "111111";
					when "11000110001101100" => rgb <= "101010";
					when "11000110001101101" => rgb <= "101010";
					when "11000110001101110" => rgb <= "000000";
					when "11000110001101111" => rgb <= "000000";
					when "11000110001110000" => rgb <= "000000";
					when "11000110001110001" => rgb <= "000000";
					when "11000110001110010" => rgb <= "000000";
					when "11000110001110011" => rgb <= "000000";
					when "11000110001110100" => rgb <= "000000";
					when "11000110001110101" => rgb <= "000000";
					when "11000110001110110" => rgb <= "000000";
					when "11000110001110111" => rgb <= "000000";
					when "11000110001111000" => rgb <= "000000";
					when "11000110001111001" => rgb <= "000000";
					when "11000110001111010" => rgb <= "000000";
					when "11000110001111011" => rgb <= "000000";
					when "11000110001111100" => rgb <= "000000";
					when "11000110001111101" => rgb <= "101010";
					when "11000110001111110" => rgb <= "111111";
					when "11000110001111111" => rgb <= "111111";
					when "11000110010000000" => rgb <= "111111";
					when "11000110010000001" => rgb <= "111111";
					when "11000110010000010" => rgb <= "111111";
					when "11000110010000011" => rgb <= "111111";
					when "11000110010000100" => rgb <= "111111";
					when "11000110010000101" => rgb <= "111111";
					when "11000110010000110" => rgb <= "111111";
					when "11000110010000111" => rgb <= "111111";
					when "11000110010001000" => rgb <= "111111";
					when "11000110010001001" => rgb <= "111111";
					when "11000110010001010" => rgb <= "111111";
					when "11000110010001011" => rgb <= "101010";
					when "11000110010001100" => rgb <= "000000";
					when "11000110010001101" => rgb <= "000000";
					when "11000110010001110" => rgb <= "000000";
					when "11000110010001111" => rgb <= "000000";
					when "11000110010010000" => rgb <= "000000";
					when "11000110010010001" => rgb <= "000000";
					when "11000110010010010" => rgb <= "000000";
					when "11000110010010011" => rgb <= "000000";
					when "11000110010010100" => rgb <= "000000";
					when "11000110010010101" => rgb <= "000000";
					when "11000110010010110" => rgb <= "000000";
					when "11000110010010111" => rgb <= "000000";
					when "11000110010011000" => rgb <= "000000";
					when "11000110010011001" => rgb <= "000000";
					when "11000110010011010" => rgb <= "000000";
					when "11000110010011011" => rgb <= "000000";
					when "11000110010011100" => rgb <= "000000";
					when "11000110010011101" => rgb <= "000000";
					when "11000110010011110" => rgb <= "000000";
					when "11000110010011111" => rgb <= "000000";
					when "11000110010100000" => rgb <= "000000";
					when "11000110010100001" => rgb <= "000000";
					when "11000110010100010" => rgb <= "010101";
					when "11000110010100011" => rgb <= "111111";
					when "11000110010100100" => rgb <= "101010";
					when "11000110010100101" => rgb <= "111111";
					when "11000110010100110" => rgb <= "111111";
					when "11000110010100111" => rgb <= "111111";
					when "11000110010101000" => rgb <= "111111";
					when "11000110010101001" => rgb <= "111111";
					when "11000110010101010" => rgb <= "000000";
					when "11000110010101011" => rgb <= "000000";
					when "11000110010101100" => rgb <= "000000";
					when "11000110010101101" => rgb <= "000000";
					when "11000110010101110" => rgb <= "000000";
					when "11000110010101111" => rgb <= "000000";
					when "11000110010110000" => rgb <= "000000";
					when "11000110010110001" => rgb <= "010101";
					when "11000110010110010" => rgb <= "101010";
					when "11000110010110011" => rgb <= "101010";
					when "11000110010110100" => rgb <= "111111";
					when "11000110010110101" => rgb <= "111111";
					when "11000110010110110" => rgb <= "101010";
					when "11000110010110111" => rgb <= "111111";
					when "11000110010111000" => rgb <= "101010";
					when "11000110010111001" => rgb <= "000000";
					when "11000110010111010" => rgb <= "000000";
					when "11000110010111011" => rgb <= "000000";
					when "11000110010111100" => rgb <= "000000";
					when "11000110010111101" => rgb <= "000000";
					when "11000110010111110" => rgb <= "000000";
					when "11000110010111111" => rgb <= "000000";
					when "11000110011000000" => rgb <= "010101";
					when "11000110011000001" => rgb <= "111111";
					when "11000110011000010" => rgb <= "101010";
					when "11000110011000011" => rgb <= "111111";
					when "11000110011000100" => rgb <= "101010";
					when "11000110011000101" => rgb <= "111111";
					when "11000110011000110" => rgb <= "111111";
					when "11000110011000111" => rgb <= "111111";
					when "11000110011001000" => rgb <= "111111";
					when "11000110011001001" => rgb <= "111111";
					when "11000110011001010" => rgb <= "111111";
					when "11000110011001011" => rgb <= "101010";
					when "11000110011001100" => rgb <= "111111";
					when "11000110011001101" => rgb <= "101010";
					when "11000110011001110" => rgb <= "111111";
					when "11000110011001111" => rgb <= "101010";
					when "11000110011010000" => rgb <= "000000";
					when "11000110011010001" => rgb <= "000000";
					when "11000110011010010" => rgb <= "000000";
					when "11000110011010011" => rgb <= "000000";
					when "11000110011010100" => rgb <= "000000";
					when "11000110011010101" => rgb <= "000000";
					when "11000110011010110" => rgb <= "000000";
					when "11000110011010111" => rgb <= "101010";
					when "11000110011011000" => rgb <= "101010";
					when "11000110011011001" => rgb <= "101010";
					when "11000110011011010" => rgb <= "101010";
					when "11000110011011011" => rgb <= "111111";
					when "11000110011011100" => rgb <= "111111";
					when "11000110011011101" => rgb <= "111111";
					when "11000110011011110" => rgb <= "111111";
					when "11000110011011111" => rgb <= "111111";
					when "11000110011100000" => rgb <= "111111";
					when "11000110011100001" => rgb <= "111111";
					when "11000110011100010" => rgb <= "111111";
					when "11000110011100011" => rgb <= "101010";
					when "11000110011100100" => rgb <= "111111";
					when "11000110011100101" => rgb <= "111111";
					when "11000110011100110" => rgb <= "000000";
					when "11000110011100111" => rgb <= "000000";
					when "11000110011101000" => rgb <= "000000";
					when "11000110011101001" => rgb <= "000000";
					when "11000110011101010" => rgb <= "000000";
					when "11000110011101011" => rgb <= "000000";
					when "11000110011101100" => rgb <= "000000";
					when "11000110011101101" => rgb <= "010101";
					when "11000110011101110" => rgb <= "111111";
					when "11000110011101111" => rgb <= "101010";
					when "11000110011110000" => rgb <= "111111";
					when "11000110011110001" => rgb <= "111111";
					when "11000110011110010" => rgb <= "111111";
					when "11000110011110011" => rgb <= "101010";
					when "11000110011110100" => rgb <= "101010";
					when "11000110011110101" => rgb <= "000000";
					when "11000110011110110" => rgb <= "000000";
					when "11000110011110111" => rgb <= "000000";
					when "11000110011111000" => rgb <= "000000";
					when "11000110011111001" => rgb <= "000000";
					when "11000110011111010" => rgb <= "000000";
					when "11000110011111011" => rgb <= "000000";
					when "11000110011111100" => rgb <= "000000";
					when "11000110011111101" => rgb <= "000000";
					when "11000110011111110" => rgb <= "000000";
					when "11000110011111111" => rgb <= "000000";
					when "11000110100000000" => rgb <= "000000";
					when "11000110100000001" => rgb <= "000000";
					when "11000110100000010" => rgb <= "000000";
					when "11000110100000011" => rgb <= "000000";
					when "11000110100000100" => rgb <= "000000";
					when "11000110100000101" => rgb <= "000000";
					when "11000110100000110" => rgb <= "000000";
					when "11000110100000111" => rgb <= "000000";
					when "11000110100001000" => rgb <= "000000";
					when "11000110100001001" => rgb <= "000000";
					when "11000110100001010" => rgb <= "000000";
					when "11000110100001011" => rgb <= "010101";
					when "11000110100001100" => rgb <= "111111";
					when "11000110100001101" => rgb <= "101010";
					when "11000110100001110" => rgb <= "111111";
					when "11000110100001111" => rgb <= "111111";
					when "11000110100010000" => rgb <= "111111";
					when "11000110100010001" => rgb <= "111111";
					when "11000110100010010" => rgb <= "111111";
					when "11000110100010011" => rgb <= "111111";
					when "11000110100010100" => rgb <= "111111";
					when "11000110100010101" => rgb <= "111111";
					when "11000110100010110" => rgb <= "111111";
					when "11000110100010111" => rgb <= "111111";
					when "11000110100011000" => rgb <= "101010";
					when "11000110100011001" => rgb <= "111111";
					when "11000110100011010" => rgb <= "101010";
					when "11000110100011011" => rgb <= "000000";
					when "11000110100011100" => rgb <= "000000";
					when "11000110100011101" => rgb <= "000000";
					when "11000110100011110" => rgb <= "000000";
					when "11000110100011111" => rgb <= "000000";
					when "11000110100100000" => rgb <= "000000";
					when "11000110100100001" => rgb <= "000000";
					when "11000110100100010" => rgb <= "010101";
					when "11000110100100011" => rgb <= "010101";
					when "11000110100100100" => rgb <= "010101";
					when "11000110100100101" => rgb <= "010101";
					when "11000110100100110" => rgb <= "010101";
					when "11000110100100111" => rgb <= "010101";
					when "11000110100101000" => rgb <= "010101";
					when "11000110100101001" => rgb <= "010101";
					when "11000110100101010" => rgb <= "010101";
					when "11000110100101011" => rgb <= "010101";
					when "11000110100101100" => rgb <= "010101";
					when "11000110100101101" => rgb <= "010101";
					when "11000110100101110" => rgb <= "010101";
					when "11000110100101111" => rgb <= "010101";
					when "11000110100110000" => rgb <= "010101";
					when "11000110100110001" => rgb <= "000000";
					when "11000110100110010" => rgb <= "000000";
					when "11000110100110011" => rgb <= "000000";
					when "11000110100110100" => rgb <= "000000";
					when "11000110100110101" => rgb <= "000000";
					when "11000110100110110" => rgb <= "000000";
					when "11000110100110111" => rgb <= "000000";
					when "11000110100111000" => rgb <= "000000";
					when "11000110100111001" => rgb <= "000000";
					when "11000110100111010" => rgb <= "000000";
					when "11000110100111011" => rgb <= "000000";
					when "11000110100111100" => rgb <= "000000";
					when "11000110100111101" => rgb <= "000000";
					when "11000110100111110" => rgb <= "000000";
					when "11000110100111111" => rgb <= "000000";
					when "11000111000000000" => rgb <= "000000";
					when "11000111000000001" => rgb <= "000000";
					when "11000111000000010" => rgb <= "000000";
					when "11000111000000011" => rgb <= "000000";
					when "11000111000000100" => rgb <= "000000";
					when "11000111000000101" => rgb <= "000000";
					when "11000111000000110" => rgb <= "000000";
					when "11000111000000111" => rgb <= "000000";
					when "11000111000001000" => rgb <= "000000";
					when "11000111000001001" => rgb <= "000000";
					when "11000111000001010" => rgb <= "000000";
					when "11000111000001011" => rgb <= "000000";
					when "11000111000001100" => rgb <= "000000";
					when "11000111000001101" => rgb <= "000000";
					when "11000111000001110" => rgb <= "000000";
					when "11000111000001111" => rgb <= "000000";
					when "11000111000010000" => rgb <= "000000";
					when "11000111000010001" => rgb <= "000000";
					when "11000111000010010" => rgb <= "000000";
					when "11000111000010011" => rgb <= "000000";
					when "11000111000010100" => rgb <= "101010";
					when "11000111000010101" => rgb <= "111111";
					when "11000111000010110" => rgb <= "101010";
					when "11000111000010111" => rgb <= "111111";
					when "11000111000011000" => rgb <= "111111";
					when "11000111000011001" => rgb <= "111111";
					when "11000111000011010" => rgb <= "111111";
					when "11000111000011011" => rgb <= "111111";
					when "11000111000011100" => rgb <= "111111";
					when "11000111000011101" => rgb <= "111111";
					when "11000111000011110" => rgb <= "111111";
					when "11000111000011111" => rgb <= "111111";
					when "11000111000100000" => rgb <= "111111";
					when "11000111000100001" => rgb <= "111111";
					when "11000111000100010" => rgb <= "111111";
					when "11000111000100011" => rgb <= "000000";
					when "11000111000100100" => rgb <= "000000";
					when "11000111000100101" => rgb <= "000000";
					when "11000111000100110" => rgb <= "000000";
					when "11000111000100111" => rgb <= "000000";
					when "11000111000101000" => rgb <= "000000";
					when "11000111000101001" => rgb <= "000000";
					when "11000111000101010" => rgb <= "000000";
					when "11000111000101011" => rgb <= "000000";
					when "11000111000101100" => rgb <= "000000";
					when "11000111000101101" => rgb <= "000000";
					when "11000111000101110" => rgb <= "000000";
					when "11000111000101111" => rgb <= "000000";
					when "11000111000110000" => rgb <= "000000";
					when "11000111000110001" => rgb <= "000000";
					when "11000111000110010" => rgb <= "000000";
					when "11000111000110011" => rgb <= "000000";
					when "11000111000110100" => rgb <= "000000";
					when "11000111000110101" => rgb <= "000000";
					when "11000111000110110" => rgb <= "000000";
					when "11000111000110111" => rgb <= "000000";
					when "11000111000111000" => rgb <= "000000";
					when "11000111000111001" => rgb <= "010101";
					when "11000111000111010" => rgb <= "101010";
					when "11000111000111011" => rgb <= "101010";
					when "11000111000111100" => rgb <= "101010";
					when "11000111000111101" => rgb <= "111111";
					when "11000111000111110" => rgb <= "111111";
					when "11000111000111111" => rgb <= "111111";
					when "11000111001000000" => rgb <= "101010";
					when "11000111001000001" => rgb <= "000000";
					when "11000111001000010" => rgb <= "000000";
					when "11000111001000011" => rgb <= "000000";
					when "11000111001000100" => rgb <= "000000";
					when "11000111001000101" => rgb <= "000000";
					when "11000111001000110" => rgb <= "000000";
					when "11000111001000111" => rgb <= "000000";
					when "11000111001001000" => rgb <= "000000";
					when "11000111001001001" => rgb <= "000000";
					when "11000111001001010" => rgb <= "000000";
					when "11000111001001011" => rgb <= "000000";
					when "11000111001001100" => rgb <= "000000";
					when "11000111001001101" => rgb <= "000000";
					when "11000111001001110" => rgb <= "000000";
					when "11000111001001111" => rgb <= "000000";
					when "11000111001010000" => rgb <= "101010";
					when "11000111001010001" => rgb <= "101010";
					when "11000111001010010" => rgb <= "101010";
					when "11000111001010011" => rgb <= "101010";
					when "11000111001010100" => rgb <= "111111";
					when "11000111001010101" => rgb <= "111111";
					when "11000111001010110" => rgb <= "101010";
					when "11000111001010111" => rgb <= "111111";
					when "11000111001011000" => rgb <= "111111";
					when "11000111001011001" => rgb <= "111111";
					when "11000111001011010" => rgb <= "111111";
					when "11000111001011011" => rgb <= "101010";
					when "11000111001011100" => rgb <= "111111";
					when "11000111001011101" => rgb <= "101010";
					when "11000111001011110" => rgb <= "101010";
					when "11000111001011111" => rgb <= "000000";
					when "11000111001100000" => rgb <= "000000";
					when "11000111001100001" => rgb <= "000000";
					when "11000111001100010" => rgb <= "000000";
					when "11000111001100011" => rgb <= "000000";
					when "11000111001100100" => rgb <= "000000";
					when "11000111001100101" => rgb <= "000000";
					when "11000111001100110" => rgb <= "010101";
					when "11000111001100111" => rgb <= "111111";
					when "11000111001101000" => rgb <= "101010";
					when "11000111001101001" => rgb <= "111111";
					when "11000111001101010" => rgb <= "101010";
					when "11000111001101011" => rgb <= "111111";
					when "11000111001101100" => rgb <= "101010";
					when "11000111001101101" => rgb <= "101010";
					when "11000111001101110" => rgb <= "000000";
					when "11000111001101111" => rgb <= "000000";
					when "11000111001110000" => rgb <= "000000";
					when "11000111001110001" => rgb <= "000000";
					when "11000111001110010" => rgb <= "000000";
					when "11000111001110011" => rgb <= "000000";
					when "11000111001110100" => rgb <= "000000";
					when "11000111001110101" => rgb <= "000000";
					when "11000111001110110" => rgb <= "000000";
					when "11000111001110111" => rgb <= "000000";
					when "11000111001111000" => rgb <= "000000";
					when "11000111001111001" => rgb <= "000000";
					when "11000111001111010" => rgb <= "000000";
					when "11000111001111011" => rgb <= "000000";
					when "11000111001111100" => rgb <= "000000";
					when "11000111001111101" => rgb <= "101010";
					when "11000111001111110" => rgb <= "111111";
					when "11000111001111111" => rgb <= "111111";
					when "11000111010000000" => rgb <= "111111";
					when "11000111010000001" => rgb <= "111111";
					when "11000111010000010" => rgb <= "111111";
					when "11000111010000011" => rgb <= "111111";
					when "11000111010000100" => rgb <= "111111";
					when "11000111010000101" => rgb <= "111111";
					when "11000111010000110" => rgb <= "111111";
					when "11000111010000111" => rgb <= "111111";
					when "11000111010001000" => rgb <= "111111";
					when "11000111010001001" => rgb <= "111111";
					when "11000111010001010" => rgb <= "111111";
					when "11000111010001011" => rgb <= "101010";
					when "11000111010001100" => rgb <= "000000";
					when "11000111010001101" => rgb <= "000000";
					when "11000111010001110" => rgb <= "000000";
					when "11000111010001111" => rgb <= "000000";
					when "11000111010010000" => rgb <= "000000";
					when "11000111010010001" => rgb <= "000000";
					when "11000111010010010" => rgb <= "000000";
					when "11000111010010011" => rgb <= "000000";
					when "11000111010010100" => rgb <= "000000";
					when "11000111010010101" => rgb <= "000000";
					when "11000111010010110" => rgb <= "000000";
					when "11000111010010111" => rgb <= "000000";
					when "11000111010011000" => rgb <= "000000";
					when "11000111010011001" => rgb <= "000000";
					when "11000111010011010" => rgb <= "000000";
					when "11000111010011011" => rgb <= "000000";
					when "11000111010011100" => rgb <= "000000";
					when "11000111010011101" => rgb <= "000000";
					when "11000111010011110" => rgb <= "000000";
					when "11000111010011111" => rgb <= "000000";
					when "11000111010100000" => rgb <= "000000";
					when "11000111010100001" => rgb <= "000000";
					when "11000111010100010" => rgb <= "010101";
					when "11000111010100011" => rgb <= "111111";
					when "11000111010100100" => rgb <= "101010";
					when "11000111010100101" => rgb <= "111111";
					when "11000111010100110" => rgb <= "111111";
					when "11000111010100111" => rgb <= "111111";
					when "11000111010101000" => rgb <= "111111";
					when "11000111010101001" => rgb <= "111111";
					when "11000111010101010" => rgb <= "000000";
					when "11000111010101011" => rgb <= "000000";
					when "11000111010101100" => rgb <= "000000";
					when "11000111010101101" => rgb <= "000000";
					when "11000111010101110" => rgb <= "000000";
					when "11000111010101111" => rgb <= "000000";
					when "11000111010110000" => rgb <= "000000";
					when "11000111010110001" => rgb <= "010101";
					when "11000111010110010" => rgb <= "101010";
					when "11000111010110011" => rgb <= "101010";
					when "11000111010110100" => rgb <= "111111";
					when "11000111010110101" => rgb <= "111111";
					when "11000111010110110" => rgb <= "101010";
					when "11000111010110111" => rgb <= "111111";
					when "11000111010111000" => rgb <= "101010";
					when "11000111010111001" => rgb <= "000000";
					when "11000111010111010" => rgb <= "000000";
					when "11000111010111011" => rgb <= "000000";
					when "11000111010111100" => rgb <= "000000";
					when "11000111010111101" => rgb <= "000000";
					when "11000111010111110" => rgb <= "000000";
					when "11000111010111111" => rgb <= "000000";
					when "11000111011000000" => rgb <= "010101";
					when "11000111011000001" => rgb <= "111111";
					when "11000111011000010" => rgb <= "101010";
					when "11000111011000011" => rgb <= "111111";
					when "11000111011000100" => rgb <= "101010";
					when "11000111011000101" => rgb <= "111111";
					when "11000111011000110" => rgb <= "111111";
					when "11000111011000111" => rgb <= "111111";
					when "11000111011001000" => rgb <= "111111";
					when "11000111011001001" => rgb <= "111111";
					when "11000111011001010" => rgb <= "111111";
					when "11000111011001011" => rgb <= "101010";
					when "11000111011001100" => rgb <= "111111";
					when "11000111011001101" => rgb <= "101010";
					when "11000111011001110" => rgb <= "111111";
					when "11000111011001111" => rgb <= "101010";
					when "11000111011010000" => rgb <= "000000";
					when "11000111011010001" => rgb <= "000000";
					when "11000111011010010" => rgb <= "000000";
					when "11000111011010011" => rgb <= "000000";
					when "11000111011010100" => rgb <= "000000";
					when "11000111011010101" => rgb <= "000000";
					when "11000111011010110" => rgb <= "000000";
					when "11000111011010111" => rgb <= "101010";
					when "11000111011011000" => rgb <= "101010";
					when "11000111011011001" => rgb <= "101010";
					when "11000111011011010" => rgb <= "101010";
					when "11000111011011011" => rgb <= "111111";
					when "11000111011011100" => rgb <= "111111";
					when "11000111011011101" => rgb <= "111111";
					when "11000111011011110" => rgb <= "111111";
					when "11000111011011111" => rgb <= "111111";
					when "11000111011100000" => rgb <= "111111";
					when "11000111011100001" => rgb <= "111111";
					when "11000111011100010" => rgb <= "111111";
					when "11000111011100011" => rgb <= "101010";
					when "11000111011100100" => rgb <= "111111";
					when "11000111011100101" => rgb <= "111111";
					when "11000111011100110" => rgb <= "000000";
					when "11000111011100111" => rgb <= "000000";
					when "11000111011101000" => rgb <= "000000";
					when "11000111011101001" => rgb <= "000000";
					when "11000111011101010" => rgb <= "000000";
					when "11000111011101011" => rgb <= "000000";
					when "11000111011101100" => rgb <= "000000";
					when "11000111011101101" => rgb <= "010101";
					when "11000111011101110" => rgb <= "111111";
					when "11000111011101111" => rgb <= "101010";
					when "11000111011110000" => rgb <= "111111";
					when "11000111011110001" => rgb <= "111111";
					when "11000111011110010" => rgb <= "111111";
					when "11000111011110011" => rgb <= "101010";
					when "11000111011110100" => rgb <= "101010";
					when "11000111011110101" => rgb <= "000000";
					when "11000111011110110" => rgb <= "000000";
					when "11000111011110111" => rgb <= "000000";
					when "11000111011111000" => rgb <= "000000";
					when "11000111011111001" => rgb <= "000000";
					when "11000111011111010" => rgb <= "000000";
					when "11000111011111011" => rgb <= "000000";
					when "11000111011111100" => rgb <= "000000";
					when "11000111011111101" => rgb <= "000000";
					when "11000111011111110" => rgb <= "000000";
					when "11000111011111111" => rgb <= "000000";
					when "11000111100000000" => rgb <= "000000";
					when "11000111100000001" => rgb <= "000000";
					when "11000111100000010" => rgb <= "000000";
					when "11000111100000011" => rgb <= "000000";
					when "11000111100000100" => rgb <= "000000";
					when "11000111100000101" => rgb <= "000000";
					when "11000111100000110" => rgb <= "000000";
					when "11000111100000111" => rgb <= "000000";
					when "11000111100001000" => rgb <= "000000";
					when "11000111100001001" => rgb <= "000000";
					when "11000111100001010" => rgb <= "000000";
					when "11000111100001011" => rgb <= "010101";
					when "11000111100001100" => rgb <= "111111";
					when "11000111100001101" => rgb <= "101010";
					when "11000111100001110" => rgb <= "111111";
					when "11000111100001111" => rgb <= "111111";
					when "11000111100010000" => rgb <= "111111";
					when "11000111100010001" => rgb <= "111111";
					when "11000111100010010" => rgb <= "111111";
					when "11000111100010011" => rgb <= "111111";
					when "11000111100010100" => rgb <= "111111";
					when "11000111100010101" => rgb <= "111111";
					when "11000111100010110" => rgb <= "111111";
					when "11000111100010111" => rgb <= "111111";
					when "11000111100011000" => rgb <= "101010";
					when "11000111100011001" => rgb <= "111111";
					when "11000111100011010" => rgb <= "101010";
					when "11000111100011011" => rgb <= "000000";
					when "11000111100011100" => rgb <= "000000";
					when "11000111100011101" => rgb <= "000000";
					when "11000111100011110" => rgb <= "000000";
					when "11000111100011111" => rgb <= "000000";
					when "11000111100100000" => rgb <= "000000";
					when "11000111100100001" => rgb <= "000000";
					when "11000111100100010" => rgb <= "000000";
					when "11000111100100011" => rgb <= "000000";
					when "11000111100100100" => rgb <= "000000";
					when "11000111100100101" => rgb <= "000000";
					when "11000111100100110" => rgb <= "000000";
					when "11000111100100111" => rgb <= "000000";
					when "11000111100101000" => rgb <= "000000";
					when "11000111100101001" => rgb <= "000000";
					when "11000111100101010" => rgb <= "000000";
					when "11000111100101011" => rgb <= "000000";
					when "11000111100101100" => rgb <= "000000";
					when "11000111100101101" => rgb <= "000000";
					when "11000111100101110" => rgb <= "000000";
					when "11000111100101111" => rgb <= "000000";
					when "11000111100110000" => rgb <= "000000";
					when "11000111100110001" => rgb <= "000000";
					when "11000111100110010" => rgb <= "000000";
					when "11000111100110011" => rgb <= "000000";
					when "11000111100110100" => rgb <= "000000";
					when "11000111100110101" => rgb <= "000000";
					when "11000111100110110" => rgb <= "000000";
					when "11000111100110111" => rgb <= "000000";
					when "11000111100111000" => rgb <= "000000";
					when "11000111100111001" => rgb <= "000000";
					when "11000111100111010" => rgb <= "000000";
					when "11000111100111011" => rgb <= "000000";
					when "11000111100111100" => rgb <= "000000";
					when "11000111100111101" => rgb <= "000000";
					when "11000111100111110" => rgb <= "000000";
					when "11000111100111111" => rgb <= "000000";
					when "11001000000000000" => rgb <= "000000";
					when "11001000000000001" => rgb <= "000000";
					when "11001000000000010" => rgb <= "000000";
					when "11001000000000011" => rgb <= "000000";
					when "11001000000000100" => rgb <= "000000";
					when "11001000000000101" => rgb <= "000000";
					when "11001000000000110" => rgb <= "000000";
					when "11001000000000111" => rgb <= "000000";
					when "11001000000001000" => rgb <= "000000";
					when "11001000000001001" => rgb <= "000000";
					when "11001000000001010" => rgb <= "000000";
					when "11001000000001011" => rgb <= "000000";
					when "11001000000001100" => rgb <= "000000";
					when "11001000000001101" => rgb <= "000000";
					when "11001000000001110" => rgb <= "000000";
					when "11001000000001111" => rgb <= "000000";
					when "11001000000010000" => rgb <= "000000";
					when "11001000000010001" => rgb <= "000000";
					when "11001000000010010" => rgb <= "000000";
					when "11001000000010011" => rgb <= "000000";
					when "11001000000010100" => rgb <= "101010";
					when "11001000000010101" => rgb <= "111111";
					when "11001000000010110" => rgb <= "101010";
					when "11001000000010111" => rgb <= "111111";
					when "11001000000011000" => rgb <= "111111";
					when "11001000000011001" => rgb <= "111111";
					when "11001000000011010" => rgb <= "111111";
					when "11001000000011011" => rgb <= "111111";
					when "11001000000011100" => rgb <= "111111";
					when "11001000000011101" => rgb <= "111111";
					when "11001000000011110" => rgb <= "111111";
					when "11001000000011111" => rgb <= "111111";
					when "11001000000100000" => rgb <= "111111";
					when "11001000000100001" => rgb <= "101010";
					when "11001000000100010" => rgb <= "111111";
					when "11001000000100011" => rgb <= "000000";
					when "11001000000100100" => rgb <= "000000";
					when "11001000000100101" => rgb <= "000000";
					when "11001000000100110" => rgb <= "000000";
					when "11001000000100111" => rgb <= "000000";
					when "11001000000101000" => rgb <= "000000";
					when "11001000000101001" => rgb <= "000000";
					when "11001000000101010" => rgb <= "000000";
					when "11001000000101011" => rgb <= "000000";
					when "11001000000101100" => rgb <= "000000";
					when "11001000000101101" => rgb <= "000000";
					when "11001000000101110" => rgb <= "000000";
					when "11001000000101111" => rgb <= "000000";
					when "11001000000110000" => rgb <= "000000";
					when "11001000000110001" => rgb <= "000000";
					when "11001000000110010" => rgb <= "000000";
					when "11001000000110011" => rgb <= "000000";
					when "11001000000110100" => rgb <= "000000";
					when "11001000000110101" => rgb <= "000000";
					when "11001000000110110" => rgb <= "000000";
					when "11001000000110111" => rgb <= "000000";
					when "11001000000111000" => rgb <= "000000";
					when "11001000000111001" => rgb <= "010101";
					when "11001000000111010" => rgb <= "101010";
					when "11001000000111011" => rgb <= "101010";
					when "11001000000111100" => rgb <= "101010";
					when "11001000000111101" => rgb <= "111111";
					when "11001000000111110" => rgb <= "111111";
					when "11001000000111111" => rgb <= "101010";
					when "11001000001000000" => rgb <= "101010";
					when "11001000001000001" => rgb <= "000000";
					when "11001000001000010" => rgb <= "000000";
					when "11001000001000011" => rgb <= "000000";
					when "11001000001000100" => rgb <= "000000";
					when "11001000001000101" => rgb <= "000000";
					when "11001000001000110" => rgb <= "000000";
					when "11001000001000111" => rgb <= "000000";
					when "11001000001001000" => rgb <= "000000";
					when "11001000001001001" => rgb <= "000000";
					when "11001000001001010" => rgb <= "000000";
					when "11001000001001011" => rgb <= "000000";
					when "11001000001001100" => rgb <= "000000";
					when "11001000001001101" => rgb <= "000000";
					when "11001000001001110" => rgb <= "000000";
					when "11001000001001111" => rgb <= "000000";
					when "11001000001010000" => rgb <= "101010";
					when "11001000001010001" => rgb <= "101010";
					when "11001000001010010" => rgb <= "101010";
					when "11001000001010011" => rgb <= "101010";
					when "11001000001010100" => rgb <= "111111";
					when "11001000001010101" => rgb <= "101010";
					when "11001000001010110" => rgb <= "101010";
					when "11001000001010111" => rgb <= "111111";
					when "11001000001011000" => rgb <= "111111";
					when "11001000001011001" => rgb <= "111111";
					when "11001000001011010" => rgb <= "111111";
					when "11001000001011011" => rgb <= "101010";
					when "11001000001011100" => rgb <= "111111";
					when "11001000001011101" => rgb <= "101010";
					when "11001000001011110" => rgb <= "101010";
					when "11001000001011111" => rgb <= "000000";
					when "11001000001100000" => rgb <= "000000";
					when "11001000001100001" => rgb <= "000000";
					when "11001000001100010" => rgb <= "000000";
					when "11001000001100011" => rgb <= "000000";
					when "11001000001100100" => rgb <= "000000";
					when "11001000001100101" => rgb <= "000000";
					when "11001000001100110" => rgb <= "010101";
					when "11001000001100111" => rgb <= "111111";
					when "11001000001101000" => rgb <= "101010";
					when "11001000001101001" => rgb <= "101010";
					when "11001000001101010" => rgb <= "101010";
					when "11001000001101011" => rgb <= "111111";
					when "11001000001101100" => rgb <= "111111";
					when "11001000001101101" => rgb <= "111111";
					when "11001000001101110" => rgb <= "000000";
					when "11001000001101111" => rgb <= "000000";
					when "11001000001110000" => rgb <= "000000";
					when "11001000001110001" => rgb <= "000000";
					when "11001000001110010" => rgb <= "000000";
					when "11001000001110011" => rgb <= "000000";
					when "11001000001110100" => rgb <= "000000";
					when "11001000001110101" => rgb <= "000000";
					when "11001000001110110" => rgb <= "000000";
					when "11001000001110111" => rgb <= "000000";
					when "11001000001111000" => rgb <= "000000";
					when "11001000001111001" => rgb <= "000000";
					when "11001000001111010" => rgb <= "000000";
					when "11001000001111011" => rgb <= "000000";
					when "11001000001111100" => rgb <= "000000";
					when "11001000001111101" => rgb <= "101010";
					when "11001000001111110" => rgb <= "111111";
					when "11001000001111111" => rgb <= "101010";
					when "11001000010000000" => rgb <= "111111";
					when "11001000010000001" => rgb <= "111111";
					when "11001000010000010" => rgb <= "111111";
					when "11001000010000011" => rgb <= "111111";
					when "11001000010000100" => rgb <= "101010";
					when "11001000010000101" => rgb <= "111111";
					when "11001000010000110" => rgb <= "111111";
					when "11001000010000111" => rgb <= "101010";
					when "11001000010001000" => rgb <= "111111";
					when "11001000010001001" => rgb <= "101010";
					when "11001000010001010" => rgb <= "101010";
					when "11001000010001011" => rgb <= "101010";
					when "11001000010001100" => rgb <= "000000";
					when "11001000010001101" => rgb <= "000000";
					when "11001000010001110" => rgb <= "000000";
					when "11001000010001111" => rgb <= "000000";
					when "11001000010010000" => rgb <= "000000";
					when "11001000010010001" => rgb <= "000000";
					when "11001000010010010" => rgb <= "000000";
					when "11001000010010011" => rgb <= "000000";
					when "11001000010010100" => rgb <= "000000";
					when "11001000010010101" => rgb <= "000000";
					when "11001000010010110" => rgb <= "000000";
					when "11001000010010111" => rgb <= "000000";
					when "11001000010011000" => rgb <= "000000";
					when "11001000010011001" => rgb <= "000000";
					when "11001000010011010" => rgb <= "000000";
					when "11001000010011011" => rgb <= "000000";
					when "11001000010011100" => rgb <= "000000";
					when "11001000010011101" => rgb <= "000000";
					when "11001000010011110" => rgb <= "000000";
					when "11001000010011111" => rgb <= "000000";
					when "11001000010100000" => rgb <= "000000";
					when "11001000010100001" => rgb <= "000000";
					when "11001000010100010" => rgb <= "010101";
					when "11001000010100011" => rgb <= "111111";
					when "11001000010100100" => rgb <= "101010";
					when "11001000010100101" => rgb <= "111111";
					when "11001000010100110" => rgb <= "111111";
					when "11001000010100111" => rgb <= "111111";
					when "11001000010101000" => rgb <= "101010";
					when "11001000010101001" => rgb <= "111111";
					when "11001000010101010" => rgb <= "000000";
					when "11001000010101011" => rgb <= "000000";
					when "11001000010101100" => rgb <= "000000";
					when "11001000010101101" => rgb <= "000000";
					when "11001000010101110" => rgb <= "000000";
					when "11001000010101111" => rgb <= "000000";
					when "11001000010110000" => rgb <= "000000";
					when "11001000010110001" => rgb <= "010101";
					when "11001000010110010" => rgb <= "111111";
					when "11001000010110011" => rgb <= "101010";
					when "11001000010110100" => rgb <= "111111";
					when "11001000010110101" => rgb <= "111111";
					when "11001000010110110" => rgb <= "101010";
					when "11001000010110111" => rgb <= "101010";
					when "11001000010111000" => rgb <= "101010";
					when "11001000010111001" => rgb <= "000000";
					when "11001000010111010" => rgb <= "000000";
					when "11001000010111011" => rgb <= "000000";
					when "11001000010111100" => rgb <= "000000";
					when "11001000010111101" => rgb <= "000000";
					when "11001000010111110" => rgb <= "000000";
					when "11001000010111111" => rgb <= "000000";
					when "11001000011000000" => rgb <= "010101";
					when "11001000011000001" => rgb <= "111111";
					when "11001000011000010" => rgb <= "101010";
					when "11001000011000011" => rgb <= "111111";
					when "11001000011000100" => rgb <= "111111";
					when "11001000011000101" => rgb <= "101010";
					when "11001000011000110" => rgb <= "101010";
					when "11001000011000111" => rgb <= "111111";
					when "11001000011001000" => rgb <= "101010";
					when "11001000011001001" => rgb <= "111111";
					when "11001000011001010" => rgb <= "101010";
					when "11001000011001011" => rgb <= "101010";
					when "11001000011001100" => rgb <= "111111";
					when "11001000011001101" => rgb <= "101010";
					when "11001000011001110" => rgb <= "111111";
					when "11001000011001111" => rgb <= "101010";
					when "11001000011010000" => rgb <= "000000";
					when "11001000011010001" => rgb <= "000000";
					when "11001000011010010" => rgb <= "000000";
					when "11001000011010011" => rgb <= "000000";
					when "11001000011010100" => rgb <= "000000";
					when "11001000011010101" => rgb <= "000000";
					when "11001000011010110" => rgb <= "000000";
					when "11001000011010111" => rgb <= "101010";
					when "11001000011011000" => rgb <= "101010";
					when "11001000011011001" => rgb <= "101010";
					when "11001000011011010" => rgb <= "101010";
					when "11001000011011011" => rgb <= "111111";
					when "11001000011011100" => rgb <= "111111";
					when "11001000011011101" => rgb <= "111111";
					when "11001000011011110" => rgb <= "111111";
					when "11001000011011111" => rgb <= "111111";
					when "11001000011100000" => rgb <= "111111";
					when "11001000011100001" => rgb <= "111111";
					when "11001000011100010" => rgb <= "111111";
					when "11001000011100011" => rgb <= "101010";
					when "11001000011100100" => rgb <= "111111";
					when "11001000011100101" => rgb <= "111111";
					when "11001000011100110" => rgb <= "000000";
					when "11001000011100111" => rgb <= "000000";
					when "11001000011101000" => rgb <= "000000";
					when "11001000011101001" => rgb <= "000000";
					when "11001000011101010" => rgb <= "000000";
					when "11001000011101011" => rgb <= "000000";
					when "11001000011101100" => rgb <= "000000";
					when "11001000011101101" => rgb <= "010101";
					when "11001000011101110" => rgb <= "111111";
					when "11001000011101111" => rgb <= "101010";
					when "11001000011110000" => rgb <= "111111";
					when "11001000011110001" => rgb <= "111111";
					when "11001000011110010" => rgb <= "111111";
					when "11001000011110011" => rgb <= "101010";
					when "11001000011110100" => rgb <= "101010";
					when "11001000011110101" => rgb <= "000000";
					when "11001000011110110" => rgb <= "000000";
					when "11001000011110111" => rgb <= "000000";
					when "11001000011111000" => rgb <= "000000";
					when "11001000011111001" => rgb <= "000000";
					when "11001000011111010" => rgb <= "000000";
					when "11001000011111011" => rgb <= "000000";
					when "11001000011111100" => rgb <= "000000";
					when "11001000011111101" => rgb <= "000000";
					when "11001000011111110" => rgb <= "000000";
					when "11001000011111111" => rgb <= "000000";
					when "11001000100000000" => rgb <= "000000";
					when "11001000100000001" => rgb <= "000000";
					when "11001000100000010" => rgb <= "000000";
					when "11001000100000011" => rgb <= "000000";
					when "11001000100000100" => rgb <= "000000";
					when "11001000100000101" => rgb <= "000000";
					when "11001000100000110" => rgb <= "000000";
					when "11001000100000111" => rgb <= "000000";
					when "11001000100001000" => rgb <= "000000";
					when "11001000100001001" => rgb <= "000000";
					when "11001000100001010" => rgb <= "000000";
					when "11001000100001011" => rgb <= "010101";
					when "11001000100001100" => rgb <= "111111";
					when "11001000100001101" => rgb <= "101010";
					when "11001000100001110" => rgb <= "111111";
					when "11001000100001111" => rgb <= "111111";
					when "11001000100010000" => rgb <= "111111";
					when "11001000100010001" => rgb <= "111111";
					when "11001000100010010" => rgb <= "111111";
					when "11001000100010011" => rgb <= "111111";
					when "11001000100010100" => rgb <= "111111";
					when "11001000100010101" => rgb <= "111111";
					when "11001000100010110" => rgb <= "111111";
					when "11001000100010111" => rgb <= "111111";
					when "11001000100011000" => rgb <= "101010";
					when "11001000100011001" => rgb <= "101010";
					when "11001000100011010" => rgb <= "101010";
					when "11001000100011011" => rgb <= "000000";
					when "11001000100011100" => rgb <= "000000";
					when "11001000100011101" => rgb <= "000000";
					when "11001000100011110" => rgb <= "000000";
					when "11001000100011111" => rgb <= "000000";
					when "11001000100100000" => rgb <= "000000";
					when "11001000100100001" => rgb <= "000000";
					when "11001000100100010" => rgb <= "000000";
					when "11001000100100011" => rgb <= "000000";
					when "11001000100100100" => rgb <= "000000";
					when "11001000100100101" => rgb <= "000000";
					when "11001000100100110" => rgb <= "000000";
					when "11001000100100111" => rgb <= "000000";
					when "11001000100101000" => rgb <= "000000";
					when "11001000100101001" => rgb <= "000000";
					when "11001000100101010" => rgb <= "000000";
					when "11001000100101011" => rgb <= "000000";
					when "11001000100101100" => rgb <= "000000";
					when "11001000100101101" => rgb <= "000000";
					when "11001000100101110" => rgb <= "000000";
					when "11001000100101111" => rgb <= "000000";
					when "11001000100110000" => rgb <= "000000";
					when "11001000100110001" => rgb <= "000000";
					when "11001000100110010" => rgb <= "000000";
					when "11001000100110011" => rgb <= "000000";
					when "11001000100110100" => rgb <= "000000";
					when "11001000100110101" => rgb <= "000000";
					when "11001000100110110" => rgb <= "000000";
					when "11001000100110111" => rgb <= "000000";
					when "11001000100111000" => rgb <= "000000";
					when "11001000100111001" => rgb <= "000000";
					when "11001000100111010" => rgb <= "000000";
					when "11001000100111011" => rgb <= "000000";
					when "11001000100111100" => rgb <= "000000";
					when "11001000100111101" => rgb <= "000000";
					when "11001000100111110" => rgb <= "000000";
					when "11001000100111111" => rgb <= "000000";
					when "11001001000000000" => rgb <= "000000";
					when "11001001000000001" => rgb <= "000000";
					when "11001001000000010" => rgb <= "000000";
					when "11001001000000011" => rgb <= "000000";
					when "11001001000000100" => rgb <= "000000";
					when "11001001000000101" => rgb <= "000000";
					when "11001001000000110" => rgb <= "000000";
					when "11001001000000111" => rgb <= "000000";
					when "11001001000001000" => rgb <= "000000";
					when "11001001000001001" => rgb <= "000000";
					when "11001001000001010" => rgb <= "000000";
					when "11001001000001011" => rgb <= "000000";
					when "11001001000001100" => rgb <= "000000";
					when "11001001000001101" => rgb <= "000000";
					when "11001001000001110" => rgb <= "000000";
					when "11001001000001111" => rgb <= "000000";
					when "11001001000010000" => rgb <= "000000";
					when "11001001000010001" => rgb <= "000000";
					when "11001001000010010" => rgb <= "000000";
					when "11001001000010011" => rgb <= "000000";
					when "11001001000010100" => rgb <= "101010";
					when "11001001000010101" => rgb <= "111111";
					when "11001001000010110" => rgb <= "101010";
					when "11001001000010111" => rgb <= "111111";
					when "11001001000011000" => rgb <= "111111";
					when "11001001000011001" => rgb <= "111111";
					when "11001001000011010" => rgb <= "111111";
					when "11001001000011011" => rgb <= "111111";
					when "11001001000011100" => rgb <= "111111";
					when "11001001000011101" => rgb <= "111111";
					when "11001001000011110" => rgb <= "111111";
					when "11001001000011111" => rgb <= "111111";
					when "11001001000100000" => rgb <= "111111";
					when "11001001000100001" => rgb <= "101010";
					when "11001001000100010" => rgb <= "111111";
					when "11001001000100011" => rgb <= "000000";
					when "11001001000100100" => rgb <= "000000";
					when "11001001000100101" => rgb <= "000000";
					when "11001001000100110" => rgb <= "000000";
					when "11001001000100111" => rgb <= "000000";
					when "11001001000101000" => rgb <= "000000";
					when "11001001000101001" => rgb <= "000000";
					when "11001001000101010" => rgb <= "000000";
					when "11001001000101011" => rgb <= "000000";
					when "11001001000101100" => rgb <= "000000";
					when "11001001000101101" => rgb <= "000000";
					when "11001001000101110" => rgb <= "000000";
					when "11001001000101111" => rgb <= "000000";
					when "11001001000110000" => rgb <= "000000";
					when "11001001000110001" => rgb <= "000000";
					when "11001001000110010" => rgb <= "000000";
					when "11001001000110011" => rgb <= "000000";
					when "11001001000110100" => rgb <= "000000";
					when "11001001000110101" => rgb <= "000000";
					when "11001001000110110" => rgb <= "000000";
					when "11001001000110111" => rgb <= "000000";
					when "11001001000111000" => rgb <= "000000";
					when "11001001000111001" => rgb <= "010101";
					when "11001001000111010" => rgb <= "111111";
					when "11001001000111011" => rgb <= "101010";
					when "11001001000111100" => rgb <= "101010";
					when "11001001000111101" => rgb <= "101010";
					when "11001001000111110" => rgb <= "101010";
					when "11001001000111111" => rgb <= "111111";
					when "11001001001000000" => rgb <= "111111";
					when "11001001001000001" => rgb <= "000000";
					when "11001001001000010" => rgb <= "000000";
					when "11001001001000011" => rgb <= "000000";
					when "11001001001000100" => rgb <= "000000";
					when "11001001001000101" => rgb <= "000000";
					when "11001001001000110" => rgb <= "000000";
					when "11001001001000111" => rgb <= "000000";
					when "11001001001001000" => rgb <= "000000";
					when "11001001001001001" => rgb <= "000000";
					when "11001001001001010" => rgb <= "000000";
					when "11001001001001011" => rgb <= "000000";
					when "11001001001001100" => rgb <= "000000";
					when "11001001001001101" => rgb <= "000000";
					when "11001001001001110" => rgb <= "000000";
					when "11001001001001111" => rgb <= "000000";
					when "11001001001010000" => rgb <= "101010";
					when "11001001001010001" => rgb <= "101010";
					when "11001001001010010" => rgb <= "101010";
					when "11001001001010011" => rgb <= "101010";
					when "11001001001010100" => rgb <= "111111";
					when "11001001001010101" => rgb <= "111111";
					when "11001001001010110" => rgb <= "111111";
					when "11001001001010111" => rgb <= "101010";
					when "11001001001011000" => rgb <= "101010";
					when "11001001001011001" => rgb <= "101010";
					when "11001001001011010" => rgb <= "111111";
					when "11001001001011011" => rgb <= "111111";
					when "11001001001011100" => rgb <= "111111";
					when "11001001001011101" => rgb <= "101010";
					when "11001001001011110" => rgb <= "101010";
					when "11001001001011111" => rgb <= "000000";
					when "11001001001100000" => rgb <= "000000";
					when "11001001001100001" => rgb <= "000000";
					when "11001001001100010" => rgb <= "000000";
					when "11001001001100011" => rgb <= "000000";
					when "11001001001100100" => rgb <= "000000";
					when "11001001001100101" => rgb <= "000000";
					when "11001001001100110" => rgb <= "010101";
					when "11001001001100111" => rgb <= "101010";
					when "11001001001101000" => rgb <= "101010";
					when "11001001001101001" => rgb <= "101010";
					when "11001001001101010" => rgb <= "101010";
					when "11001001001101011" => rgb <= "111111";
					when "11001001001101100" => rgb <= "101010";
					when "11001001001101101" => rgb <= "101010";
					when "11001001001101110" => rgb <= "000000";
					when "11001001001101111" => rgb <= "000000";
					when "11001001001110000" => rgb <= "000000";
					when "11001001001110001" => rgb <= "000000";
					when "11001001001110010" => rgb <= "000000";
					when "11001001001110011" => rgb <= "000000";
					when "11001001001110100" => rgb <= "000000";
					when "11001001001110101" => rgb <= "000000";
					when "11001001001110110" => rgb <= "000000";
					when "11001001001110111" => rgb <= "000000";
					when "11001001001111000" => rgb <= "000000";
					when "11001001001111001" => rgb <= "000000";
					when "11001001001111010" => rgb <= "000000";
					when "11001001001111011" => rgb <= "000000";
					when "11001001001111100" => rgb <= "000000";
					when "11001001001111101" => rgb <= "101010";
					when "11001001001111110" => rgb <= "101010";
					when "11001001001111111" => rgb <= "111111";
					when "11001001010000000" => rgb <= "101010";
					when "11001001010000001" => rgb <= "111111";
					when "11001001010000010" => rgb <= "101010";
					when "11001001010000011" => rgb <= "111111";
					when "11001001010000100" => rgb <= "111111";
					when "11001001010000101" => rgb <= "101010";
					when "11001001010000110" => rgb <= "101010";
					when "11001001010000111" => rgb <= "111111";
					when "11001001010001000" => rgb <= "111111";
					when "11001001010001001" => rgb <= "111111";
					when "11001001010001010" => rgb <= "111111";
					when "11001001010001011" => rgb <= "101010";
					when "11001001010001100" => rgb <= "000000";
					when "11001001010001101" => rgb <= "000000";
					when "11001001010001110" => rgb <= "000000";
					when "11001001010001111" => rgb <= "000000";
					when "11001001010010000" => rgb <= "000000";
					when "11001001010010001" => rgb <= "000000";
					when "11001001010010010" => rgb <= "000000";
					when "11001001010010011" => rgb <= "000000";
					when "11001001010010100" => rgb <= "000000";
					when "11001001010010101" => rgb <= "000000";
					when "11001001010010110" => rgb <= "000000";
					when "11001001010010111" => rgb <= "000000";
					when "11001001010011000" => rgb <= "000000";
					when "11001001010011001" => rgb <= "000000";
					when "11001001010011010" => rgb <= "000000";
					when "11001001010011011" => rgb <= "000000";
					when "11001001010011100" => rgb <= "000000";
					when "11001001010011101" => rgb <= "000000";
					when "11001001010011110" => rgb <= "000000";
					when "11001001010011111" => rgb <= "000000";
					when "11001001010100000" => rgb <= "000000";
					when "11001001010100001" => rgb <= "000000";
					when "11001001010100010" => rgb <= "010101";
					when "11001001010100011" => rgb <= "101010";
					when "11001001010100100" => rgb <= "101010";
					when "11001001010100101" => rgb <= "111111";
					when "11001001010100110" => rgb <= "111111";
					when "11001001010100111" => rgb <= "101010";
					when "11001001010101000" => rgb <= "111111";
					when "11001001010101001" => rgb <= "101010";
					when "11001001010101010" => rgb <= "000000";
					when "11001001010101011" => rgb <= "000000";
					when "11001001010101100" => rgb <= "000000";
					when "11001001010101101" => rgb <= "000000";
					when "11001001010101110" => rgb <= "000000";
					when "11001001010101111" => rgb <= "000000";
					when "11001001010110000" => rgb <= "000000";
					when "11001001010110001" => rgb <= "010101";
					when "11001001010110010" => rgb <= "101010";
					when "11001001010110011" => rgb <= "111111";
					when "11001001010110100" => rgb <= "101010";
					when "11001001010110101" => rgb <= "111111";
					when "11001001010110110" => rgb <= "111111";
					when "11001001010110111" => rgb <= "111111";
					when "11001001010111000" => rgb <= "101010";
					when "11001001010111001" => rgb <= "000000";
					when "11001001010111010" => rgb <= "000000";
					when "11001001010111011" => rgb <= "000000";
					when "11001001010111100" => rgb <= "000000";
					when "11001001010111101" => rgb <= "000000";
					when "11001001010111110" => rgb <= "000000";
					when "11001001010111111" => rgb <= "000000";
					when "11001001011000000" => rgb <= "010101";
					when "11001001011000001" => rgb <= "111111";
					when "11001001011000010" => rgb <= "101010";
					when "11001001011000011" => rgb <= "101010";
					when "11001001011000100" => rgb <= "101010";
					when "11001001011000101" => rgb <= "111111";
					when "11001001011000110" => rgb <= "111111";
					when "11001001011000111" => rgb <= "101010";
					when "11001001011001000" => rgb <= "111111";
					when "11001001011001001" => rgb <= "111111";
					when "11001001011001010" => rgb <= "101010";
					when "11001001011001011" => rgb <= "101010";
					when "11001001011001100" => rgb <= "111111";
					when "11001001011001101" => rgb <= "101010";
					when "11001001011001110" => rgb <= "101010";
					when "11001001011001111" => rgb <= "101010";
					when "11001001011010000" => rgb <= "000000";
					when "11001001011010001" => rgb <= "000000";
					when "11001001011010010" => rgb <= "000000";
					when "11001001011010011" => rgb <= "000000";
					when "11001001011010100" => rgb <= "000000";
					when "11001001011010101" => rgb <= "000000";
					when "11001001011010110" => rgb <= "000000";
					when "11001001011010111" => rgb <= "101010";
					when "11001001011011000" => rgb <= "101010";
					when "11001001011011001" => rgb <= "101010";
					when "11001001011011010" => rgb <= "101010";
					when "11001001011011011" => rgb <= "111111";
					when "11001001011011100" => rgb <= "111111";
					when "11001001011011101" => rgb <= "111111";
					when "11001001011011110" => rgb <= "111111";
					when "11001001011011111" => rgb <= "111111";
					when "11001001011100000" => rgb <= "111111";
					when "11001001011100001" => rgb <= "111111";
					when "11001001011100010" => rgb <= "111111";
					when "11001001011100011" => rgb <= "101010";
					when "11001001011100100" => rgb <= "111111";
					when "11001001011100101" => rgb <= "111111";
					when "11001001011100110" => rgb <= "000000";
					when "11001001011100111" => rgb <= "000000";
					when "11001001011101000" => rgb <= "000000";
					when "11001001011101001" => rgb <= "000000";
					when "11001001011101010" => rgb <= "000000";
					when "11001001011101011" => rgb <= "000000";
					when "11001001011101100" => rgb <= "000000";
					when "11001001011101101" => rgb <= "010101";
					when "11001001011101110" => rgb <= "111111";
					when "11001001011101111" => rgb <= "101010";
					when "11001001011110000" => rgb <= "111111";
					when "11001001011110001" => rgb <= "111111";
					when "11001001011110010" => rgb <= "111111";
					when "11001001011110011" => rgb <= "101010";
					when "11001001011110100" => rgb <= "101010";
					when "11001001011110101" => rgb <= "000000";
					when "11001001011110110" => rgb <= "000000";
					when "11001001011110111" => rgb <= "000000";
					when "11001001011111000" => rgb <= "000000";
					when "11001001011111001" => rgb <= "000000";
					when "11001001011111010" => rgb <= "000000";
					when "11001001011111011" => rgb <= "000000";
					when "11001001011111100" => rgb <= "000000";
					when "11001001011111101" => rgb <= "000000";
					when "11001001011111110" => rgb <= "000000";
					when "11001001011111111" => rgb <= "000000";
					when "11001001100000000" => rgb <= "000000";
					when "11001001100000001" => rgb <= "000000";
					when "11001001100000010" => rgb <= "000000";
					when "11001001100000011" => rgb <= "000000";
					when "11001001100000100" => rgb <= "000000";
					when "11001001100000101" => rgb <= "000000";
					when "11001001100000110" => rgb <= "000000";
					when "11001001100000111" => rgb <= "000000";
					when "11001001100001000" => rgb <= "000000";
					when "11001001100001001" => rgb <= "000000";
					when "11001001100001010" => rgb <= "000000";
					when "11001001100001011" => rgb <= "010101";
					when "11001001100001100" => rgb <= "111111";
					when "11001001100001101" => rgb <= "101010";
					when "11001001100001110" => rgb <= "111111";
					when "11001001100001111" => rgb <= "111111";
					when "11001001100010000" => rgb <= "111111";
					when "11001001100010001" => rgb <= "111111";
					when "11001001100010010" => rgb <= "111111";
					when "11001001100010011" => rgb <= "111111";
					when "11001001100010100" => rgb <= "111111";
					when "11001001100010101" => rgb <= "111111";
					when "11001001100010110" => rgb <= "111111";
					when "11001001100010111" => rgb <= "111111";
					when "11001001100011000" => rgb <= "101010";
					when "11001001100011001" => rgb <= "101010";
					when "11001001100011010" => rgb <= "101010";
					when "11001001100011011" => rgb <= "000000";
					when "11001001100011100" => rgb <= "000000";
					when "11001001100011101" => rgb <= "000000";
					when "11001001100011110" => rgb <= "000000";
					when "11001001100011111" => rgb <= "000000";
					when "11001001100100000" => rgb <= "000000";
					when "11001001100100001" => rgb <= "000000";
					when "11001001100100010" => rgb <= "000000";
					when "11001001100100011" => rgb <= "000000";
					when "11001001100100100" => rgb <= "000000";
					when "11001001100100101" => rgb <= "000000";
					when "11001001100100110" => rgb <= "000000";
					when "11001001100100111" => rgb <= "000000";
					when "11001001100101000" => rgb <= "000000";
					when "11001001100101001" => rgb <= "000000";
					when "11001001100101010" => rgb <= "000000";
					when "11001001100101011" => rgb <= "000000";
					when "11001001100101100" => rgb <= "000000";
					when "11001001100101101" => rgb <= "000000";
					when "11001001100101110" => rgb <= "000000";
					when "11001001100101111" => rgb <= "000000";
					when "11001001100110000" => rgb <= "000000";
					when "11001001100110001" => rgb <= "000000";
					when "11001001100110010" => rgb <= "000000";
					when "11001001100110011" => rgb <= "000000";
					when "11001001100110100" => rgb <= "000000";
					when "11001001100110101" => rgb <= "000000";
					when "11001001100110110" => rgb <= "000000";
					when "11001001100110111" => rgb <= "000000";
					when "11001001100111000" => rgb <= "000000";
					when "11001001100111001" => rgb <= "000000";
					when "11001001100111010" => rgb <= "000000";
					when "11001001100111011" => rgb <= "000000";
					when "11001001100111100" => rgb <= "000000";
					when "11001001100111101" => rgb <= "000000";
					when "11001001100111110" => rgb <= "000000";
					when "11001001100111111" => rgb <= "000000";
					when "11001010000000000" => rgb <= "000000";
					when "11001010000000001" => rgb <= "000000";
					when "11001010000000010" => rgb <= "000000";
					when "11001010000000011" => rgb <= "000000";
					when "11001010000000100" => rgb <= "000000";
					when "11001010000000101" => rgb <= "000000";
					when "11001010000000110" => rgb <= "000000";
					when "11001010000000111" => rgb <= "000000";
					when "11001010000001000" => rgb <= "000000";
					when "11001010000001001" => rgb <= "000000";
					when "11001010000001010" => rgb <= "000000";
					when "11001010000001011" => rgb <= "000000";
					when "11001010000001100" => rgb <= "000000";
					when "11001010000001101" => rgb <= "000000";
					when "11001010000001110" => rgb <= "000000";
					when "11001010000001111" => rgb <= "000000";
					when "11001010000010000" => rgb <= "000000";
					when "11001010000010001" => rgb <= "000000";
					when "11001010000010010" => rgb <= "000000";
					when "11001010000010011" => rgb <= "000000";
					when "11001010000010100" => rgb <= "101010";
					when "11001010000010101" => rgb <= "111111";
					when "11001010000010110" => rgb <= "101010";
					when "11001010000010111" => rgb <= "111111";
					when "11001010000011000" => rgb <= "111111";
					when "11001010000011001" => rgb <= "111111";
					when "11001010000011010" => rgb <= "111111";
					when "11001010000011011" => rgb <= "111111";
					when "11001010000011100" => rgb <= "111111";
					when "11001010000011101" => rgb <= "111111";
					when "11001010000011110" => rgb <= "111111";
					when "11001010000011111" => rgb <= "111111";
					when "11001010000100000" => rgb <= "111111";
					when "11001010000100001" => rgb <= "101010";
					when "11001010000100010" => rgb <= "111111";
					when "11001010000100011" => rgb <= "000000";
					when "11001010000100100" => rgb <= "000000";
					when "11001010000100101" => rgb <= "000000";
					when "11001010000100110" => rgb <= "000000";
					when "11001010000100111" => rgb <= "000000";
					when "11001010000101000" => rgb <= "000000";
					when "11001010000101001" => rgb <= "000000";
					when "11001010000101010" => rgb <= "000000";
					when "11001010000101011" => rgb <= "000000";
					when "11001010000101100" => rgb <= "000000";
					when "11001010000101101" => rgb <= "000000";
					when "11001010000101110" => rgb <= "000000";
					when "11001010000101111" => rgb <= "000000";
					when "11001010000110000" => rgb <= "000000";
					when "11001010000110001" => rgb <= "000000";
					when "11001010000110010" => rgb <= "000000";
					when "11001010000110011" => rgb <= "000000";
					when "11001010000110100" => rgb <= "000000";
					when "11001010000110101" => rgb <= "000000";
					when "11001010000110110" => rgb <= "000000";
					when "11001010000110111" => rgb <= "000000";
					when "11001010000111000" => rgb <= "000000";
					when "11001010000111001" => rgb <= "010101";
					when "11001010000111010" => rgb <= "101010";
					when "11001010000111011" => rgb <= "101010";
					when "11001010000111100" => rgb <= "111111";
					when "11001010000111101" => rgb <= "111111";
					when "11001010000111110" => rgb <= "111111";
					when "11001010000111111" => rgb <= "111111";
					when "11001010001000000" => rgb <= "101010";
					when "11001010001000001" => rgb <= "000000";
					when "11001010001000010" => rgb <= "000000";
					when "11001010001000011" => rgb <= "000000";
					when "11001010001000100" => rgb <= "000000";
					when "11001010001000101" => rgb <= "000000";
					when "11001010001000110" => rgb <= "000000";
					when "11001010001000111" => rgb <= "000000";
					when "11001010001001000" => rgb <= "000000";
					when "11001010001001001" => rgb <= "000000";
					when "11001010001001010" => rgb <= "000000";
					when "11001010001001011" => rgb <= "000000";
					when "11001010001001100" => rgb <= "000000";
					when "11001010001001101" => rgb <= "000000";
					when "11001010001001110" => rgb <= "000000";
					when "11001010001001111" => rgb <= "000000";
					when "11001010001010000" => rgb <= "101010";
					when "11001010001010001" => rgb <= "101010";
					when "11001010001010010" => rgb <= "111111";
					when "11001010001010011" => rgb <= "111111";
					when "11001010001010100" => rgb <= "101010";
					when "11001010001010101" => rgb <= "111111";
					when "11001010001010110" => rgb <= "111111";
					when "11001010001010111" => rgb <= "111111";
					when "11001010001011000" => rgb <= "111111";
					when "11001010001011001" => rgb <= "111111";
					when "11001010001011010" => rgb <= "111111";
					when "11001010001011011" => rgb <= "101010";
					when "11001010001011100" => rgb <= "101010";
					when "11001010001011101" => rgb <= "111111";
					when "11001010001011110" => rgb <= "101010";
					when "11001010001011111" => rgb <= "000000";
					when "11001010001100000" => rgb <= "000000";
					when "11001010001100001" => rgb <= "000000";
					when "11001010001100010" => rgb <= "000000";
					when "11001010001100011" => rgb <= "000000";
					when "11001010001100100" => rgb <= "000000";
					when "11001010001100101" => rgb <= "000000";
					when "11001010001100110" => rgb <= "010101";
					when "11001010001100111" => rgb <= "111111";
					when "11001010001101000" => rgb <= "111111";
					when "11001010001101001" => rgb <= "111111";
					when "11001010001101010" => rgb <= "101010";
					when "11001010001101011" => rgb <= "111111";
					when "11001010001101100" => rgb <= "101010";
					when "11001010001101101" => rgb <= "111111";
					when "11001010001101110" => rgb <= "000000";
					when "11001010001101111" => rgb <= "000000";
					when "11001010001110000" => rgb <= "000000";
					when "11001010001110001" => rgb <= "000000";
					when "11001010001110010" => rgb <= "000000";
					when "11001010001110011" => rgb <= "000000";
					when "11001010001110100" => rgb <= "000000";
					when "11001010001110101" => rgb <= "000000";
					when "11001010001110110" => rgb <= "000000";
					when "11001010001110111" => rgb <= "000000";
					when "11001010001111000" => rgb <= "000000";
					when "11001010001111001" => rgb <= "000000";
					when "11001010001111010" => rgb <= "000000";
					when "11001010001111011" => rgb <= "000000";
					when "11001010001111100" => rgb <= "000000";
					when "11001010001111101" => rgb <= "101010";
					when "11001010001111110" => rgb <= "101010";
					when "11001010001111111" => rgb <= "101010";
					when "11001010010000000" => rgb <= "111111";
					when "11001010010000001" => rgb <= "111111";
					when "11001010010000010" => rgb <= "101010";
					when "11001010010000011" => rgb <= "101010";
					when "11001010010000100" => rgb <= "101010";
					when "11001010010000101" => rgb <= "111111";
					when "11001010010000110" => rgb <= "111111";
					when "11001010010000111" => rgb <= "101010";
					when "11001010010001000" => rgb <= "101010";
					when "11001010010001001" => rgb <= "111111";
					when "11001010010001010" => rgb <= "101010";
					when "11001010010001011" => rgb <= "101010";
					when "11001010010001100" => rgb <= "000000";
					when "11001010010001101" => rgb <= "000000";
					when "11001010010001110" => rgb <= "000000";
					when "11001010010001111" => rgb <= "000000";
					when "11001010010010000" => rgb <= "000000";
					when "11001010010010001" => rgb <= "000000";
					when "11001010010010010" => rgb <= "000000";
					when "11001010010010011" => rgb <= "000000";
					when "11001010010010100" => rgb <= "000000";
					when "11001010010010101" => rgb <= "000000";
					when "11001010010010110" => rgb <= "000000";
					when "11001010010010111" => rgb <= "000000";
					when "11001010010011000" => rgb <= "000000";
					when "11001010010011001" => rgb <= "000000";
					when "11001010010011010" => rgb <= "000000";
					when "11001010010011011" => rgb <= "000000";
					when "11001010010011100" => rgb <= "000000";
					when "11001010010011101" => rgb <= "000000";
					when "11001010010011110" => rgb <= "000000";
					when "11001010010011111" => rgb <= "000000";
					when "11001010010100000" => rgb <= "000000";
					when "11001010010100001" => rgb <= "000000";
					when "11001010010100010" => rgb <= "010101";
					when "11001010010100011" => rgb <= "101010";
					when "11001010010100100" => rgb <= "111111";
					when "11001010010100101" => rgb <= "111111";
					when "11001010010100110" => rgb <= "101010";
					when "11001010010100111" => rgb <= "111111";
					when "11001010010101000" => rgb <= "101010";
					when "11001010010101001" => rgb <= "101010";
					when "11001010010101010" => rgb <= "000000";
					when "11001010010101011" => rgb <= "000000";
					when "11001010010101100" => rgb <= "000000";
					when "11001010010101101" => rgb <= "000000";
					when "11001010010101110" => rgb <= "000000";
					when "11001010010101111" => rgb <= "000000";
					when "11001010010110000" => rgb <= "000000";
					when "11001010010110001" => rgb <= "010101";
					when "11001010010110010" => rgb <= "111111";
					when "11001010010110011" => rgb <= "101010";
					when "11001010010110100" => rgb <= "111111";
					when "11001010010110101" => rgb <= "111111";
					when "11001010010110110" => rgb <= "101010";
					when "11001010010110111" => rgb <= "111111";
					when "11001010010111000" => rgb <= "101010";
					when "11001010010111001" => rgb <= "000000";
					when "11001010010111010" => rgb <= "000000";
					when "11001010010111011" => rgb <= "000000";
					when "11001010010111100" => rgb <= "000000";
					when "11001010010111101" => rgb <= "000000";
					when "11001010010111110" => rgb <= "000000";
					when "11001010010111111" => rgb <= "000000";
					when "11001010011000000" => rgb <= "010101";
					when "11001010011000001" => rgb <= "101010";
					when "11001010011000010" => rgb <= "111111";
					when "11001010011000011" => rgb <= "111111";
					when "11001010011000100" => rgb <= "101010";
					when "11001010011000101" => rgb <= "111111";
					when "11001010011000110" => rgb <= "101010";
					when "11001010011000111" => rgb <= "111111";
					when "11001010011001000" => rgb <= "101010";
					when "11001010011001001" => rgb <= "101010";
					when "11001010011001010" => rgb <= "111111";
					when "11001010011001011" => rgb <= "101010";
					when "11001010011001100" => rgb <= "111111";
					when "11001010011001101" => rgb <= "111111";
					when "11001010011001110" => rgb <= "111111";
					when "11001010011001111" => rgb <= "010101";
					when "11001010011010000" => rgb <= "000000";
					when "11001010011010001" => rgb <= "000000";
					when "11001010011010010" => rgb <= "000000";
					when "11001010011010011" => rgb <= "000000";
					when "11001010011010100" => rgb <= "000000";
					when "11001010011010101" => rgb <= "000000";
					when "11001010011010110" => rgb <= "000000";
					when "11001010011010111" => rgb <= "101010";
					when "11001010011011000" => rgb <= "101010";
					when "11001010011011001" => rgb <= "101010";
					when "11001010011011010" => rgb <= "101010";
					when "11001010011011011" => rgb <= "111111";
					when "11001010011011100" => rgb <= "111111";
					when "11001010011011101" => rgb <= "111111";
					when "11001010011011110" => rgb <= "111111";
					when "11001010011011111" => rgb <= "111111";
					when "11001010011100000" => rgb <= "111111";
					when "11001010011100001" => rgb <= "111111";
					when "11001010011100010" => rgb <= "111111";
					when "11001010011100011" => rgb <= "101010";
					when "11001010011100100" => rgb <= "111111";
					when "11001010011100101" => rgb <= "111111";
					when "11001010011100110" => rgb <= "000000";
					when "11001010011100111" => rgb <= "000000";
					when "11001010011101000" => rgb <= "000000";
					when "11001010011101001" => rgb <= "000000";
					when "11001010011101010" => rgb <= "000000";
					when "11001010011101011" => rgb <= "000000";
					when "11001010011101100" => rgb <= "000000";
					when "11001010011101101" => rgb <= "010101";
					when "11001010011101110" => rgb <= "111111";
					when "11001010011101111" => rgb <= "101010";
					when "11001010011110000" => rgb <= "111111";
					when "11001010011110001" => rgb <= "111111";
					when "11001010011110010" => rgb <= "111111";
					when "11001010011110011" => rgb <= "101010";
					when "11001010011110100" => rgb <= "101010";
					when "11001010011110101" => rgb <= "000000";
					when "11001010011110110" => rgb <= "000000";
					when "11001010011110111" => rgb <= "000000";
					when "11001010011111000" => rgb <= "000000";
					when "11001010011111001" => rgb <= "000000";
					when "11001010011111010" => rgb <= "000000";
					when "11001010011111011" => rgb <= "000000";
					when "11001010011111100" => rgb <= "000000";
					when "11001010011111101" => rgb <= "000000";
					when "11001010011111110" => rgb <= "000000";
					when "11001010011111111" => rgb <= "000000";
					when "11001010100000000" => rgb <= "000000";
					when "11001010100000001" => rgb <= "000000";
					when "11001010100000010" => rgb <= "000000";
					when "11001010100000011" => rgb <= "000000";
					when "11001010100000100" => rgb <= "000000";
					when "11001010100000101" => rgb <= "000000";
					when "11001010100000110" => rgb <= "000000";
					when "11001010100000111" => rgb <= "000000";
					when "11001010100001000" => rgb <= "000000";
					when "11001010100001001" => rgb <= "000000";
					when "11001010100001010" => rgb <= "000000";
					when "11001010100001011" => rgb <= "010101";
					when "11001010100001100" => rgb <= "111111";
					when "11001010100001101" => rgb <= "101010";
					when "11001010100001110" => rgb <= "111111";
					when "11001010100001111" => rgb <= "111111";
					when "11001010100010000" => rgb <= "111111";
					when "11001010100010001" => rgb <= "111111";
					when "11001010100010010" => rgb <= "111111";
					when "11001010100010011" => rgb <= "111111";
					when "11001010100010100" => rgb <= "111111";
					when "11001010100010101" => rgb <= "111111";
					when "11001010100010110" => rgb <= "111111";
					when "11001010100010111" => rgb <= "111111";
					when "11001010100011000" => rgb <= "101010";
					when "11001010100011001" => rgb <= "101010";
					when "11001010100011010" => rgb <= "101010";
					when "11001010100011011" => rgb <= "000000";
					when "11001010100011100" => rgb <= "000000";
					when "11001010100011101" => rgb <= "000000";
					when "11001010100011110" => rgb <= "000000";
					when "11001010100011111" => rgb <= "000000";
					when "11001010100100000" => rgb <= "000000";
					when "11001010100100001" => rgb <= "000000";
					when "11001010100100010" => rgb <= "000000";
					when "11001010100100011" => rgb <= "000000";
					when "11001010100100100" => rgb <= "000000";
					when "11001010100100101" => rgb <= "000000";
					when "11001010100100110" => rgb <= "000000";
					when "11001010100100111" => rgb <= "000000";
					when "11001010100101000" => rgb <= "000000";
					when "11001010100101001" => rgb <= "000000";
					when "11001010100101010" => rgb <= "000000";
					when "11001010100101011" => rgb <= "000000";
					when "11001010100101100" => rgb <= "000000";
					when "11001010100101101" => rgb <= "000000";
					when "11001010100101110" => rgb <= "000000";
					when "11001010100101111" => rgb <= "000000";
					when "11001010100110000" => rgb <= "000000";
					when "11001010100110001" => rgb <= "000000";
					when "11001010100110010" => rgb <= "000000";
					when "11001010100110011" => rgb <= "000000";
					when "11001010100110100" => rgb <= "000000";
					when "11001010100110101" => rgb <= "000000";
					when "11001010100110110" => rgb <= "000000";
					when "11001010100110111" => rgb <= "000000";
					when "11001010100111000" => rgb <= "000000";
					when "11001010100111001" => rgb <= "000000";
					when "11001010100111010" => rgb <= "000000";
					when "11001010100111011" => rgb <= "000000";
					when "11001010100111100" => rgb <= "000000";
					when "11001010100111101" => rgb <= "000000";
					when "11001010100111110" => rgb <= "000000";
					when "11001010100111111" => rgb <= "000000";
					when "11001011000000000" => rgb <= "000000";
					when "11001011000000001" => rgb <= "000000";
					when "11001011000000010" => rgb <= "000000";
					when "11001011000000011" => rgb <= "000000";
					when "11001011000000100" => rgb <= "000000";
					when "11001011000000101" => rgb <= "000000";
					when "11001011000000110" => rgb <= "000000";
					when "11001011000000111" => rgb <= "000000";
					when "11001011000001000" => rgb <= "000000";
					when "11001011000001001" => rgb <= "000000";
					when "11001011000001010" => rgb <= "000000";
					when "11001011000001011" => rgb <= "000000";
					when "11001011000001100" => rgb <= "000000";
					when "11001011000001101" => rgb <= "000000";
					when "11001011000001110" => rgb <= "000000";
					when "11001011000001111" => rgb <= "000000";
					when "11001011000010000" => rgb <= "000000";
					when "11001011000010001" => rgb <= "000000";
					when "11001011000010010" => rgb <= "000000";
					when "11001011000010011" => rgb <= "000000";
					when "11001011000010100" => rgb <= "101010";
					when "11001011000010101" => rgb <= "111111";
					when "11001011000010110" => rgb <= "101010";
					when "11001011000010111" => rgb <= "111111";
					when "11001011000011000" => rgb <= "111111";
					when "11001011000011001" => rgb <= "111111";
					when "11001011000011010" => rgb <= "111111";
					when "11001011000011011" => rgb <= "111111";
					when "11001011000011100" => rgb <= "111111";
					when "11001011000011101" => rgb <= "111111";
					when "11001011000011110" => rgb <= "111111";
					when "11001011000011111" => rgb <= "111111";
					when "11001011000100000" => rgb <= "111111";
					when "11001011000100001" => rgb <= "101010";
					when "11001011000100010" => rgb <= "111111";
					when "11001011000100011" => rgb <= "000000";
					when "11001011000100100" => rgb <= "000000";
					when "11001011000100101" => rgb <= "000000";
					when "11001011000100110" => rgb <= "000000";
					when "11001011000100111" => rgb <= "000000";
					when "11001011000101000" => rgb <= "000000";
					when "11001011000101001" => rgb <= "000000";
					when "11001011000101010" => rgb <= "000000";
					when "11001011000101011" => rgb <= "000000";
					when "11001011000101100" => rgb <= "000000";
					when "11001011000101101" => rgb <= "000000";
					when "11001011000101110" => rgb <= "000000";
					when "11001011000101111" => rgb <= "000000";
					when "11001011000110000" => rgb <= "000000";
					when "11001011000110001" => rgb <= "000000";
					when "11001011000110010" => rgb <= "000000";
					when "11001011000110011" => rgb <= "000000";
					when "11001011000110100" => rgb <= "000000";
					when "11001011000110101" => rgb <= "000000";
					when "11001011000110110" => rgb <= "000000";
					when "11001011000110111" => rgb <= "000000";
					when "11001011000111000" => rgb <= "000000";
					when "11001011000111001" => rgb <= "010101";
					when "11001011000111010" => rgb <= "111111";
					when "11001011000111011" => rgb <= "101010";
					when "11001011000111100" => rgb <= "101010";
					when "11001011000111101" => rgb <= "101010";
					when "11001011000111110" => rgb <= "101010";
					when "11001011000111111" => rgb <= "111111";
					when "11001011001000000" => rgb <= "101010";
					when "11001011001000001" => rgb <= "000000";
					when "11001011001000010" => rgb <= "000000";
					when "11001011001000011" => rgb <= "000000";
					when "11001011001000100" => rgb <= "000000";
					when "11001011001000101" => rgb <= "000000";
					when "11001011001000110" => rgb <= "000000";
					when "11001011001000111" => rgb <= "000000";
					when "11001011001001000" => rgb <= "000000";
					when "11001011001001001" => rgb <= "000000";
					when "11001011001001010" => rgb <= "000000";
					when "11001011001001011" => rgb <= "000000";
					when "11001011001001100" => rgb <= "000000";
					when "11001011001001101" => rgb <= "000000";
					when "11001011001001110" => rgb <= "000000";
					when "11001011001001111" => rgb <= "000000";
					when "11001011001010000" => rgb <= "101010";
					when "11001011001010001" => rgb <= "111111";
					when "11001011001010010" => rgb <= "101010";
					when "11001011001010011" => rgb <= "101010";
					when "11001011001010100" => rgb <= "111111";
					when "11001011001010101" => rgb <= "111111";
					when "11001011001010110" => rgb <= "101010";
					when "11001011001010111" => rgb <= "101010";
					when "11001011001011000" => rgb <= "101010";
					when "11001011001011001" => rgb <= "101010";
					when "11001011001011010" => rgb <= "111111";
					when "11001011001011011" => rgb <= "111111";
					when "11001011001011100" => rgb <= "111111";
					when "11001011001011101" => rgb <= "101010";
					when "11001011001011110" => rgb <= "101010";
					when "11001011001011111" => rgb <= "000000";
					when "11001011001100000" => rgb <= "000000";
					when "11001011001100001" => rgb <= "000000";
					when "11001011001100010" => rgb <= "000000";
					when "11001011001100011" => rgb <= "000000";
					when "11001011001100100" => rgb <= "000000";
					when "11001011001100101" => rgb <= "000000";
					when "11001011001100110" => rgb <= "010101";
					when "11001011001100111" => rgb <= "101010";
					when "11001011001101000" => rgb <= "101010";
					when "11001011001101001" => rgb <= "101010";
					when "11001011001101010" => rgb <= "101010";
					when "11001011001101011" => rgb <= "101010";
					when "11001011001101100" => rgb <= "111111";
					when "11001011001101101" => rgb <= "101010";
					when "11001011001101110" => rgb <= "000000";
					when "11001011001101111" => rgb <= "000000";
					when "11001011001110000" => rgb <= "000000";
					when "11001011001110001" => rgb <= "000000";
					when "11001011001110010" => rgb <= "000000";
					when "11001011001110011" => rgb <= "000000";
					when "11001011001110100" => rgb <= "000000";
					when "11001011001110101" => rgb <= "000000";
					when "11001011001110110" => rgb <= "000000";
					when "11001011001110111" => rgb <= "000000";
					when "11001011001111000" => rgb <= "000000";
					when "11001011001111001" => rgb <= "000000";
					when "11001011001111010" => rgb <= "000000";
					when "11001011001111011" => rgb <= "000000";
					when "11001011001111100" => rgb <= "000000";
					when "11001011001111101" => rgb <= "101010";
					when "11001011001111110" => rgb <= "111111";
					when "11001011001111111" => rgb <= "111111";
					when "11001011010000000" => rgb <= "101010";
					when "11001011010000001" => rgb <= "101010";
					when "11001011010000010" => rgb <= "101010";
					when "11001011010000011" => rgb <= "111111";
					when "11001011010000100" => rgb <= "111111";
					when "11001011010000101" => rgb <= "101010";
					when "11001011010000110" => rgb <= "101010";
					when "11001011010000111" => rgb <= "111111";
					when "11001011010001000" => rgb <= "101010";
					when "11001011010001001" => rgb <= "111111";
					when "11001011010001010" => rgb <= "101010";
					when "11001011010001011" => rgb <= "111111";
					when "11001011010001100" => rgb <= "000000";
					when "11001011010001101" => rgb <= "000000";
					when "11001011010001110" => rgb <= "000000";
					when "11001011010001111" => rgb <= "000000";
					when "11001011010010000" => rgb <= "000000";
					when "11001011010010001" => rgb <= "000000";
					when "11001011010010010" => rgb <= "000000";
					when "11001011010010011" => rgb <= "000000";
					when "11001011010010100" => rgb <= "000000";
					when "11001011010010101" => rgb <= "000000";
					when "11001011010010110" => rgb <= "000000";
					when "11001011010010111" => rgb <= "000000";
					when "11001011010011000" => rgb <= "000000";
					when "11001011010011001" => rgb <= "000000";
					when "11001011010011010" => rgb <= "000000";
					when "11001011010011011" => rgb <= "000000";
					when "11001011010011100" => rgb <= "000000";
					when "11001011010011101" => rgb <= "000000";
					when "11001011010011110" => rgb <= "000000";
					when "11001011010011111" => rgb <= "000000";
					when "11001011010100000" => rgb <= "000000";
					when "11001011010100001" => rgb <= "000000";
					when "11001011010100010" => rgb <= "010101";
					when "11001011010100011" => rgb <= "101010";
					when "11001011010100100" => rgb <= "101010";
					when "11001011010100101" => rgb <= "111111";
					when "11001011010100110" => rgb <= "111111";
					when "11001011010100111" => rgb <= "101010";
					when "11001011010101000" => rgb <= "111111";
					when "11001011010101001" => rgb <= "101010";
					when "11001011010101010" => rgb <= "000000";
					when "11001011010101011" => rgb <= "000000";
					when "11001011010101100" => rgb <= "000000";
					when "11001011010101101" => rgb <= "000000";
					when "11001011010101110" => rgb <= "000000";
					when "11001011010101111" => rgb <= "000000";
					when "11001011010110000" => rgb <= "000000";
					when "11001011010110001" => rgb <= "010101";
					when "11001011010110010" => rgb <= "101010";
					when "11001011010110011" => rgb <= "101010";
					when "11001011010110100" => rgb <= "101010";
					when "11001011010110101" => rgb <= "111111";
					when "11001011010110110" => rgb <= "111111";
					when "11001011010110111" => rgb <= "101010";
					when "11001011010111000" => rgb <= "101010";
					when "11001011010111001" => rgb <= "000000";
					when "11001011010111010" => rgb <= "000000";
					when "11001011010111011" => rgb <= "000000";
					when "11001011010111100" => rgb <= "000000";
					when "11001011010111101" => rgb <= "000000";
					when "11001011010111110" => rgb <= "000000";
					when "11001011010111111" => rgb <= "000000";
					when "11001011011000000" => rgb <= "010101";
					when "11001011011000001" => rgb <= "111111";
					when "11001011011000010" => rgb <= "101010";
					when "11001011011000011" => rgb <= "111111";
					when "11001011011000100" => rgb <= "101010";
					when "11001011011000101" => rgb <= "111111";
					when "11001011011000110" => rgb <= "101010";
					when "11001011011000111" => rgb <= "111111";
					when "11001011011001000" => rgb <= "111111";
					when "11001011011001001" => rgb <= "101010";
					when "11001011011001010" => rgb <= "101010";
					when "11001011011001011" => rgb <= "101010";
					when "11001011011001100" => rgb <= "101010";
					when "11001011011001101" => rgb <= "101010";
					when "11001011011001110" => rgb <= "101010";
					when "11001011011001111" => rgb <= "101010";
					when "11001011011010000" => rgb <= "000000";
					when "11001011011010001" => rgb <= "000000";
					when "11001011011010010" => rgb <= "000000";
					when "11001011011010011" => rgb <= "000000";
					when "11001011011010100" => rgb <= "000000";
					when "11001011011010101" => rgb <= "000000";
					when "11001011011010110" => rgb <= "000000";
					when "11001011011010111" => rgb <= "101010";
					when "11001011011011000" => rgb <= "101010";
					when "11001011011011001" => rgb <= "101010";
					when "11001011011011010" => rgb <= "101010";
					when "11001011011011011" => rgb <= "111111";
					when "11001011011011100" => rgb <= "111111";
					when "11001011011011101" => rgb <= "111111";
					when "11001011011011110" => rgb <= "111111";
					when "11001011011011111" => rgb <= "111111";
					when "11001011011100000" => rgb <= "111111";
					when "11001011011100001" => rgb <= "111111";
					when "11001011011100010" => rgb <= "111111";
					when "11001011011100011" => rgb <= "101010";
					when "11001011011100100" => rgb <= "111111";
					when "11001011011100101" => rgb <= "111111";
					when "11001011011100110" => rgb <= "000000";
					when "11001011011100111" => rgb <= "000000";
					when "11001011011101000" => rgb <= "000000";
					when "11001011011101001" => rgb <= "000000";
					when "11001011011101010" => rgb <= "000000";
					when "11001011011101011" => rgb <= "000000";
					when "11001011011101100" => rgb <= "000000";
					when "11001011011101101" => rgb <= "010101";
					when "11001011011101110" => rgb <= "111111";
					when "11001011011101111" => rgb <= "101010";
					when "11001011011110000" => rgb <= "111111";
					when "11001011011110001" => rgb <= "111111";
					when "11001011011110010" => rgb <= "111111";
					when "11001011011110011" => rgb <= "101010";
					when "11001011011110100" => rgb <= "101010";
					when "11001011011110101" => rgb <= "000000";
					when "11001011011110110" => rgb <= "000000";
					when "11001011011110111" => rgb <= "000000";
					when "11001011011111000" => rgb <= "000000";
					when "11001011011111001" => rgb <= "000000";
					when "11001011011111010" => rgb <= "000000";
					when "11001011011111011" => rgb <= "000000";
					when "11001011011111100" => rgb <= "000000";
					when "11001011011111101" => rgb <= "000000";
					when "11001011011111110" => rgb <= "000000";
					when "11001011011111111" => rgb <= "000000";
					when "11001011100000000" => rgb <= "000000";
					when "11001011100000001" => rgb <= "000000";
					when "11001011100000010" => rgb <= "000000";
					when "11001011100000011" => rgb <= "000000";
					when "11001011100000100" => rgb <= "000000";
					when "11001011100000101" => rgb <= "000000";
					when "11001011100000110" => rgb <= "000000";
					when "11001011100000111" => rgb <= "000000";
					when "11001011100001000" => rgb <= "000000";
					when "11001011100001001" => rgb <= "000000";
					when "11001011100001010" => rgb <= "000000";
					when "11001011100001011" => rgb <= "010101";
					when "11001011100001100" => rgb <= "111111";
					when "11001011100001101" => rgb <= "101010";
					when "11001011100001110" => rgb <= "111111";
					when "11001011100001111" => rgb <= "111111";
					when "11001011100010000" => rgb <= "111111";
					when "11001011100010001" => rgb <= "111111";
					when "11001011100010010" => rgb <= "111111";
					when "11001011100010011" => rgb <= "111111";
					when "11001011100010100" => rgb <= "111111";
					when "11001011100010101" => rgb <= "111111";
					when "11001011100010110" => rgb <= "111111";
					when "11001011100010111" => rgb <= "111111";
					when "11001011100011000" => rgb <= "101010";
					when "11001011100011001" => rgb <= "101010";
					when "11001011100011010" => rgb <= "101010";
					when "11001011100011011" => rgb <= "000000";
					when "11001011100011100" => rgb <= "000000";
					when "11001011100011101" => rgb <= "000000";
					when "11001011100011110" => rgb <= "000000";
					when "11001011100011111" => rgb <= "000000";
					when "11001011100100000" => rgb <= "000000";
					when "11001011100100001" => rgb <= "000000";
					when "11001011100100010" => rgb <= "000000";
					when "11001011100100011" => rgb <= "000000";
					when "11001011100100100" => rgb <= "000000";
					when "11001011100100101" => rgb <= "000000";
					when "11001011100100110" => rgb <= "000000";
					when "11001011100100111" => rgb <= "000000";
					when "11001011100101000" => rgb <= "000000";
					when "11001011100101001" => rgb <= "000000";
					when "11001011100101010" => rgb <= "000000";
					when "11001011100101011" => rgb <= "000000";
					when "11001011100101100" => rgb <= "000000";
					when "11001011100101101" => rgb <= "000000";
					when "11001011100101110" => rgb <= "000000";
					when "11001011100101111" => rgb <= "000000";
					when "11001011100110000" => rgb <= "000000";
					when "11001011100110001" => rgb <= "000000";
					when "11001011100110010" => rgb <= "000000";
					when "11001011100110011" => rgb <= "000000";
					when "11001011100110100" => rgb <= "000000";
					when "11001011100110101" => rgb <= "000000";
					when "11001011100110110" => rgb <= "000000";
					when "11001011100110111" => rgb <= "000000";
					when "11001011100111000" => rgb <= "000000";
					when "11001011100111001" => rgb <= "000000";
					when "11001011100111010" => rgb <= "000000";
					when "11001011100111011" => rgb <= "000000";
					when "11001011100111100" => rgb <= "000000";
					when "11001011100111101" => rgb <= "000000";
					when "11001011100111110" => rgb <= "000000";
					when "11001011100111111" => rgb <= "000000";
					when "11001100000000000" => rgb <= "000000";
					when "11001100000000001" => rgb <= "000000";
					when "11001100000000010" => rgb <= "000000";
					when "11001100000000011" => rgb <= "000000";
					when "11001100000000100" => rgb <= "000000";
					when "11001100000000101" => rgb <= "000000";
					when "11001100000000110" => rgb <= "000000";
					when "11001100000000111" => rgb <= "000000";
					when "11001100000001000" => rgb <= "000000";
					when "11001100000001001" => rgb <= "000000";
					when "11001100000001010" => rgb <= "000000";
					when "11001100000001011" => rgb <= "000000";
					when "11001100000001100" => rgb <= "000000";
					when "11001100000001101" => rgb <= "000000";
					when "11001100000001110" => rgb <= "000000";
					when "11001100000001111" => rgb <= "000000";
					when "11001100000010000" => rgb <= "000000";
					when "11001100000010001" => rgb <= "000000";
					when "11001100000010010" => rgb <= "000000";
					when "11001100000010011" => rgb <= "000000";
					when "11001100000010100" => rgb <= "101010";
					when "11001100000010101" => rgb <= "111111";
					when "11001100000010110" => rgb <= "101010";
					when "11001100000010111" => rgb <= "111111";
					when "11001100000011000" => rgb <= "111111";
					when "11001100000011001" => rgb <= "111111";
					when "11001100000011010" => rgb <= "111111";
					when "11001100000011011" => rgb <= "111111";
					when "11001100000011100" => rgb <= "111111";
					when "11001100000011101" => rgb <= "111111";
					when "11001100000011110" => rgb <= "111111";
					when "11001100000011111" => rgb <= "111111";
					when "11001100000100000" => rgb <= "111111";
					when "11001100000100001" => rgb <= "101010";
					when "11001100000100010" => rgb <= "111111";
					when "11001100000100011" => rgb <= "000000";
					when "11001100000100100" => rgb <= "000000";
					when "11001100000100101" => rgb <= "000000";
					when "11001100000100110" => rgb <= "000000";
					when "11001100000100111" => rgb <= "000000";
					when "11001100000101000" => rgb <= "000000";
					when "11001100000101001" => rgb <= "000000";
					when "11001100000101010" => rgb <= "000000";
					when "11001100000101011" => rgb <= "000000";
					when "11001100000101100" => rgb <= "000000";
					when "11001100000101101" => rgb <= "000000";
					when "11001100000101110" => rgb <= "000000";
					when "11001100000101111" => rgb <= "000000";
					when "11001100000110000" => rgb <= "000000";
					when "11001100000110001" => rgb <= "000000";
					when "11001100000110010" => rgb <= "000000";
					when "11001100000110011" => rgb <= "000000";
					when "11001100000110100" => rgb <= "000000";
					when "11001100000110101" => rgb <= "000000";
					when "11001100000110110" => rgb <= "000000";
					when "11001100000110111" => rgb <= "000000";
					when "11001100000111000" => rgb <= "000000";
					when "11001100000111001" => rgb <= "010101";
					when "11001100000111010" => rgb <= "111111";
					when "11001100000111011" => rgb <= "101010";
					when "11001100000111100" => rgb <= "111111";
					when "11001100000111101" => rgb <= "111111";
					when "11001100000111110" => rgb <= "111111";
					when "11001100000111111" => rgb <= "111111";
					when "11001100001000000" => rgb <= "111111";
					when "11001100001000001" => rgb <= "000000";
					when "11001100001000010" => rgb <= "000000";
					when "11001100001000011" => rgb <= "000000";
					when "11001100001000100" => rgb <= "000000";
					when "11001100001000101" => rgb <= "000000";
					when "11001100001000110" => rgb <= "000000";
					when "11001100001000111" => rgb <= "000000";
					when "11001100001001000" => rgb <= "000000";
					when "11001100001001001" => rgb <= "000000";
					when "11001100001001010" => rgb <= "000000";
					when "11001100001001011" => rgb <= "000000";
					when "11001100001001100" => rgb <= "000000";
					when "11001100001001101" => rgb <= "000000";
					when "11001100001001110" => rgb <= "000000";
					when "11001100001001111" => rgb <= "000000";
					when "11001100001010000" => rgb <= "101010";
					when "11001100001010001" => rgb <= "111111";
					when "11001100001010010" => rgb <= "101010";
					when "11001100001010011" => rgb <= "111111";
					when "11001100001010100" => rgb <= "111111";
					when "11001100001010101" => rgb <= "111111";
					when "11001100001010110" => rgb <= "111111";
					when "11001100001010111" => rgb <= "111111";
					when "11001100001011000" => rgb <= "111111";
					when "11001100001011001" => rgb <= "111111";
					when "11001100001011010" => rgb <= "101010";
					when "11001100001011011" => rgb <= "101010";
					when "11001100001011100" => rgb <= "101010";
					when "11001100001011101" => rgb <= "111111";
					when "11001100001011110" => rgb <= "111111";
					when "11001100001011111" => rgb <= "000000";
					when "11001100001100000" => rgb <= "000000";
					when "11001100001100001" => rgb <= "000000";
					when "11001100001100010" => rgb <= "000000";
					when "11001100001100011" => rgb <= "000000";
					when "11001100001100100" => rgb <= "000000";
					when "11001100001100101" => rgb <= "000000";
					when "11001100001100110" => rgb <= "010101";
					when "11001100001100111" => rgb <= "111111";
					when "11001100001101000" => rgb <= "111111";
					when "11001100001101001" => rgb <= "111111";
					when "11001100001101010" => rgb <= "111111";
					when "11001100001101011" => rgb <= "111111";
					when "11001100001101100" => rgb <= "101010";
					when "11001100001101101" => rgb <= "111111";
					when "11001100001101110" => rgb <= "000000";
					when "11001100001101111" => rgb <= "000000";
					when "11001100001110000" => rgb <= "000000";
					when "11001100001110001" => rgb <= "000000";
					when "11001100001110010" => rgb <= "000000";
					when "11001100001110011" => rgb <= "000000";
					when "11001100001110100" => rgb <= "000000";
					when "11001100001110101" => rgb <= "000000";
					when "11001100001110110" => rgb <= "000000";
					when "11001100001110111" => rgb <= "000000";
					when "11001100001111000" => rgb <= "000000";
					when "11001100001111001" => rgb <= "000000";
					when "11001100001111010" => rgb <= "000000";
					when "11001100001111011" => rgb <= "000000";
					when "11001100001111100" => rgb <= "000000";
					when "11001100001111101" => rgb <= "101010";
					when "11001100001111110" => rgb <= "111111";
					when "11001100001111111" => rgb <= "101010";
					when "11001100010000000" => rgb <= "111111";
					when "11001100010000001" => rgb <= "111111";
					when "11001100010000010" => rgb <= "111111";
					when "11001100010000011" => rgb <= "101010";
					when "11001100010000100" => rgb <= "101010";
					when "11001100010000101" => rgb <= "111111";
					when "11001100010000110" => rgb <= "111111";
					when "11001100010000111" => rgb <= "111111";
					when "11001100010001000" => rgb <= "111111";
					when "11001100010001001" => rgb <= "111111";
					when "11001100010001010" => rgb <= "101010";
					when "11001100010001011" => rgb <= "111111";
					when "11001100010001100" => rgb <= "000000";
					when "11001100010001101" => rgb <= "000000";
					when "11001100010001110" => rgb <= "000000";
					when "11001100010001111" => rgb <= "000000";
					when "11001100010010000" => rgb <= "000000";
					when "11001100010010001" => rgb <= "000000";
					when "11001100010010010" => rgb <= "000000";
					when "11001100010010011" => rgb <= "000000";
					when "11001100010010100" => rgb <= "000000";
					when "11001100010010101" => rgb <= "000000";
					when "11001100010010110" => rgb <= "000000";
					when "11001100010010111" => rgb <= "000000";
					when "11001100010011000" => rgb <= "000000";
					when "11001100010011001" => rgb <= "000000";
					when "11001100010011010" => rgb <= "000000";
					when "11001100010011011" => rgb <= "000000";
					when "11001100010011100" => rgb <= "000000";
					when "11001100010011101" => rgb <= "000000";
					when "11001100010011110" => rgb <= "000000";
					when "11001100010011111" => rgb <= "000000";
					when "11001100010100000" => rgb <= "000000";
					when "11001100010100001" => rgb <= "000000";
					when "11001100010100010" => rgb <= "010101";
					when "11001100010100011" => rgb <= "111111";
					when "11001100010100100" => rgb <= "101010";
					when "11001100010100101" => rgb <= "111111";
					when "11001100010100110" => rgb <= "101010";
					when "11001100010100111" => rgb <= "111111";
					when "11001100010101000" => rgb <= "111111";
					when "11001100010101001" => rgb <= "111111";
					when "11001100010101010" => rgb <= "000000";
					when "11001100010101011" => rgb <= "000000";
					when "11001100010101100" => rgb <= "000000";
					when "11001100010101101" => rgb <= "000000";
					when "11001100010101110" => rgb <= "000000";
					when "11001100010101111" => rgb <= "000000";
					when "11001100010110000" => rgb <= "000000";
					when "11001100010110001" => rgb <= "010101";
					when "11001100010110010" => rgb <= "101010";
					when "11001100010110011" => rgb <= "111111";
					when "11001100010110100" => rgb <= "111111";
					when "11001100010110101" => rgb <= "101010";
					when "11001100010110110" => rgb <= "111111";
					when "11001100010110111" => rgb <= "111111";
					when "11001100010111000" => rgb <= "101010";
					when "11001100010111001" => rgb <= "000000";
					when "11001100010111010" => rgb <= "000000";
					when "11001100010111011" => rgb <= "000000";
					when "11001100010111100" => rgb <= "000000";
					when "11001100010111101" => rgb <= "000000";
					when "11001100010111110" => rgb <= "000000";
					when "11001100010111111" => rgb <= "000000";
					when "11001100011000000" => rgb <= "010101";
					when "11001100011000001" => rgb <= "101010";
					when "11001100011000010" => rgb <= "101010";
					when "11001100011000011" => rgb <= "101010";
					when "11001100011000100" => rgb <= "101010";
					when "11001100011000101" => rgb <= "111111";
					when "11001100011000110" => rgb <= "111111";
					when "11001100011000111" => rgb <= "101010";
					when "11001100011001000" => rgb <= "111111";
					when "11001100011001001" => rgb <= "111111";
					when "11001100011001010" => rgb <= "111111";
					when "11001100011001011" => rgb <= "111111";
					when "11001100011001100" => rgb <= "111111";
					when "11001100011001101" => rgb <= "111111";
					when "11001100011001110" => rgb <= "111111";
					when "11001100011001111" => rgb <= "010101";
					when "11001100011010000" => rgb <= "000000";
					when "11001100011010001" => rgb <= "000000";
					when "11001100011010010" => rgb <= "000000";
					when "11001100011010011" => rgb <= "000000";
					when "11001100011010100" => rgb <= "000000";
					when "11001100011010101" => rgb <= "000000";
					when "11001100011010110" => rgb <= "000000";
					when "11001100011010111" => rgb <= "101010";
					when "11001100011011000" => rgb <= "101010";
					when "11001100011011001" => rgb <= "101010";
					when "11001100011011010" => rgb <= "101010";
					when "11001100011011011" => rgb <= "111111";
					when "11001100011011100" => rgb <= "111111";
					when "11001100011011101" => rgb <= "111111";
					when "11001100011011110" => rgb <= "111111";
					when "11001100011011111" => rgb <= "111111";
					when "11001100011100000" => rgb <= "111111";
					when "11001100011100001" => rgb <= "111111";
					when "11001100011100010" => rgb <= "111111";
					when "11001100011100011" => rgb <= "101010";
					when "11001100011100100" => rgb <= "111111";
					when "11001100011100101" => rgb <= "111111";
					when "11001100011100110" => rgb <= "000000";
					when "11001100011100111" => rgb <= "000000";
					when "11001100011101000" => rgb <= "000000";
					when "11001100011101001" => rgb <= "000000";
					when "11001100011101010" => rgb <= "000000";
					when "11001100011101011" => rgb <= "000000";
					when "11001100011101100" => rgb <= "000000";
					when "11001100011101101" => rgb <= "010101";
					when "11001100011101110" => rgb <= "111111";
					when "11001100011101111" => rgb <= "101010";
					when "11001100011110000" => rgb <= "111111";
					when "11001100011110001" => rgb <= "111111";
					when "11001100011110010" => rgb <= "111111";
					when "11001100011110011" => rgb <= "101010";
					when "11001100011110100" => rgb <= "101010";
					when "11001100011110101" => rgb <= "000000";
					when "11001100011110110" => rgb <= "000000";
					when "11001100011110111" => rgb <= "000000";
					when "11001100011111000" => rgb <= "000000";
					when "11001100011111001" => rgb <= "000000";
					when "11001100011111010" => rgb <= "000000";
					when "11001100011111011" => rgb <= "000000";
					when "11001100011111100" => rgb <= "000000";
					when "11001100011111101" => rgb <= "000000";
					when "11001100011111110" => rgb <= "000000";
					when "11001100011111111" => rgb <= "000000";
					when "11001100100000000" => rgb <= "000000";
					when "11001100100000001" => rgb <= "000000";
					when "11001100100000010" => rgb <= "000000";
					when "11001100100000011" => rgb <= "000000";
					when "11001100100000100" => rgb <= "000000";
					when "11001100100000101" => rgb <= "000000";
					when "11001100100000110" => rgb <= "000000";
					when "11001100100000111" => rgb <= "000000";
					when "11001100100001000" => rgb <= "000000";
					when "11001100100001001" => rgb <= "000000";
					when "11001100100001010" => rgb <= "000000";
					when "11001100100001011" => rgb <= "010101";
					when "11001100100001100" => rgb <= "111111";
					when "11001100100001101" => rgb <= "101010";
					when "11001100100001110" => rgb <= "111111";
					when "11001100100001111" => rgb <= "111111";
					when "11001100100010000" => rgb <= "111111";
					when "11001100100010001" => rgb <= "111111";
					when "11001100100010010" => rgb <= "111111";
					when "11001100100010011" => rgb <= "111111";
					when "11001100100010100" => rgb <= "111111";
					when "11001100100010101" => rgb <= "111111";
					when "11001100100010110" => rgb <= "111111";
					when "11001100100010111" => rgb <= "111111";
					when "11001100100011000" => rgb <= "101010";
					when "11001100100011001" => rgb <= "101010";
					when "11001100100011010" => rgb <= "101010";
					when "11001100100011011" => rgb <= "000000";
					when "11001100100011100" => rgb <= "000000";
					when "11001100100011101" => rgb <= "000000";
					when "11001100100011110" => rgb <= "000000";
					when "11001100100011111" => rgb <= "000000";
					when "11001100100100000" => rgb <= "000000";
					when "11001100100100001" => rgb <= "000000";
					when "11001100100100010" => rgb <= "000000";
					when "11001100100100011" => rgb <= "000000";
					when "11001100100100100" => rgb <= "000000";
					when "11001100100100101" => rgb <= "000000";
					when "11001100100100110" => rgb <= "000000";
					when "11001100100100111" => rgb <= "000000";
					when "11001100100101000" => rgb <= "000000";
					when "11001100100101001" => rgb <= "000000";
					when "11001100100101010" => rgb <= "000000";
					when "11001100100101011" => rgb <= "000000";
					when "11001100100101100" => rgb <= "000000";
					when "11001100100101101" => rgb <= "000000";
					when "11001100100101110" => rgb <= "000000";
					when "11001100100101111" => rgb <= "000000";
					when "11001100100110000" => rgb <= "000000";
					when "11001100100110001" => rgb <= "000000";
					when "11001100100110010" => rgb <= "000000";
					when "11001100100110011" => rgb <= "000000";
					when "11001100100110100" => rgb <= "000000";
					when "11001100100110101" => rgb <= "000000";
					when "11001100100110110" => rgb <= "000000";
					when "11001100100110111" => rgb <= "000000";
					when "11001100100111000" => rgb <= "000000";
					when "11001100100111001" => rgb <= "000000";
					when "11001100100111010" => rgb <= "000000";
					when "11001100100111011" => rgb <= "000000";
					when "11001100100111100" => rgb <= "000000";
					when "11001100100111101" => rgb <= "000000";
					when "11001100100111110" => rgb <= "000000";
					when "11001100100111111" => rgb <= "000000";
					when "11001101000000000" => rgb <= "000000";
					when "11001101000000001" => rgb <= "000000";
					when "11001101000000010" => rgb <= "000000";
					when "11001101000000011" => rgb <= "000000";
					when "11001101000000100" => rgb <= "000000";
					when "11001101000000101" => rgb <= "000000";
					when "11001101000000110" => rgb <= "000000";
					when "11001101000000111" => rgb <= "000000";
					when "11001101000001000" => rgb <= "000000";
					when "11001101000001001" => rgb <= "000000";
					when "11001101000001010" => rgb <= "000000";
					when "11001101000001011" => rgb <= "000000";
					when "11001101000001100" => rgb <= "000000";
					when "11001101000001101" => rgb <= "000000";
					when "11001101000001110" => rgb <= "000000";
					when "11001101000001111" => rgb <= "000000";
					when "11001101000010000" => rgb <= "000000";
					when "11001101000010001" => rgb <= "000000";
					when "11001101000010010" => rgb <= "000000";
					when "11001101000010011" => rgb <= "000000";
					when "11001101000010100" => rgb <= "101010";
					when "11001101000010101" => rgb <= "111111";
					when "11001101000010110" => rgb <= "101010";
					when "11001101000010111" => rgb <= "111111";
					when "11001101000011000" => rgb <= "111111";
					when "11001101000011001" => rgb <= "111111";
					when "11001101000011010" => rgb <= "111111";
					when "11001101000011011" => rgb <= "111111";
					when "11001101000011100" => rgb <= "111111";
					when "11001101000011101" => rgb <= "111111";
					when "11001101000011110" => rgb <= "111111";
					when "11001101000011111" => rgb <= "111111";
					when "11001101000100000" => rgb <= "111111";
					when "11001101000100001" => rgb <= "101010";
					when "11001101000100010" => rgb <= "111111";
					when "11001101000100011" => rgb <= "000000";
					when "11001101000100100" => rgb <= "000000";
					when "11001101000100101" => rgb <= "000000";
					when "11001101000100110" => rgb <= "000000";
					when "11001101000100111" => rgb <= "000000";
					when "11001101000101000" => rgb <= "000000";
					when "11001101000101001" => rgb <= "000000";
					when "11001101000101010" => rgb <= "000000";
					when "11001101000101011" => rgb <= "000000";
					when "11001101000101100" => rgb <= "000000";
					when "11001101000101101" => rgb <= "000000";
					when "11001101000101110" => rgb <= "000000";
					when "11001101000101111" => rgb <= "000000";
					when "11001101000110000" => rgb <= "000000";
					when "11001101000110001" => rgb <= "000000";
					when "11001101000110010" => rgb <= "000000";
					when "11001101000110011" => rgb <= "000000";
					when "11001101000110100" => rgb <= "000000";
					when "11001101000110101" => rgb <= "000000";
					when "11001101000110110" => rgb <= "000000";
					when "11001101000110111" => rgb <= "000000";
					when "11001101000111000" => rgb <= "000000";
					when "11001101000111001" => rgb <= "010101";
					when "11001101000111010" => rgb <= "101010";
					when "11001101000111011" => rgb <= "101010";
					when "11001101000111100" => rgb <= "101010";
					when "11001101000111101" => rgb <= "101010";
					when "11001101000111110" => rgb <= "101010";
					when "11001101000111111" => rgb <= "101010";
					when "11001101001000000" => rgb <= "101010";
					when "11001101001000001" => rgb <= "000000";
					when "11001101001000010" => rgb <= "000000";
					when "11001101001000011" => rgb <= "000000";
					when "11001101001000100" => rgb <= "000000";
					when "11001101001000101" => rgb <= "000000";
					when "11001101001000110" => rgb <= "000000";
					when "11001101001000111" => rgb <= "000000";
					when "11001101001001000" => rgb <= "000000";
					when "11001101001001001" => rgb <= "000000";
					when "11001101001001010" => rgb <= "000000";
					when "11001101001001011" => rgb <= "000000";
					when "11001101001001100" => rgb <= "000000";
					when "11001101001001101" => rgb <= "000000";
					when "11001101001001110" => rgb <= "000000";
					when "11001101001001111" => rgb <= "000000";
					when "11001101001010000" => rgb <= "101010";
					when "11001101001010001" => rgb <= "101010";
					when "11001101001010010" => rgb <= "101010";
					when "11001101001010011" => rgb <= "111111";
					when "11001101001010100" => rgb <= "111111";
					when "11001101001010101" => rgb <= "101010";
					when "11001101001010110" => rgb <= "111111";
					when "11001101001010111" => rgb <= "101010";
					when "11001101001011000" => rgb <= "101010";
					when "11001101001011001" => rgb <= "101010";
					when "11001101001011010" => rgb <= "101010";
					when "11001101001011011" => rgb <= "101010";
					when "11001101001011100" => rgb <= "101010";
					when "11001101001011101" => rgb <= "101010";
					when "11001101001011110" => rgb <= "101010";
					when "11001101001011111" => rgb <= "000000";
					when "11001101001100000" => rgb <= "000000";
					when "11001101001100001" => rgb <= "000000";
					when "11001101001100010" => rgb <= "000000";
					when "11001101001100011" => rgb <= "000000";
					when "11001101001100100" => rgb <= "000000";
					when "11001101001100101" => rgb <= "000000";
					when "11001101001100110" => rgb <= "010101";
					when "11001101001100111" => rgb <= "101010";
					when "11001101001101000" => rgb <= "101010";
					when "11001101001101001" => rgb <= "101010";
					when "11001101001101010" => rgb <= "101010";
					when "11001101001101011" => rgb <= "101010";
					when "11001101001101100" => rgb <= "101010";
					when "11001101001101101" => rgb <= "101010";
					when "11001101001101110" => rgb <= "000000";
					when "11001101001101111" => rgb <= "000000";
					when "11001101001110000" => rgb <= "000000";
					when "11001101001110001" => rgb <= "000000";
					when "11001101001110010" => rgb <= "000000";
					when "11001101001110011" => rgb <= "000000";
					when "11001101001110100" => rgb <= "000000";
					when "11001101001110101" => rgb <= "000000";
					when "11001101001110110" => rgb <= "000000";
					when "11001101001110111" => rgb <= "000000";
					when "11001101001111000" => rgb <= "000000";
					when "11001101001111001" => rgb <= "000000";
					when "11001101001111010" => rgb <= "000000";
					when "11001101001111011" => rgb <= "000000";
					when "11001101001111100" => rgb <= "000000";
					when "11001101001111101" => rgb <= "101010";
					when "11001101001111110" => rgb <= "111111";
					when "11001101001111111" => rgb <= "111111";
					when "11001101010000000" => rgb <= "101010";
					when "11001101010000001" => rgb <= "101010";
					when "11001101010000010" => rgb <= "111111";
					when "11001101010000011" => rgb <= "101010";
					when "11001101010000100" => rgb <= "101010";
					when "11001101010000101" => rgb <= "101010";
					when "11001101010000110" => rgb <= "101010";
					when "11001101010000111" => rgb <= "101010";
					when "11001101010001000" => rgb <= "101010";
					when "11001101010001001" => rgb <= "101010";
					when "11001101010001010" => rgb <= "101010";
					when "11001101010001011" => rgb <= "101010";
					when "11001101010001100" => rgb <= "000000";
					when "11001101010001101" => rgb <= "000000";
					when "11001101010001110" => rgb <= "000000";
					when "11001101010001111" => rgb <= "000000";
					when "11001101010010000" => rgb <= "000000";
					when "11001101010010001" => rgb <= "000000";
					when "11001101010010010" => rgb <= "000000";
					when "11001101010010011" => rgb <= "000000";
					when "11001101010010100" => rgb <= "000000";
					when "11001101010010101" => rgb <= "000000";
					when "11001101010010110" => rgb <= "000000";
					when "11001101010010111" => rgb <= "000000";
					when "11001101010011000" => rgb <= "000000";
					when "11001101010011001" => rgb <= "000000";
					when "11001101010011010" => rgb <= "000000";
					when "11001101010011011" => rgb <= "000000";
					when "11001101010011100" => rgb <= "000000";
					when "11001101010011101" => rgb <= "000000";
					when "11001101010011110" => rgb <= "000000";
					when "11001101010011111" => rgb <= "000000";
					when "11001101010100000" => rgb <= "000000";
					when "11001101010100001" => rgb <= "000000";
					when "11001101010100010" => rgb <= "010101";
					when "11001101010100011" => rgb <= "101010";
					when "11001101010100100" => rgb <= "101010";
					when "11001101010100101" => rgb <= "101010";
					when "11001101010100110" => rgb <= "101010";
					when "11001101010100111" => rgb <= "101010";
					when "11001101010101000" => rgb <= "101010";
					when "11001101010101001" => rgb <= "101010";
					when "11001101010101010" => rgb <= "000000";
					when "11001101010101011" => rgb <= "000000";
					when "11001101010101100" => rgb <= "000000";
					when "11001101010101101" => rgb <= "000000";
					when "11001101010101110" => rgb <= "000000";
					when "11001101010101111" => rgb <= "000000";
					when "11001101010110000" => rgb <= "000000";
					when "11001101010110001" => rgb <= "010101";
					when "11001101010110010" => rgb <= "101010";
					when "11001101010110011" => rgb <= "101010";
					when "11001101010110100" => rgb <= "101010";
					when "11001101010110101" => rgb <= "101010";
					when "11001101010110110" => rgb <= "101010";
					when "11001101010110111" => rgb <= "101010";
					when "11001101010111000" => rgb <= "101010";
					when "11001101010111001" => rgb <= "000000";
					when "11001101010111010" => rgb <= "000000";
					when "11001101010111011" => rgb <= "000000";
					when "11001101010111100" => rgb <= "000000";
					when "11001101010111101" => rgb <= "000000";
					when "11001101010111110" => rgb <= "000000";
					when "11001101010111111" => rgb <= "000000";
					when "11001101011000000" => rgb <= "010101";
					when "11001101011000001" => rgb <= "101010";
					when "11001101011000010" => rgb <= "101010";
					when "11001101011000011" => rgb <= "111111";
					when "11001101011000100" => rgb <= "111111";
					when "11001101011000101" => rgb <= "101010";
					when "11001101011000110" => rgb <= "101010";
					when "11001101011000111" => rgb <= "111111";
					when "11001101011001000" => rgb <= "101010";
					when "11001101011001001" => rgb <= "101010";
					when "11001101011001010" => rgb <= "101010";
					when "11001101011001011" => rgb <= "101010";
					when "11001101011001100" => rgb <= "101010";
					when "11001101011001101" => rgb <= "101010";
					when "11001101011001110" => rgb <= "101010";
					when "11001101011001111" => rgb <= "010101";
					when "11001101011010000" => rgb <= "000000";
					when "11001101011010001" => rgb <= "000000";
					when "11001101011010010" => rgb <= "000000";
					when "11001101011010011" => rgb <= "000000";
					when "11001101011010100" => rgb <= "000000";
					when "11001101011010101" => rgb <= "000000";
					when "11001101011010110" => rgb <= "000000";
					when "11001101011010111" => rgb <= "101010";
					when "11001101011011000" => rgb <= "101010";
					when "11001101011011001" => rgb <= "101010";
					when "11001101011011010" => rgb <= "101010";
					when "11001101011011011" => rgb <= "111111";
					when "11001101011011100" => rgb <= "111111";
					when "11001101011011101" => rgb <= "111111";
					when "11001101011011110" => rgb <= "111111";
					when "11001101011011111" => rgb <= "111111";
					when "11001101011100000" => rgb <= "111111";
					when "11001101011100001" => rgb <= "111111";
					when "11001101011100010" => rgb <= "111111";
					when "11001101011100011" => rgb <= "101010";
					when "11001101011100100" => rgb <= "111111";
					when "11001101011100101" => rgb <= "111111";
					when "11001101011100110" => rgb <= "000000";
					when "11001101011100111" => rgb <= "000000";
					when "11001101011101000" => rgb <= "000000";
					when "11001101011101001" => rgb <= "000000";
					when "11001101011101010" => rgb <= "000000";
					when "11001101011101011" => rgb <= "000000";
					when "11001101011101100" => rgb <= "000000";
					when "11001101011101101" => rgb <= "010101";
					when "11001101011101110" => rgb <= "111111";
					when "11001101011101111" => rgb <= "101010";
					when "11001101011110000" => rgb <= "111111";
					when "11001101011110001" => rgb <= "111111";
					when "11001101011110010" => rgb <= "111111";
					when "11001101011110011" => rgb <= "101010";
					when "11001101011110100" => rgb <= "101010";
					when "11001101011110101" => rgb <= "000000";
					when "11001101011110110" => rgb <= "000000";
					when "11001101011110111" => rgb <= "000000";
					when "11001101011111000" => rgb <= "000000";
					when "11001101011111001" => rgb <= "000000";
					when "11001101011111010" => rgb <= "000000";
					when "11001101011111011" => rgb <= "000000";
					when "11001101011111100" => rgb <= "000000";
					when "11001101011111101" => rgb <= "000000";
					when "11001101011111110" => rgb <= "000000";
					when "11001101011111111" => rgb <= "000000";
					when "11001101100000000" => rgb <= "000000";
					when "11001101100000001" => rgb <= "000000";
					when "11001101100000010" => rgb <= "000000";
					when "11001101100000011" => rgb <= "000000";
					when "11001101100000100" => rgb <= "000000";
					when "11001101100000101" => rgb <= "000000";
					when "11001101100000110" => rgb <= "000000";
					when "11001101100000111" => rgb <= "000000";
					when "11001101100001000" => rgb <= "000000";
					when "11001101100001001" => rgb <= "000000";
					when "11001101100001010" => rgb <= "000000";
					when "11001101100001011" => rgb <= "010101";
					when "11001101100001100" => rgb <= "111111";
					when "11001101100001101" => rgb <= "101010";
					when "11001101100001110" => rgb <= "111111";
					when "11001101100001111" => rgb <= "111111";
					when "11001101100010000" => rgb <= "111111";
					when "11001101100010001" => rgb <= "111111";
					when "11001101100010010" => rgb <= "111111";
					when "11001101100010011" => rgb <= "111111";
					when "11001101100010100" => rgb <= "111111";
					when "11001101100010101" => rgb <= "111111";
					when "11001101100010110" => rgb <= "111111";
					when "11001101100010111" => rgb <= "111111";
					when "11001101100011000" => rgb <= "101010";
					when "11001101100011001" => rgb <= "101010";
					when "11001101100011010" => rgb <= "101010";
					when "11001101100011011" => rgb <= "000000";
					when "11001101100011100" => rgb <= "000000";
					when "11001101100011101" => rgb <= "000000";
					when "11001101100011110" => rgb <= "000000";
					when "11001101100011111" => rgb <= "000000";
					when "11001101100100000" => rgb <= "000000";
					when "11001101100100001" => rgb <= "000000";
					when "11001101100100010" => rgb <= "000000";
					when "11001101100100011" => rgb <= "000000";
					when "11001101100100100" => rgb <= "000000";
					when "11001101100100101" => rgb <= "000000";
					when "11001101100100110" => rgb <= "000000";
					when "11001101100100111" => rgb <= "000000";
					when "11001101100101000" => rgb <= "000000";
					when "11001101100101001" => rgb <= "000000";
					when "11001101100101010" => rgb <= "000000";
					when "11001101100101011" => rgb <= "000000";
					when "11001101100101100" => rgb <= "000000";
					when "11001101100101101" => rgb <= "000000";
					when "11001101100101110" => rgb <= "000000";
					when "11001101100101111" => rgb <= "000000";
					when "11001101100110000" => rgb <= "000000";
					when "11001101100110001" => rgb <= "000000";
					when "11001101100110010" => rgb <= "000000";
					when "11001101100110011" => rgb <= "000000";
					when "11001101100110100" => rgb <= "000000";
					when "11001101100110101" => rgb <= "000000";
					when "11001101100110110" => rgb <= "000000";
					when "11001101100110111" => rgb <= "000000";
					when "11001101100111000" => rgb <= "000000";
					when "11001101100111001" => rgb <= "000000";
					when "11001101100111010" => rgb <= "000000";
					when "11001101100111011" => rgb <= "000000";
					when "11001101100111100" => rgb <= "000000";
					when "11001101100111101" => rgb <= "000000";
					when "11001101100111110" => rgb <= "000000";
					when "11001101100111111" => rgb <= "000000";
					when "11001110000000000" => rgb <= "000000";
					when "11001110000000001" => rgb <= "000000";
					when "11001110000000010" => rgb <= "000000";
					when "11001110000000011" => rgb <= "000000";
					when "11001110000000100" => rgb <= "000000";
					when "11001110000000101" => rgb <= "000000";
					when "11001110000000110" => rgb <= "000000";
					when "11001110000000111" => rgb <= "000000";
					when "11001110000001000" => rgb <= "000000";
					when "11001110000001001" => rgb <= "000000";
					when "11001110000001010" => rgb <= "000000";
					when "11001110000001011" => rgb <= "000000";
					when "11001110000001100" => rgb <= "000000";
					when "11001110000001101" => rgb <= "000000";
					when "11001110000001110" => rgb <= "000000";
					when "11001110000001111" => rgb <= "000000";
					when "11001110000010000" => rgb <= "000000";
					when "11001110000010001" => rgb <= "000000";
					when "11001110000010010" => rgb <= "000000";
					when "11001110000010011" => rgb <= "000000";
					when "11001110000010100" => rgb <= "101010";
					when "11001110000010101" => rgb <= "111111";
					when "11001110000010110" => rgb <= "101010";
					when "11001110000010111" => rgb <= "111111";
					when "11001110000011000" => rgb <= "111111";
					when "11001110000011001" => rgb <= "111111";
					when "11001110000011010" => rgb <= "111111";
					when "11001110000011011" => rgb <= "111111";
					when "11001110000011100" => rgb <= "111111";
					when "11001110000011101" => rgb <= "111111";
					when "11001110000011110" => rgb <= "111111";
					when "11001110000011111" => rgb <= "111111";
					when "11001110000100000" => rgb <= "111111";
					when "11001110000100001" => rgb <= "101010";
					when "11001110000100010" => rgb <= "111111";
					when "11001110000100011" => rgb <= "000000";
					when "11001110000100100" => rgb <= "000000";
					when "11001110000100101" => rgb <= "000000";
					when "11001110000100110" => rgb <= "000000";
					when "11001110000100111" => rgb <= "000000";
					when "11001110000101000" => rgb <= "000000";
					when "11001110000101001" => rgb <= "000000";
					when "11001110000101010" => rgb <= "000000";
					when "11001110000101011" => rgb <= "000000";
					when "11001110000101100" => rgb <= "000000";
					when "11001110000101101" => rgb <= "000000";
					when "11001110000101110" => rgb <= "000000";
					when "11001110000101111" => rgb <= "000000";
					when "11001110000110000" => rgb <= "000000";
					when "11001110000110001" => rgb <= "000000";
					when "11001110000110010" => rgb <= "000000";
					when "11001110000110011" => rgb <= "000000";
					when "11001110000110100" => rgb <= "000000";
					when "11001110000110101" => rgb <= "000000";
					when "11001110000110110" => rgb <= "000000";
					when "11001110000110111" => rgb <= "000000";
					when "11001110000111000" => rgb <= "000000";
					when "11001110000111001" => rgb <= "000000";
					when "11001110000111010" => rgb <= "000000";
					when "11001110000111011" => rgb <= "000000";
					when "11001110000111100" => rgb <= "000000";
					when "11001110000111101" => rgb <= "000000";
					when "11001110000111110" => rgb <= "000000";
					when "11001110000111111" => rgb <= "000000";
					when "11001110001000000" => rgb <= "000000";
					when "11001110001000001" => rgb <= "101010";
					when "11001110001000010" => rgb <= "101010";
					when "11001110001000011" => rgb <= "101010";
					when "11001110001000100" => rgb <= "101010";
					when "11001110001000101" => rgb <= "101010";
					when "11001110001000110" => rgb <= "101010";
					when "11001110001000111" => rgb <= "101010";
					when "11001110001001000" => rgb <= "101010";
					when "11001110001001001" => rgb <= "101010";
					when "11001110001001010" => rgb <= "101010";
					when "11001110001001011" => rgb <= "101010";
					when "11001110001001100" => rgb <= "101010";
					when "11001110001001101" => rgb <= "101010";
					when "11001110001001110" => rgb <= "101010";
					when "11001110001001111" => rgb <= "101010";
					when "11001110001010000" => rgb <= "101010";
					when "11001110001010001" => rgb <= "111111";
					when "11001110001010010" => rgb <= "101010";
					when "11001110001010011" => rgb <= "101010";
					when "11001110001010100" => rgb <= "111111";
					when "11001110001010101" => rgb <= "101010";
					when "11001110001010110" => rgb <= "101010";
					when "11001110001010111" => rgb <= "101010";
					when "11001110001011000" => rgb <= "000000";
					when "11001110001011001" => rgb <= "000000";
					when "11001110001011010" => rgb <= "000000";
					when "11001110001011011" => rgb <= "000000";
					when "11001110001011100" => rgb <= "000000";
					when "11001110001011101" => rgb <= "000000";
					when "11001110001011110" => rgb <= "000000";
					when "11001110001011111" => rgb <= "000000";
					when "11001110001100000" => rgb <= "000000";
					when "11001110001100001" => rgb <= "000000";
					when "11001110001100010" => rgb <= "000000";
					when "11001110001100011" => rgb <= "000000";
					when "11001110001100100" => rgb <= "000000";
					when "11001110001100101" => rgb <= "000000";
					when "11001110001100110" => rgb <= "000000";
					when "11001110001100111" => rgb <= "000000";
					when "11001110001101000" => rgb <= "000000";
					when "11001110001101001" => rgb <= "000000";
					when "11001110001101010" => rgb <= "000000";
					when "11001110001101011" => rgb <= "000000";
					when "11001110001101100" => rgb <= "000000";
					when "11001110001101101" => rgb <= "000000";
					when "11001110001101110" => rgb <= "101010";
					when "11001110001101111" => rgb <= "101010";
					when "11001110001110000" => rgb <= "101010";
					when "11001110001110001" => rgb <= "101010";
					when "11001110001110010" => rgb <= "101010";
					when "11001110001110011" => rgb <= "101010";
					when "11001110001110100" => rgb <= "101010";
					when "11001110001110101" => rgb <= "101010";
					when "11001110001110110" => rgb <= "101010";
					when "11001110001110111" => rgb <= "101010";
					when "11001110001111000" => rgb <= "101010";
					when "11001110001111001" => rgb <= "101010";
					when "11001110001111010" => rgb <= "101010";
					when "11001110001111011" => rgb <= "101010";
					when "11001110001111100" => rgb <= "101010";
					when "11001110001111101" => rgb <= "111111";
					when "11001110001111110" => rgb <= "101010";
					when "11001110001111111" => rgb <= "101010";
					when "11001110010000000" => rgb <= "111111";
					when "11001110010000001" => rgb <= "101010";
					when "11001110010000010" => rgb <= "101010";
					when "11001110010000011" => rgb <= "111111";
					when "11001110010000100" => rgb <= "101010";
					when "11001110010000101" => rgb <= "000000";
					when "11001110010000110" => rgb <= "000000";
					when "11001110010000111" => rgb <= "000000";
					when "11001110010001000" => rgb <= "000000";
					when "11001110010001001" => rgb <= "000000";
					when "11001110010001010" => rgb <= "000000";
					when "11001110010001011" => rgb <= "000000";
					when "11001110010001100" => rgb <= "000000";
					when "11001110010001101" => rgb <= "000000";
					when "11001110010001110" => rgb <= "000000";
					when "11001110010001111" => rgb <= "000000";
					when "11001110010010000" => rgb <= "000000";
					when "11001110010010001" => rgb <= "000000";
					when "11001110010010010" => rgb <= "000000";
					when "11001110010010011" => rgb <= "000000";
					when "11001110010010100" => rgb <= "000000";
					when "11001110010010101" => rgb <= "000000";
					when "11001110010010110" => rgb <= "000000";
					when "11001110010010111" => rgb <= "000000";
					when "11001110010011000" => rgb <= "000000";
					when "11001110010011001" => rgb <= "000000";
					when "11001110010011010" => rgb <= "000000";
					when "11001110010011011" => rgb <= "000000";
					when "11001110010011100" => rgb <= "000000";
					when "11001110010011101" => rgb <= "000000";
					when "11001110010011110" => rgb <= "000000";
					when "11001110010011111" => rgb <= "000000";
					when "11001110010100000" => rgb <= "000000";
					when "11001110010100001" => rgb <= "000000";
					when "11001110010100010" => rgb <= "000000";
					when "11001110010100011" => rgb <= "000000";
					when "11001110010100100" => rgb <= "000000";
					when "11001110010100101" => rgb <= "000000";
					when "11001110010100110" => rgb <= "000000";
					when "11001110010100111" => rgb <= "000000";
					when "11001110010101000" => rgb <= "000000";
					when "11001110010101001" => rgb <= "000000";
					when "11001110010101010" => rgb <= "101010";
					when "11001110010101011" => rgb <= "101010";
					when "11001110010101100" => rgb <= "101010";
					when "11001110010101101" => rgb <= "101010";
					when "11001110010101110" => rgb <= "101010";
					when "11001110010101111" => rgb <= "101010";
					when "11001110010110000" => rgb <= "111111";
					when "11001110010110001" => rgb <= "010101";
					when "11001110010110010" => rgb <= "000000";
					when "11001110010110011" => rgb <= "000000";
					when "11001110010110100" => rgb <= "000000";
					when "11001110010110101" => rgb <= "000000";
					when "11001110010110110" => rgb <= "000000";
					when "11001110010110111" => rgb <= "000000";
					when "11001110010111000" => rgb <= "000000";
					when "11001110010111001" => rgb <= "101010";
					when "11001110010111010" => rgb <= "101010";
					when "11001110010111011" => rgb <= "101010";
					when "11001110010111100" => rgb <= "101010";
					when "11001110010111101" => rgb <= "101010";
					when "11001110010111110" => rgb <= "101010";
					when "11001110010111111" => rgb <= "101010";
					when "11001110011000000" => rgb <= "101010";
					when "11001110011000001" => rgb <= "111111";
					when "11001110011000010" => rgb <= "101010";
					when "11001110011000011" => rgb <= "101010";
					when "11001110011000100" => rgb <= "111111";
					when "11001110011000101" => rgb <= "111111";
					when "11001110011000110" => rgb <= "101010";
					when "11001110011000111" => rgb <= "111111";
					when "11001110011001000" => rgb <= "000000";
					when "11001110011001001" => rgb <= "000000";
					when "11001110011001010" => rgb <= "000000";
					when "11001110011001011" => rgb <= "000000";
					when "11001110011001100" => rgb <= "000000";
					when "11001110011001101" => rgb <= "000000";
					when "11001110011001110" => rgb <= "000000";
					when "11001110011001111" => rgb <= "000000";
					when "11001110011010000" => rgb <= "000000";
					when "11001110011010001" => rgb <= "000000";
					when "11001110011010010" => rgb <= "000000";
					when "11001110011010011" => rgb <= "000000";
					when "11001110011010100" => rgb <= "000000";
					when "11001110011010101" => rgb <= "000000";
					when "11001110011010110" => rgb <= "000000";
					when "11001110011010111" => rgb <= "101010";
					when "11001110011011000" => rgb <= "101010";
					when "11001110011011001" => rgb <= "101010";
					when "11001110011011010" => rgb <= "101010";
					when "11001110011011011" => rgb <= "111111";
					when "11001110011011100" => rgb <= "111111";
					when "11001110011011101" => rgb <= "111111";
					when "11001110011011110" => rgb <= "111111";
					when "11001110011011111" => rgb <= "111111";
					when "11001110011100000" => rgb <= "111111";
					when "11001110011100001" => rgb <= "111111";
					when "11001110011100010" => rgb <= "111111";
					when "11001110011100011" => rgb <= "101010";
					when "11001110011100100" => rgb <= "111111";
					when "11001110011100101" => rgb <= "111111";
					when "11001110011100110" => rgb <= "000000";
					when "11001110011100111" => rgb <= "000000";
					when "11001110011101000" => rgb <= "000000";
					when "11001110011101001" => rgb <= "000000";
					when "11001110011101010" => rgb <= "000000";
					when "11001110011101011" => rgb <= "000000";
					when "11001110011101100" => rgb <= "000000";
					when "11001110011101101" => rgb <= "010101";
					when "11001110011101110" => rgb <= "111111";
					when "11001110011101111" => rgb <= "101010";
					when "11001110011110000" => rgb <= "111111";
					when "11001110011110001" => rgb <= "111111";
					when "11001110011110010" => rgb <= "111111";
					when "11001110011110011" => rgb <= "101010";
					when "11001110011110100" => rgb <= "101010";
					when "11001110011110101" => rgb <= "000000";
					when "11001110011110110" => rgb <= "000000";
					when "11001110011110111" => rgb <= "000000";
					when "11001110011111000" => rgb <= "000000";
					when "11001110011111001" => rgb <= "000000";
					when "11001110011111010" => rgb <= "000000";
					when "11001110011111011" => rgb <= "000000";
					when "11001110011111100" => rgb <= "000000";
					when "11001110011111101" => rgb <= "000000";
					when "11001110011111110" => rgb <= "000000";
					when "11001110011111111" => rgb <= "000000";
					when "11001110100000000" => rgb <= "000000";
					when "11001110100000001" => rgb <= "000000";
					when "11001110100000010" => rgb <= "000000";
					when "11001110100000011" => rgb <= "000000";
					when "11001110100000100" => rgb <= "000000";
					when "11001110100000101" => rgb <= "000000";
					when "11001110100000110" => rgb <= "000000";
					when "11001110100000111" => rgb <= "000000";
					when "11001110100001000" => rgb <= "000000";
					when "11001110100001001" => rgb <= "000000";
					when "11001110100001010" => rgb <= "000000";
					when "11001110100001011" => rgb <= "010101";
					when "11001110100001100" => rgb <= "111111";
					when "11001110100001101" => rgb <= "101010";
					when "11001110100001110" => rgb <= "111111";
					when "11001110100001111" => rgb <= "111111";
					when "11001110100010000" => rgb <= "111111";
					when "11001110100010001" => rgb <= "111111";
					when "11001110100010010" => rgb <= "111111";
					when "11001110100010011" => rgb <= "111111";
					when "11001110100010100" => rgb <= "111111";
					when "11001110100010101" => rgb <= "111111";
					when "11001110100010110" => rgb <= "111111";
					when "11001110100010111" => rgb <= "111111";
					when "11001110100011000" => rgb <= "101010";
					when "11001110100011001" => rgb <= "101010";
					when "11001110100011010" => rgb <= "101010";
					when "11001110100011011" => rgb <= "000000";
					when "11001110100011100" => rgb <= "000000";
					when "11001110100011101" => rgb <= "000000";
					when "11001110100011110" => rgb <= "000000";
					when "11001110100011111" => rgb <= "000000";
					when "11001110100100000" => rgb <= "000000";
					when "11001110100100001" => rgb <= "000000";
					when "11001110100100010" => rgb <= "101010";
					when "11001110100100011" => rgb <= "101010";
					when "11001110100100100" => rgb <= "101010";
					when "11001110100100101" => rgb <= "101010";
					when "11001110100100110" => rgb <= "101010";
					when "11001110100100111" => rgb <= "101010";
					when "11001110100101000" => rgb <= "101010";
					when "11001110100101001" => rgb <= "101010";
					when "11001110100101010" => rgb <= "101010";
					when "11001110100101011" => rgb <= "101010";
					when "11001110100101100" => rgb <= "101010";
					when "11001110100101101" => rgb <= "101010";
					when "11001110100101110" => rgb <= "101010";
					when "11001110100101111" => rgb <= "101010";
					when "11001110100110000" => rgb <= "101010";
					when "11001110100110001" => rgb <= "000000";
					when "11001110100110010" => rgb <= "000000";
					when "11001110100110011" => rgb <= "000000";
					when "11001110100110100" => rgb <= "000000";
					when "11001110100110101" => rgb <= "000000";
					when "11001110100110110" => rgb <= "000000";
					when "11001110100110111" => rgb <= "000000";
					when "11001110100111000" => rgb <= "000000";
					when "11001110100111001" => rgb <= "000000";
					when "11001110100111010" => rgb <= "000000";
					when "11001110100111011" => rgb <= "000000";
					when "11001110100111100" => rgb <= "000000";
					when "11001110100111101" => rgb <= "000000";
					when "11001110100111110" => rgb <= "000000";
					when "11001110100111111" => rgb <= "000000";
					when "11001111000000000" => rgb <= "000000";
					when "11001111000000001" => rgb <= "000000";
					when "11001111000000010" => rgb <= "000000";
					when "11001111000000011" => rgb <= "000000";
					when "11001111000000100" => rgb <= "000000";
					when "11001111000000101" => rgb <= "000000";
					when "11001111000000110" => rgb <= "000000";
					when "11001111000000111" => rgb <= "000000";
					when "11001111000001000" => rgb <= "000000";
					when "11001111000001001" => rgb <= "000000";
					when "11001111000001010" => rgb <= "000000";
					when "11001111000001011" => rgb <= "000000";
					when "11001111000001100" => rgb <= "000000";
					when "11001111000001101" => rgb <= "000000";
					when "11001111000001110" => rgb <= "000000";
					when "11001111000001111" => rgb <= "000000";
					when "11001111000010000" => rgb <= "000000";
					when "11001111000010001" => rgb <= "000000";
					when "11001111000010010" => rgb <= "000000";
					when "11001111000010011" => rgb <= "000000";
					when "11001111000010100" => rgb <= "101010";
					when "11001111000010101" => rgb <= "111111";
					when "11001111000010110" => rgb <= "101010";
					when "11001111000010111" => rgb <= "111111";
					when "11001111000011000" => rgb <= "111111";
					when "11001111000011001" => rgb <= "111111";
					when "11001111000011010" => rgb <= "111111";
					when "11001111000011011" => rgb <= "111111";
					when "11001111000011100" => rgb <= "111111";
					when "11001111000011101" => rgb <= "111111";
					when "11001111000011110" => rgb <= "111111";
					when "11001111000011111" => rgb <= "111111";
					when "11001111000100000" => rgb <= "111111";
					when "11001111000100001" => rgb <= "101010";
					when "11001111000100010" => rgb <= "111111";
					when "11001111000100011" => rgb <= "000000";
					when "11001111000100100" => rgb <= "000000";
					when "11001111000100101" => rgb <= "000000";
					when "11001111000100110" => rgb <= "000000";
					when "11001111000100111" => rgb <= "000000";
					when "11001111000101000" => rgb <= "000000";
					when "11001111000101001" => rgb <= "000000";
					when "11001111000101010" => rgb <= "000000";
					when "11001111000101011" => rgb <= "000000";
					when "11001111000101100" => rgb <= "000000";
					when "11001111000101101" => rgb <= "000000";
					when "11001111000101110" => rgb <= "000000";
					when "11001111000101111" => rgb <= "000000";
					when "11001111000110000" => rgb <= "000000";
					when "11001111000110001" => rgb <= "000000";
					when "11001111000110010" => rgb <= "000000";
					when "11001111000110011" => rgb <= "000000";
					when "11001111000110100" => rgb <= "000000";
					when "11001111000110101" => rgb <= "000000";
					when "11001111000110110" => rgb <= "000000";
					when "11001111000110111" => rgb <= "000000";
					when "11001111000111000" => rgb <= "000000";
					when "11001111000111001" => rgb <= "000000";
					when "11001111000111010" => rgb <= "000000";
					when "11001111000111011" => rgb <= "000000";
					when "11001111000111100" => rgb <= "000000";
					when "11001111000111101" => rgb <= "000000";
					when "11001111000111110" => rgb <= "000000";
					when "11001111000111111" => rgb <= "000000";
					when "11001111001000000" => rgb <= "000000";
					when "11001111001000001" => rgb <= "101010";
					when "11001111001000010" => rgb <= "101010";
					when "11001111001000011" => rgb <= "111111";
					when "11001111001000100" => rgb <= "111111";
					when "11001111001000101" => rgb <= "111111";
					when "11001111001000110" => rgb <= "111111";
					when "11001111001000111" => rgb <= "101010";
					when "11001111001001000" => rgb <= "111111";
					when "11001111001001001" => rgb <= "111111";
					when "11001111001001010" => rgb <= "111111";
					when "11001111001001011" => rgb <= "111111";
					when "11001111001001100" => rgb <= "111111";
					when "11001111001001101" => rgb <= "111111";
					when "11001111001001110" => rgb <= "111111";
					when "11001111001001111" => rgb <= "111111";
					when "11001111001010000" => rgb <= "101010";
					when "11001111001010001" => rgb <= "101010";
					when "11001111001010010" => rgb <= "111111";
					when "11001111001010011" => rgb <= "111111";
					when "11001111001010100" => rgb <= "101010";
					when "11001111001010101" => rgb <= "101010";
					when "11001111001010110" => rgb <= "111111";
					when "11001111001010111" => rgb <= "010101";
					when "11001111001011000" => rgb <= "000000";
					when "11001111001011001" => rgb <= "000000";
					when "11001111001011010" => rgb <= "000000";
					when "11001111001011011" => rgb <= "000000";
					when "11001111001011100" => rgb <= "000000";
					when "11001111001011101" => rgb <= "000000";
					when "11001111001011110" => rgb <= "000000";
					when "11001111001011111" => rgb <= "000000";
					when "11001111001100000" => rgb <= "000000";
					when "11001111001100001" => rgb <= "000000";
					when "11001111001100010" => rgb <= "000000";
					when "11001111001100011" => rgb <= "000000";
					when "11001111001100100" => rgb <= "000000";
					when "11001111001100101" => rgb <= "000000";
					when "11001111001100110" => rgb <= "000000";
					when "11001111001100111" => rgb <= "000000";
					when "11001111001101000" => rgb <= "000000";
					when "11001111001101001" => rgb <= "000000";
					when "11001111001101010" => rgb <= "000000";
					when "11001111001101011" => rgb <= "000000";
					when "11001111001101100" => rgb <= "000000";
					when "11001111001101101" => rgb <= "000000";
					when "11001111001101110" => rgb <= "101010";
					when "11001111001101111" => rgb <= "111111";
					when "11001111001110000" => rgb <= "101010";
					when "11001111001110001" => rgb <= "111111";
					when "11001111001110010" => rgb <= "111111";
					when "11001111001110011" => rgb <= "111111";
					when "11001111001110100" => rgb <= "111111";
					when "11001111001110101" => rgb <= "111111";
					when "11001111001110110" => rgb <= "101010";
					when "11001111001110111" => rgb <= "111111";
					when "11001111001111000" => rgb <= "101010";
					when "11001111001111001" => rgb <= "111111";
					when "11001111001111010" => rgb <= "111111";
					when "11001111001111011" => rgb <= "101010";
					when "11001111001111100" => rgb <= "111111";
					when "11001111001111101" => rgb <= "111111";
					when "11001111001111110" => rgb <= "101010";
					when "11001111001111111" => rgb <= "111111";
					when "11001111010000000" => rgb <= "111111";
					when "11001111010000001" => rgb <= "111111";
					when "11001111010000010" => rgb <= "101010";
					when "11001111010000011" => rgb <= "111111";
					when "11001111010000100" => rgb <= "101010";
					when "11001111010000101" => rgb <= "000000";
					when "11001111010000110" => rgb <= "000000";
					when "11001111010000111" => rgb <= "000000";
					when "11001111010001000" => rgb <= "000000";
					when "11001111010001001" => rgb <= "000000";
					when "11001111010001010" => rgb <= "000000";
					when "11001111010001011" => rgb <= "000000";
					when "11001111010001100" => rgb <= "000000";
					when "11001111010001101" => rgb <= "000000";
					when "11001111010001110" => rgb <= "000000";
					when "11001111010001111" => rgb <= "000000";
					when "11001111010010000" => rgb <= "000000";
					when "11001111010010001" => rgb <= "000000";
					when "11001111010010010" => rgb <= "000000";
					when "11001111010010011" => rgb <= "000000";
					when "11001111010010100" => rgb <= "000000";
					when "11001111010010101" => rgb <= "000000";
					when "11001111010010110" => rgb <= "000000";
					when "11001111010010111" => rgb <= "000000";
					when "11001111010011000" => rgb <= "000000";
					when "11001111010011001" => rgb <= "000000";
					when "11001111010011010" => rgb <= "000000";
					when "11001111010011011" => rgb <= "000000";
					when "11001111010011100" => rgb <= "000000";
					when "11001111010011101" => rgb <= "000000";
					when "11001111010011110" => rgb <= "000000";
					when "11001111010011111" => rgb <= "000000";
					when "11001111010100000" => rgb <= "000000";
					when "11001111010100001" => rgb <= "000000";
					when "11001111010100010" => rgb <= "000000";
					when "11001111010100011" => rgb <= "000000";
					when "11001111010100100" => rgb <= "000000";
					when "11001111010100101" => rgb <= "000000";
					when "11001111010100110" => rgb <= "000000";
					when "11001111010100111" => rgb <= "000000";
					when "11001111010101000" => rgb <= "000000";
					when "11001111010101001" => rgb <= "000000";
					when "11001111010101010" => rgb <= "101010";
					when "11001111010101011" => rgb <= "111111";
					when "11001111010101100" => rgb <= "111111";
					when "11001111010101101" => rgb <= "101010";
					when "11001111010101110" => rgb <= "111111";
					when "11001111010101111" => rgb <= "101010";
					when "11001111010110000" => rgb <= "101010";
					when "11001111010110001" => rgb <= "010101";
					when "11001111010110010" => rgb <= "000000";
					when "11001111010110011" => rgb <= "000000";
					when "11001111010110100" => rgb <= "000000";
					when "11001111010110101" => rgb <= "000000";
					when "11001111010110110" => rgb <= "000000";
					when "11001111010110111" => rgb <= "000000";
					when "11001111010111000" => rgb <= "000000";
					when "11001111010111001" => rgb <= "101010";
					when "11001111010111010" => rgb <= "111111";
					when "11001111010111011" => rgb <= "111111";
					when "11001111010111100" => rgb <= "101010";
					when "11001111010111101" => rgb <= "111111";
					when "11001111010111110" => rgb <= "111111";
					when "11001111010111111" => rgb <= "111111";
					when "11001111011000000" => rgb <= "111111";
					when "11001111011000001" => rgb <= "101010";
					when "11001111011000010" => rgb <= "111111";
					when "11001111011000011" => rgb <= "111111";
					when "11001111011000100" => rgb <= "101010";
					when "11001111011000101" => rgb <= "111111";
					when "11001111011000110" => rgb <= "101010";
					when "11001111011000111" => rgb <= "101010";
					when "11001111011001000" => rgb <= "000000";
					when "11001111011001001" => rgb <= "000000";
					when "11001111011001010" => rgb <= "000000";
					when "11001111011001011" => rgb <= "000000";
					when "11001111011001100" => rgb <= "000000";
					when "11001111011001101" => rgb <= "000000";
					when "11001111011001110" => rgb <= "000000";
					when "11001111011001111" => rgb <= "000000";
					when "11001111011010000" => rgb <= "000000";
					when "11001111011010001" => rgb <= "000000";
					when "11001111011010010" => rgb <= "000000";
					when "11001111011010011" => rgb <= "000000";
					when "11001111011010100" => rgb <= "000000";
					when "11001111011010101" => rgb <= "000000";
					when "11001111011010110" => rgb <= "000000";
					when "11001111011010111" => rgb <= "101010";
					when "11001111011011000" => rgb <= "101010";
					when "11001111011011001" => rgb <= "101010";
					when "11001111011011010" => rgb <= "101010";
					when "11001111011011011" => rgb <= "111111";
					when "11001111011011100" => rgb <= "111111";
					when "11001111011011101" => rgb <= "111111";
					when "11001111011011110" => rgb <= "111111";
					when "11001111011011111" => rgb <= "111111";
					when "11001111011100000" => rgb <= "111111";
					when "11001111011100001" => rgb <= "111111";
					when "11001111011100010" => rgb <= "111111";
					when "11001111011100011" => rgb <= "101010";
					when "11001111011100100" => rgb <= "111111";
					when "11001111011100101" => rgb <= "111111";
					when "11001111011100110" => rgb <= "000000";
					when "11001111011100111" => rgb <= "000000";
					when "11001111011101000" => rgb <= "000000";
					when "11001111011101001" => rgb <= "000000";
					when "11001111011101010" => rgb <= "000000";
					when "11001111011101011" => rgb <= "000000";
					when "11001111011101100" => rgb <= "000000";
					when "11001111011101101" => rgb <= "010101";
					when "11001111011101110" => rgb <= "111111";
					when "11001111011101111" => rgb <= "101010";
					when "11001111011110000" => rgb <= "111111";
					when "11001111011110001" => rgb <= "111111";
					when "11001111011110010" => rgb <= "111111";
					when "11001111011110011" => rgb <= "101010";
					when "11001111011110100" => rgb <= "101010";
					when "11001111011110101" => rgb <= "000000";
					when "11001111011110110" => rgb <= "000000";
					when "11001111011110111" => rgb <= "000000";
					when "11001111011111000" => rgb <= "000000";
					when "11001111011111001" => rgb <= "000000";
					when "11001111011111010" => rgb <= "000000";
					when "11001111011111011" => rgb <= "000000";
					when "11001111011111100" => rgb <= "000000";
					when "11001111011111101" => rgb <= "000000";
					when "11001111011111110" => rgb <= "000000";
					when "11001111011111111" => rgb <= "000000";
					when "11001111100000000" => rgb <= "000000";
					when "11001111100000001" => rgb <= "000000";
					when "11001111100000010" => rgb <= "000000";
					when "11001111100000011" => rgb <= "000000";
					when "11001111100000100" => rgb <= "000000";
					when "11001111100000101" => rgb <= "000000";
					when "11001111100000110" => rgb <= "000000";
					when "11001111100000111" => rgb <= "000000";
					when "11001111100001000" => rgb <= "000000";
					when "11001111100001001" => rgb <= "000000";
					when "11001111100001010" => rgb <= "000000";
					when "11001111100001011" => rgb <= "010101";
					when "11001111100001100" => rgb <= "111111";
					when "11001111100001101" => rgb <= "101010";
					when "11001111100001110" => rgb <= "111111";
					when "11001111100001111" => rgb <= "111111";
					when "11001111100010000" => rgb <= "111111";
					when "11001111100010001" => rgb <= "111111";
					when "11001111100010010" => rgb <= "111111";
					when "11001111100010011" => rgb <= "111111";
					when "11001111100010100" => rgb <= "111111";
					when "11001111100010101" => rgb <= "111111";
					when "11001111100010110" => rgb <= "111111";
					when "11001111100010111" => rgb <= "111111";
					when "11001111100011000" => rgb <= "101010";
					when "11001111100011001" => rgb <= "101010";
					when "11001111100011010" => rgb <= "101010";
					when "11001111100011011" => rgb <= "000000";
					when "11001111100011100" => rgb <= "000000";
					when "11001111100011101" => rgb <= "000000";
					when "11001111100011110" => rgb <= "000000";
					when "11001111100011111" => rgb <= "000000";
					when "11001111100100000" => rgb <= "000000";
					when "11001111100100001" => rgb <= "000000";
					when "11001111100100010" => rgb <= "101010";
					when "11001111100100011" => rgb <= "101010";
					when "11001111100100100" => rgb <= "111111";
					when "11001111100100101" => rgb <= "111111";
					when "11001111100100110" => rgb <= "111111";
					when "11001111100100111" => rgb <= "111111";
					when "11001111100101000" => rgb <= "111111";
					when "11001111100101001" => rgb <= "111111";
					when "11001111100101010" => rgb <= "111111";
					when "11001111100101011" => rgb <= "101010";
					when "11001111100101100" => rgb <= "111111";
					when "11001111100101101" => rgb <= "111111";
					when "11001111100101110" => rgb <= "111111";
					when "11001111100101111" => rgb <= "111111";
					when "11001111100110000" => rgb <= "111111";
					when "11001111100110001" => rgb <= "000000";
					when "11001111100110010" => rgb <= "000000";
					when "11001111100110011" => rgb <= "000000";
					when "11001111100110100" => rgb <= "000000";
					when "11001111100110101" => rgb <= "000000";
					when "11001111100110110" => rgb <= "000000";
					when "11001111100110111" => rgb <= "000000";
					when "11001111100111000" => rgb <= "000000";
					when "11001111100111001" => rgb <= "000000";
					when "11001111100111010" => rgb <= "000000";
					when "11001111100111011" => rgb <= "000000";
					when "11001111100111100" => rgb <= "000000";
					when "11001111100111101" => rgb <= "000000";
					when "11001111100111110" => rgb <= "000000";
					when "11001111100111111" => rgb <= "000000";
					when "11010000000000000" => rgb <= "000000";
					when "11010000000000001" => rgb <= "000000";
					when "11010000000000010" => rgb <= "000000";
					when "11010000000000011" => rgb <= "000000";
					when "11010000000000100" => rgb <= "000000";
					when "11010000000000101" => rgb <= "000000";
					when "11010000000000110" => rgb <= "000000";
					when "11010000000000111" => rgb <= "000000";
					when "11010000000001000" => rgb <= "000000";
					when "11010000000001001" => rgb <= "000000";
					when "11010000000001010" => rgb <= "000000";
					when "11010000000001011" => rgb <= "000000";
					when "11010000000001100" => rgb <= "000000";
					when "11010000000001101" => rgb <= "000000";
					when "11010000000001110" => rgb <= "000000";
					when "11010000000001111" => rgb <= "000000";
					when "11010000000010000" => rgb <= "000000";
					when "11010000000010001" => rgb <= "000000";
					when "11010000000010010" => rgb <= "000000";
					when "11010000000010011" => rgb <= "000000";
					when "11010000000010100" => rgb <= "101010";
					when "11010000000010101" => rgb <= "111111";
					when "11010000000010110" => rgb <= "101010";
					when "11010000000010111" => rgb <= "101010";
					when "11010000000011000" => rgb <= "111111";
					when "11010000000011001" => rgb <= "111111";
					when "11010000000011010" => rgb <= "111111";
					when "11010000000011011" => rgb <= "101010";
					when "11010000000011100" => rgb <= "101010";
					when "11010000000011101" => rgb <= "111111";
					when "11010000000011110" => rgb <= "111111";
					when "11010000000011111" => rgb <= "101010";
					when "11010000000100000" => rgb <= "101010";
					when "11010000000100001" => rgb <= "111111";
					when "11010000000100010" => rgb <= "101010";
					when "11010000000100011" => rgb <= "000000";
					when "11010000000100100" => rgb <= "000000";
					when "11010000000100101" => rgb <= "000000";
					when "11010000000100110" => rgb <= "000000";
					when "11010000000100111" => rgb <= "000000";
					when "11010000000101000" => rgb <= "000000";
					when "11010000000101001" => rgb <= "000000";
					when "11010000000101010" => rgb <= "000000";
					when "11010000000101011" => rgb <= "000000";
					when "11010000000101100" => rgb <= "000000";
					when "11010000000101101" => rgb <= "000000";
					when "11010000000101110" => rgb <= "000000";
					when "11010000000101111" => rgb <= "000000";
					when "11010000000110000" => rgb <= "000000";
					when "11010000000110001" => rgb <= "000000";
					when "11010000000110010" => rgb <= "000000";
					when "11010000000110011" => rgb <= "000000";
					when "11010000000110100" => rgb <= "000000";
					when "11010000000110101" => rgb <= "000000";
					when "11010000000110110" => rgb <= "000000";
					when "11010000000110111" => rgb <= "000000";
					when "11010000000111000" => rgb <= "000000";
					when "11010000000111001" => rgb <= "000000";
					when "11010000000111010" => rgb <= "000000";
					when "11010000000111011" => rgb <= "000000";
					when "11010000000111100" => rgb <= "000000";
					when "11010000000111101" => rgb <= "000000";
					when "11010000000111110" => rgb <= "000000";
					when "11010000000111111" => rgb <= "000000";
					when "11010000001000000" => rgb <= "000000";
					when "11010000001000001" => rgb <= "101010";
					when "11010000001000010" => rgb <= "111111";
					when "11010000001000011" => rgb <= "111111";
					when "11010000001000100" => rgb <= "101010";
					when "11010000001000101" => rgb <= "101010";
					when "11010000001000110" => rgb <= "111111";
					when "11010000001000111" => rgb <= "101010";
					when "11010000001001000" => rgb <= "101010";
					when "11010000001001001" => rgb <= "101010";
					when "11010000001001010" => rgb <= "111111";
					when "11010000001001011" => rgb <= "111111";
					when "11010000001001100" => rgb <= "101010";
					when "11010000001001101" => rgb <= "101010";
					when "11010000001001110" => rgb <= "101010";
					when "11010000001001111" => rgb <= "111111";
					when "11010000001010000" => rgb <= "111111";
					when "11010000001010001" => rgb <= "101010";
					when "11010000001010010" => rgb <= "101010";
					when "11010000001010011" => rgb <= "101010";
					when "11010000001010100" => rgb <= "101010";
					when "11010000001010101" => rgb <= "101010";
					when "11010000001010110" => rgb <= "111111";
					when "11010000001010111" => rgb <= "101010";
					when "11010000001011000" => rgb <= "000000";
					when "11010000001011001" => rgb <= "000000";
					when "11010000001011010" => rgb <= "000000";
					when "11010000001011011" => rgb <= "000000";
					when "11010000001011100" => rgb <= "000000";
					when "11010000001011101" => rgb <= "000000";
					when "11010000001011110" => rgb <= "000000";
					when "11010000001011111" => rgb <= "000000";
					when "11010000001100000" => rgb <= "000000";
					when "11010000001100001" => rgb <= "000000";
					when "11010000001100010" => rgb <= "000000";
					when "11010000001100011" => rgb <= "000000";
					when "11010000001100100" => rgb <= "000000";
					when "11010000001100101" => rgb <= "000000";
					when "11010000001100110" => rgb <= "000000";
					when "11010000001100111" => rgb <= "000000";
					when "11010000001101000" => rgb <= "000000";
					when "11010000001101001" => rgb <= "000000";
					when "11010000001101010" => rgb <= "000000";
					when "11010000001101011" => rgb <= "000000";
					when "11010000001101100" => rgb <= "000000";
					when "11010000001101101" => rgb <= "000000";
					when "11010000001101110" => rgb <= "101010";
					when "11010000001101111" => rgb <= "111111";
					when "11010000001110000" => rgb <= "101010";
					when "11010000001110001" => rgb <= "101010";
					when "11010000001110010" => rgb <= "111111";
					when "11010000001110011" => rgb <= "111111";
					when "11010000001110100" => rgb <= "101010";
					when "11010000001110101" => rgb <= "111111";
					when "11010000001110110" => rgb <= "111111";
					when "11010000001110111" => rgb <= "101010";
					when "11010000001111000" => rgb <= "101010";
					when "11010000001111001" => rgb <= "101010";
					when "11010000001111010" => rgb <= "101010";
					when "11010000001111011" => rgb <= "101010";
					when "11010000001111100" => rgb <= "101010";
					when "11010000001111101" => rgb <= "101010";
					when "11010000001111110" => rgb <= "101010";
					when "11010000001111111" => rgb <= "101010";
					when "11010000010000000" => rgb <= "111111";
					when "11010000010000001" => rgb <= "101010";
					when "11010000010000010" => rgb <= "111111";
					when "11010000010000011" => rgb <= "101010";
					when "11010000010000100" => rgb <= "101010";
					when "11010000010000101" => rgb <= "000000";
					when "11010000010000110" => rgb <= "000000";
					when "11010000010000111" => rgb <= "000000";
					when "11010000010001000" => rgb <= "000000";
					when "11010000010001001" => rgb <= "000000";
					when "11010000010001010" => rgb <= "000000";
					when "11010000010001011" => rgb <= "000000";
					when "11010000010001100" => rgb <= "000000";
					when "11010000010001101" => rgb <= "000000";
					when "11010000010001110" => rgb <= "000000";
					when "11010000010001111" => rgb <= "000000";
					when "11010000010010000" => rgb <= "000000";
					when "11010000010010001" => rgb <= "000000";
					when "11010000010010010" => rgb <= "000000";
					when "11010000010010011" => rgb <= "000000";
					when "11010000010010100" => rgb <= "000000";
					when "11010000010010101" => rgb <= "000000";
					when "11010000010010110" => rgb <= "000000";
					when "11010000010010111" => rgb <= "000000";
					when "11010000010011000" => rgb <= "000000";
					when "11010000010011001" => rgb <= "000000";
					when "11010000010011010" => rgb <= "000000";
					when "11010000010011011" => rgb <= "000000";
					when "11010000010011100" => rgb <= "000000";
					when "11010000010011101" => rgb <= "000000";
					when "11010000010011110" => rgb <= "000000";
					when "11010000010011111" => rgb <= "000000";
					when "11010000010100000" => rgb <= "000000";
					when "11010000010100001" => rgb <= "000000";
					when "11010000010100010" => rgb <= "000000";
					when "11010000010100011" => rgb <= "000000";
					when "11010000010100100" => rgb <= "000000";
					when "11010000010100101" => rgb <= "000000";
					when "11010000010100110" => rgb <= "000000";
					when "11010000010100111" => rgb <= "000000";
					when "11010000010101000" => rgb <= "000000";
					when "11010000010101001" => rgb <= "000000";
					when "11010000010101010" => rgb <= "101010";
					when "11010000010101011" => rgb <= "101010";
					when "11010000010101100" => rgb <= "101010";
					when "11010000010101101" => rgb <= "111111";
					when "11010000010101110" => rgb <= "111111";
					when "11010000010101111" => rgb <= "101010";
					when "11010000010110000" => rgb <= "101010";
					when "11010000010110001" => rgb <= "010101";
					when "11010000010110010" => rgb <= "000000";
					when "11010000010110011" => rgb <= "000000";
					when "11010000010110100" => rgb <= "000000";
					when "11010000010110101" => rgb <= "000000";
					when "11010000010110110" => rgb <= "000000";
					when "11010000010110111" => rgb <= "000000";
					when "11010000010111000" => rgb <= "000000";
					when "11010000010111001" => rgb <= "101010";
					when "11010000010111010" => rgb <= "111111";
					when "11010000010111011" => rgb <= "101010";
					when "11010000010111100" => rgb <= "101010";
					when "11010000010111101" => rgb <= "101010";
					when "11010000010111110" => rgb <= "111111";
					when "11010000010111111" => rgb <= "101010";
					when "11010000011000000" => rgb <= "101010";
					when "11010000011000001" => rgb <= "111111";
					when "11010000011000010" => rgb <= "111111";
					when "11010000011000011" => rgb <= "101010";
					when "11010000011000100" => rgb <= "111111";
					when "11010000011000101" => rgb <= "111111";
					when "11010000011000110" => rgb <= "101010";
					when "11010000011000111" => rgb <= "101010";
					when "11010000011001000" => rgb <= "000000";
					when "11010000011001001" => rgb <= "000000";
					when "11010000011001010" => rgb <= "000000";
					when "11010000011001011" => rgb <= "000000";
					when "11010000011001100" => rgb <= "000000";
					when "11010000011001101" => rgb <= "000000";
					when "11010000011001110" => rgb <= "000000";
					when "11010000011001111" => rgb <= "000000";
					when "11010000011010000" => rgb <= "000000";
					when "11010000011010001" => rgb <= "000000";
					when "11010000011010010" => rgb <= "000000";
					when "11010000011010011" => rgb <= "000000";
					when "11010000011010100" => rgb <= "000000";
					when "11010000011010101" => rgb <= "000000";
					when "11010000011010110" => rgb <= "000000";
					when "11010000011010111" => rgb <= "101010";
					when "11010000011011000" => rgb <= "111111";
					when "11010000011011001" => rgb <= "111111";
					when "11010000011011010" => rgb <= "101010";
					when "11010000011011011" => rgb <= "101010";
					when "11010000011011100" => rgb <= "111111";
					when "11010000011011101" => rgb <= "111111";
					when "11010000011011110" => rgb <= "111111";
					when "11010000011011111" => rgb <= "111111";
					when "11010000011100000" => rgb <= "111111";
					when "11010000011100001" => rgb <= "111111";
					when "11010000011100010" => rgb <= "101010";
					when "11010000011100011" => rgb <= "111111";
					when "11010000011100100" => rgb <= "111111";
					when "11010000011100101" => rgb <= "111111";
					when "11010000011100110" => rgb <= "000000";
					when "11010000011100111" => rgb <= "000000";
					when "11010000011101000" => rgb <= "000000";
					when "11010000011101001" => rgb <= "000000";
					when "11010000011101010" => rgb <= "000000";
					when "11010000011101011" => rgb <= "000000";
					when "11010000011101100" => rgb <= "000000";
					when "11010000011101101" => rgb <= "010101";
					when "11010000011101110" => rgb <= "101010";
					when "11010000011101111" => rgb <= "111111";
					when "11010000011110000" => rgb <= "111111";
					when "11010000011110001" => rgb <= "101010";
					when "11010000011110010" => rgb <= "101010";
					when "11010000011110011" => rgb <= "111111";
					when "11010000011110100" => rgb <= "101010";
					when "11010000011110101" => rgb <= "000000";
					when "11010000011110110" => rgb <= "000000";
					when "11010000011110111" => rgb <= "000000";
					when "11010000011111000" => rgb <= "000000";
					when "11010000011111001" => rgb <= "000000";
					when "11010000011111010" => rgb <= "000000";
					when "11010000011111011" => rgb <= "000000";
					when "11010000011111100" => rgb <= "000000";
					when "11010000011111101" => rgb <= "000000";
					when "11010000011111110" => rgb <= "000000";
					when "11010000011111111" => rgb <= "000000";
					when "11010000100000000" => rgb <= "000000";
					when "11010000100000001" => rgb <= "000000";
					when "11010000100000010" => rgb <= "000000";
					when "11010000100000011" => rgb <= "000000";
					when "11010000100000100" => rgb <= "000000";
					when "11010000100000101" => rgb <= "000000";
					when "11010000100000110" => rgb <= "000000";
					when "11010000100000111" => rgb <= "000000";
					when "11010000100001000" => rgb <= "000000";
					when "11010000100001001" => rgb <= "000000";
					when "11010000100001010" => rgb <= "000000";
					when "11010000100001011" => rgb <= "010101";
					when "11010000100001100" => rgb <= "101010";
					when "11010000100001101" => rgb <= "101010";
					when "11010000100001110" => rgb <= "111111";
					when "11010000100001111" => rgb <= "101010";
					when "11010000100010000" => rgb <= "111111";
					when "11010000100010001" => rgb <= "111111";
					when "11010000100010010" => rgb <= "111111";
					when "11010000100010011" => rgb <= "111111";
					when "11010000100010100" => rgb <= "111111";
					when "11010000100010101" => rgb <= "111111";
					when "11010000100010110" => rgb <= "111111";
					when "11010000100010111" => rgb <= "111111";
					when "11010000100011000" => rgb <= "111111";
					when "11010000100011001" => rgb <= "101010";
					when "11010000100011010" => rgb <= "101010";
					when "11010000100011011" => rgb <= "000000";
					when "11010000100011100" => rgb <= "000000";
					when "11010000100011101" => rgb <= "000000";
					when "11010000100011110" => rgb <= "000000";
					when "11010000100011111" => rgb <= "000000";
					when "11010000100100000" => rgb <= "000000";
					when "11010000100100001" => rgb <= "000000";
					when "11010000100100010" => rgb <= "101010";
					when "11010000100100011" => rgb <= "101010";
					when "11010000100100100" => rgb <= "111111";
					when "11010000100100101" => rgb <= "101010";
					when "11010000100100110" => rgb <= "101010";
					when "11010000100100111" => rgb <= "111111";
					when "11010000100101000" => rgb <= "101010";
					when "11010000100101001" => rgb <= "101010";
					when "11010000100101010" => rgb <= "101010";
					when "11010000100101011" => rgb <= "101010";
					when "11010000100101100" => rgb <= "111111";
					when "11010000100101101" => rgb <= "111111";
					when "11010000100101110" => rgb <= "101010";
					when "11010000100101111" => rgb <= "101010";
					when "11010000100110000" => rgb <= "101010";
					when "11010000100110001" => rgb <= "000000";
					when "11010000100110010" => rgb <= "000000";
					when "11010000100110011" => rgb <= "000000";
					when "11010000100110100" => rgb <= "000000";
					when "11010000100110101" => rgb <= "000000";
					when "11010000100110110" => rgb <= "000000";
					when "11010000100110111" => rgb <= "000000";
					when "11010000100111000" => rgb <= "000000";
					when "11010000100111001" => rgb <= "000000";
					when "11010000100111010" => rgb <= "000000";
					when "11010000100111011" => rgb <= "000000";
					when "11010000100111100" => rgb <= "000000";
					when "11010000100111101" => rgb <= "000000";
					when "11010000100111110" => rgb <= "000000";
					when "11010000100111111" => rgb <= "000000";
					when "11010001000000000" => rgb <= "000000";
					when "11010001000000001" => rgb <= "000000";
					when "11010001000000010" => rgb <= "000000";
					when "11010001000000011" => rgb <= "000000";
					when "11010001000000100" => rgb <= "000000";
					when "11010001000000101" => rgb <= "000000";
					when "11010001000000110" => rgb <= "000000";
					when "11010001000000111" => rgb <= "000000";
					when "11010001000001000" => rgb <= "000000";
					when "11010001000001001" => rgb <= "000000";
					when "11010001000001010" => rgb <= "000000";
					when "11010001000001011" => rgb <= "000000";
					when "11010001000001100" => rgb <= "000000";
					when "11010001000001101" => rgb <= "000000";
					when "11010001000001110" => rgb <= "000000";
					when "11010001000001111" => rgb <= "000000";
					when "11010001000010000" => rgb <= "000000";
					when "11010001000010001" => rgb <= "000000";
					when "11010001000010010" => rgb <= "000000";
					when "11010001000010011" => rgb <= "000000";
					when "11010001000010100" => rgb <= "101010";
					when "11010001000010101" => rgb <= "111111";
					when "11010001000010110" => rgb <= "101010";
					when "11010001000010111" => rgb <= "111111";
					when "11010001000011000" => rgb <= "101010";
					when "11010001000011001" => rgb <= "101010";
					when "11010001000011010" => rgb <= "111111";
					when "11010001000011011" => rgb <= "101010";
					when "11010001000011100" => rgb <= "101010";
					when "11010001000011101" => rgb <= "111111";
					when "11010001000011110" => rgb <= "111111";
					when "11010001000011111" => rgb <= "111111";
					when "11010001000100000" => rgb <= "101010";
					when "11010001000100001" => rgb <= "111111";
					when "11010001000100010" => rgb <= "111111";
					when "11010001000100011" => rgb <= "000000";
					when "11010001000100100" => rgb <= "000000";
					when "11010001000100101" => rgb <= "000000";
					when "11010001000100110" => rgb <= "000000";
					when "11010001000100111" => rgb <= "000000";
					when "11010001000101000" => rgb <= "000000";
					when "11010001000101001" => rgb <= "000000";
					when "11010001000101010" => rgb <= "000000";
					when "11010001000101011" => rgb <= "000000";
					when "11010001000101100" => rgb <= "000000";
					when "11010001000101101" => rgb <= "000000";
					when "11010001000101110" => rgb <= "000000";
					when "11010001000101111" => rgb <= "000000";
					when "11010001000110000" => rgb <= "000000";
					when "11010001000110001" => rgb <= "000000";
					when "11010001000110010" => rgb <= "000000";
					when "11010001000110011" => rgb <= "000000";
					when "11010001000110100" => rgb <= "000000";
					when "11010001000110101" => rgb <= "000000";
					when "11010001000110110" => rgb <= "000000";
					when "11010001000110111" => rgb <= "000000";
					when "11010001000111000" => rgb <= "000000";
					when "11010001000111001" => rgb <= "000000";
					when "11010001000111010" => rgb <= "000000";
					when "11010001000111011" => rgb <= "000000";
					when "11010001000111100" => rgb <= "000000";
					when "11010001000111101" => rgb <= "000000";
					when "11010001000111110" => rgb <= "000000";
					when "11010001000111111" => rgb <= "000000";
					when "11010001001000000" => rgb <= "000000";
					when "11010001001000001" => rgb <= "101010";
					when "11010001001000010" => rgb <= "111111";
					when "11010001001000011" => rgb <= "101010";
					when "11010001001000100" => rgb <= "111111";
					when "11010001001000101" => rgb <= "111111";
					when "11010001001000110" => rgb <= "101010";
					when "11010001001000111" => rgb <= "111111";
					when "11010001001001000" => rgb <= "101010";
					when "11010001001001001" => rgb <= "101010";
					when "11010001001001010" => rgb <= "101010";
					when "11010001001001011" => rgb <= "101010";
					when "11010001001001100" => rgb <= "101010";
					when "11010001001001101" => rgb <= "101010";
					when "11010001001001110" => rgb <= "101010";
					when "11010001001001111" => rgb <= "101010";
					when "11010001001010000" => rgb <= "111111";
					when "11010001001010001" => rgb <= "101010";
					when "11010001001010010" => rgb <= "101010";
					when "11010001001010011" => rgb <= "111111";
					when "11010001001010100" => rgb <= "111111";
					when "11010001001010101" => rgb <= "101010";
					when "11010001001010110" => rgb <= "111111";
					when "11010001001010111" => rgb <= "010101";
					when "11010001001011000" => rgb <= "000000";
					when "11010001001011001" => rgb <= "000000";
					when "11010001001011010" => rgb <= "000000";
					when "11010001001011011" => rgb <= "000000";
					when "11010001001011100" => rgb <= "000000";
					when "11010001001011101" => rgb <= "000000";
					when "11010001001011110" => rgb <= "000000";
					when "11010001001011111" => rgb <= "000000";
					when "11010001001100000" => rgb <= "000000";
					when "11010001001100001" => rgb <= "000000";
					when "11010001001100010" => rgb <= "000000";
					when "11010001001100011" => rgb <= "000000";
					when "11010001001100100" => rgb <= "000000";
					when "11010001001100101" => rgb <= "000000";
					when "11010001001100110" => rgb <= "000000";
					when "11010001001100111" => rgb <= "000000";
					when "11010001001101000" => rgb <= "000000";
					when "11010001001101001" => rgb <= "000000";
					when "11010001001101010" => rgb <= "000000";
					when "11010001001101011" => rgb <= "000000";
					when "11010001001101100" => rgb <= "000000";
					when "11010001001101101" => rgb <= "000000";
					when "11010001001101110" => rgb <= "101010";
					when "11010001001101111" => rgb <= "111111";
					when "11010001001110000" => rgb <= "101010";
					when "11010001001110001" => rgb <= "111111";
					when "11010001001110010" => rgb <= "111111";
					when "11010001001110011" => rgb <= "111111";
					when "11010001001110100" => rgb <= "111111";
					when "11010001001110101" => rgb <= "111111";
					when "11010001001110110" => rgb <= "111111";
					when "11010001001110111" => rgb <= "101010";
					when "11010001001111000" => rgb <= "101010";
					when "11010001001111001" => rgb <= "101010";
					when "11010001001111010" => rgb <= "101010";
					when "11010001001111011" => rgb <= "101010";
					when "11010001001111100" => rgb <= "101010";
					when "11010001001111101" => rgb <= "101010";
					when "11010001001111110" => rgb <= "101010";
					when "11010001001111111" => rgb <= "101010";
					when "11010001010000000" => rgb <= "111111";
					when "11010001010000001" => rgb <= "101010";
					when "11010001010000010" => rgb <= "111111";
					when "11010001010000011" => rgb <= "111111";
					when "11010001010000100" => rgb <= "101010";
					when "11010001010000101" => rgb <= "000000";
					when "11010001010000110" => rgb <= "000000";
					when "11010001010000111" => rgb <= "000000";
					when "11010001010001000" => rgb <= "000000";
					when "11010001010001001" => rgb <= "000000";
					when "11010001010001010" => rgb <= "000000";
					when "11010001010001011" => rgb <= "000000";
					when "11010001010001100" => rgb <= "000000";
					when "11010001010001101" => rgb <= "000000";
					when "11010001010001110" => rgb <= "000000";
					when "11010001010001111" => rgb <= "000000";
					when "11010001010010000" => rgb <= "000000";
					when "11010001010010001" => rgb <= "000000";
					when "11010001010010010" => rgb <= "000000";
					when "11010001010010011" => rgb <= "000000";
					when "11010001010010100" => rgb <= "000000";
					when "11010001010010101" => rgb <= "000000";
					when "11010001010010110" => rgb <= "000000";
					when "11010001010010111" => rgb <= "000000";
					when "11010001010011000" => rgb <= "000000";
					when "11010001010011001" => rgb <= "000000";
					when "11010001010011010" => rgb <= "000000";
					when "11010001010011011" => rgb <= "000000";
					when "11010001010011100" => rgb <= "000000";
					when "11010001010011101" => rgb <= "000000";
					when "11010001010011110" => rgb <= "000000";
					when "11010001010011111" => rgb <= "000000";
					when "11010001010100000" => rgb <= "000000";
					when "11010001010100001" => rgb <= "000000";
					when "11010001010100010" => rgb <= "000000";
					when "11010001010100011" => rgb <= "000000";
					when "11010001010100100" => rgb <= "000000";
					when "11010001010100101" => rgb <= "000000";
					when "11010001010100110" => rgb <= "000000";
					when "11010001010100111" => rgb <= "000000";
					when "11010001010101000" => rgb <= "000000";
					when "11010001010101001" => rgb <= "000000";
					when "11010001010101010" => rgb <= "101010";
					when "11010001010101011" => rgb <= "111111";
					when "11010001010101100" => rgb <= "101010";
					when "11010001010101101" => rgb <= "111111";
					when "11010001010101110" => rgb <= "101010";
					when "11010001010101111" => rgb <= "101010";
					when "11010001010110000" => rgb <= "111111";
					when "11010001010110001" => rgb <= "101010";
					when "11010001010110010" => rgb <= "000000";
					when "11010001010110011" => rgb <= "000000";
					when "11010001010110100" => rgb <= "000000";
					when "11010001010110101" => rgb <= "000000";
					when "11010001010110110" => rgb <= "000000";
					when "11010001010110111" => rgb <= "000000";
					when "11010001010111000" => rgb <= "000000";
					when "11010001010111001" => rgb <= "101010";
					when "11010001010111010" => rgb <= "101010";
					when "11010001010111011" => rgb <= "101010";
					when "11010001010111100" => rgb <= "111111";
					when "11010001010111101" => rgb <= "111111";
					when "11010001010111110" => rgb <= "101010";
					when "11010001010111111" => rgb <= "111111";
					when "11010001011000000" => rgb <= "101010";
					when "11010001011000001" => rgb <= "111111";
					when "11010001011000010" => rgb <= "101010";
					when "11010001011000011" => rgb <= "101010";
					when "11010001011000100" => rgb <= "111111";
					when "11010001011000101" => rgb <= "111111";
					when "11010001011000110" => rgb <= "101010";
					when "11010001011000111" => rgb <= "111111";
					when "11010001011001000" => rgb <= "000000";
					when "11010001011001001" => rgb <= "000000";
					when "11010001011001010" => rgb <= "000000";
					when "11010001011001011" => rgb <= "000000";
					when "11010001011001100" => rgb <= "000000";
					when "11010001011001101" => rgb <= "000000";
					when "11010001011001110" => rgb <= "000000";
					when "11010001011001111" => rgb <= "000000";
					when "11010001011010000" => rgb <= "000000";
					when "11010001011010001" => rgb <= "000000";
					when "11010001011010010" => rgb <= "000000";
					when "11010001011010011" => rgb <= "000000";
					when "11010001011010100" => rgb <= "000000";
					when "11010001011010101" => rgb <= "000000";
					when "11010001011010110" => rgb <= "000000";
					when "11010001011010111" => rgb <= "101010";
					when "11010001011011000" => rgb <= "101010";
					when "11010001011011001" => rgb <= "101010";
					when "11010001011011010" => rgb <= "101010";
					when "11010001011011011" => rgb <= "101010";
					when "11010001011011100" => rgb <= "111111";
					when "11010001011011101" => rgb <= "111111";
					when "11010001011011110" => rgb <= "111111";
					when "11010001011011111" => rgb <= "111111";
					when "11010001011100000" => rgb <= "111111";
					when "11010001011100001" => rgb <= "111111";
					when "11010001011100010" => rgb <= "111111";
					when "11010001011100011" => rgb <= "111111";
					when "11010001011100100" => rgb <= "101010";
					when "11010001011100101" => rgb <= "111111";
					when "11010001011100110" => rgb <= "000000";
					when "11010001011100111" => rgb <= "000000";
					when "11010001011101000" => rgb <= "000000";
					when "11010001011101001" => rgb <= "000000";
					when "11010001011101010" => rgb <= "000000";
					when "11010001011101011" => rgb <= "000000";
					when "11010001011101100" => rgb <= "000000";
					when "11010001011101101" => rgb <= "010101";
					when "11010001011101110" => rgb <= "101010";
					when "11010001011101111" => rgb <= "101010";
					when "11010001011110000" => rgb <= "101010";
					when "11010001011110001" => rgb <= "101010";
					when "11010001011110010" => rgb <= "101010";
					when "11010001011110011" => rgb <= "101010";
					when "11010001011110100" => rgb <= "101010";
					when "11010001011110101" => rgb <= "000000";
					when "11010001011110110" => rgb <= "000000";
					when "11010001011110111" => rgb <= "000000";
					when "11010001011111000" => rgb <= "000000";
					when "11010001011111001" => rgb <= "000000";
					when "11010001011111010" => rgb <= "000000";
					when "11010001011111011" => rgb <= "000000";
					when "11010001011111100" => rgb <= "000000";
					when "11010001011111101" => rgb <= "000000";
					when "11010001011111110" => rgb <= "000000";
					when "11010001011111111" => rgb <= "000000";
					when "11010001100000000" => rgb <= "000000";
					when "11010001100000001" => rgb <= "000000";
					when "11010001100000010" => rgb <= "000000";
					when "11010001100000011" => rgb <= "000000";
					when "11010001100000100" => rgb <= "000000";
					when "11010001100000101" => rgb <= "000000";
					when "11010001100000110" => rgb <= "000000";
					when "11010001100000111" => rgb <= "000000";
					when "11010001100001000" => rgb <= "000000";
					when "11010001100001001" => rgb <= "000000";
					when "11010001100001010" => rgb <= "000000";
					when "11010001100001011" => rgb <= "010101";
					when "11010001100001100" => rgb <= "111111";
					when "11010001100001101" => rgb <= "101010";
					when "11010001100001110" => rgb <= "101010";
					when "11010001100001111" => rgb <= "101010";
					when "11010001100010000" => rgb <= "111111";
					when "11010001100010001" => rgb <= "111111";
					when "11010001100010010" => rgb <= "111111";
					when "11010001100010011" => rgb <= "111111";
					when "11010001100010100" => rgb <= "111111";
					when "11010001100010101" => rgb <= "111111";
					when "11010001100010110" => rgb <= "111111";
					when "11010001100010111" => rgb <= "111111";
					when "11010001100011000" => rgb <= "101010";
					when "11010001100011001" => rgb <= "101010";
					when "11010001100011010" => rgb <= "101010";
					when "11010001100011011" => rgb <= "000000";
					when "11010001100011100" => rgb <= "000000";
					when "11010001100011101" => rgb <= "000000";
					when "11010001100011110" => rgb <= "000000";
					when "11010001100011111" => rgb <= "000000";
					when "11010001100100000" => rgb <= "000000";
					when "11010001100100001" => rgb <= "000000";
					when "11010001100100010" => rgb <= "101010";
					when "11010001100100011" => rgb <= "111111";
					when "11010001100100100" => rgb <= "111111";
					when "11010001100100101" => rgb <= "111111";
					when "11010001100100110" => rgb <= "101010";
					when "11010001100100111" => rgb <= "101010";
					when "11010001100101000" => rgb <= "111111";
					when "11010001100101001" => rgb <= "111111";
					when "11010001100101010" => rgb <= "111111";
					when "11010001100101011" => rgb <= "111111";
					when "11010001100101100" => rgb <= "111111";
					when "11010001100101101" => rgb <= "111111";
					when "11010001100101110" => rgb <= "111111";
					when "11010001100101111" => rgb <= "101010";
					when "11010001100110000" => rgb <= "101010";
					when "11010001100110001" => rgb <= "000000";
					when "11010001100110010" => rgb <= "000000";
					when "11010001100110011" => rgb <= "000000";
					when "11010001100110100" => rgb <= "000000";
					when "11010001100110101" => rgb <= "000000";
					when "11010001100110110" => rgb <= "000000";
					when "11010001100110111" => rgb <= "000000";
					when "11010001100111000" => rgb <= "000000";
					when "11010001100111001" => rgb <= "000000";
					when "11010001100111010" => rgb <= "000000";
					when "11010001100111011" => rgb <= "000000";
					when "11010001100111100" => rgb <= "000000";
					when "11010001100111101" => rgb <= "000000";
					when "11010001100111110" => rgb <= "000000";
					when "11010001100111111" => rgb <= "000000";
					when "11010010000000000" => rgb <= "000000";
					when "11010010000000001" => rgb <= "000000";
					when "11010010000000010" => rgb <= "000000";
					when "11010010000000011" => rgb <= "000000";
					when "11010010000000100" => rgb <= "000000";
					when "11010010000000101" => rgb <= "000000";
					when "11010010000000110" => rgb <= "000000";
					when "11010010000000111" => rgb <= "000000";
					when "11010010000001000" => rgb <= "000000";
					when "11010010000001001" => rgb <= "000000";
					when "11010010000001010" => rgb <= "000000";
					when "11010010000001011" => rgb <= "000000";
					when "11010010000001100" => rgb <= "000000";
					when "11010010000001101" => rgb <= "000000";
					when "11010010000001110" => rgb <= "000000";
					when "11010010000001111" => rgb <= "000000";
					when "11010010000010000" => rgb <= "000000";
					when "11010010000010001" => rgb <= "000000";
					when "11010010000010010" => rgb <= "000000";
					when "11010010000010011" => rgb <= "000000";
					when "11010010000010100" => rgb <= "101010";
					when "11010010000010101" => rgb <= "111111";
					when "11010010000010110" => rgb <= "101010";
					when "11010010000010111" => rgb <= "111111";
					when "11010010000011000" => rgb <= "101010";
					when "11010010000011001" => rgb <= "111111";
					when "11010010000011010" => rgb <= "111111";
					when "11010010000011011" => rgb <= "111111";
					when "11010010000011100" => rgb <= "101010";
					when "11010010000011101" => rgb <= "111111";
					when "11010010000011110" => rgb <= "111111";
					when "11010010000011111" => rgb <= "111111";
					when "11010010000100000" => rgb <= "111111";
					when "11010010000100001" => rgb <= "101010";
					when "11010010000100010" => rgb <= "111111";
					when "11010010000100011" => rgb <= "000000";
					when "11010010000100100" => rgb <= "000000";
					when "11010010000100101" => rgb <= "000000";
					when "11010010000100110" => rgb <= "000000";
					when "11010010000100111" => rgb <= "000000";
					when "11010010000101000" => rgb <= "000000";
					when "11010010000101001" => rgb <= "000000";
					when "11010010000101010" => rgb <= "000000";
					when "11010010000101011" => rgb <= "000000";
					when "11010010000101100" => rgb <= "000000";
					when "11010010000101101" => rgb <= "000000";
					when "11010010000101110" => rgb <= "000000";
					when "11010010000101111" => rgb <= "000000";
					when "11010010000110000" => rgb <= "000000";
					when "11010010000110001" => rgb <= "000000";
					when "11010010000110010" => rgb <= "000000";
					when "11010010000110011" => rgb <= "000000";
					when "11010010000110100" => rgb <= "000000";
					when "11010010000110101" => rgb <= "000000";
					when "11010010000110110" => rgb <= "000000";
					when "11010010000110111" => rgb <= "000000";
					when "11010010000111000" => rgb <= "000000";
					when "11010010000111001" => rgb <= "000000";
					when "11010010000111010" => rgb <= "000000";
					when "11010010000111011" => rgb <= "000000";
					when "11010010000111100" => rgb <= "000000";
					when "11010010000111101" => rgb <= "000000";
					when "11010010000111110" => rgb <= "000000";
					when "11010010000111111" => rgb <= "000000";
					when "11010010001000000" => rgb <= "000000";
					when "11010010001000001" => rgb <= "101010";
					when "11010010001000010" => rgb <= "101010";
					when "11010010001000011" => rgb <= "111111";
					when "11010010001000100" => rgb <= "111111";
					when "11010010001000101" => rgb <= "111111";
					when "11010010001000110" => rgb <= "101010";
					when "11010010001000111" => rgb <= "111111";
					when "11010010001001000" => rgb <= "111111";
					when "11010010001001001" => rgb <= "111111";
					when "11010010001001010" => rgb <= "111111";
					when "11010010001001011" => rgb <= "111111";
					when "11010010001001100" => rgb <= "111111";
					when "11010010001001101" => rgb <= "111111";
					when "11010010001001110" => rgb <= "111111";
					when "11010010001001111" => rgb <= "111111";
					when "11010010001010000" => rgb <= "111111";
					when "11010010001010001" => rgb <= "111111";
					when "11010010001010010" => rgb <= "111111";
					when "11010010001010011" => rgb <= "101010";
					when "11010010001010100" => rgb <= "111111";
					when "11010010001010101" => rgb <= "101010";
					when "11010010001010110" => rgb <= "111111";
					when "11010010001010111" => rgb <= "101010";
					when "11010010001011000" => rgb <= "000000";
					when "11010010001011001" => rgb <= "000000";
					when "11010010001011010" => rgb <= "000000";
					when "11010010001011011" => rgb <= "000000";
					when "11010010001011100" => rgb <= "000000";
					when "11010010001011101" => rgb <= "000000";
					when "11010010001011110" => rgb <= "000000";
					when "11010010001011111" => rgb <= "000000";
					when "11010010001100000" => rgb <= "000000";
					when "11010010001100001" => rgb <= "000000";
					when "11010010001100010" => rgb <= "000000";
					when "11010010001100011" => rgb <= "000000";
					when "11010010001100100" => rgb <= "000000";
					when "11010010001100101" => rgb <= "000000";
					when "11010010001100110" => rgb <= "000000";
					when "11010010001100111" => rgb <= "000000";
					when "11010010001101000" => rgb <= "000000";
					when "11010010001101001" => rgb <= "000000";
					when "11010010001101010" => rgb <= "000000";
					when "11010010001101011" => rgb <= "000000";
					when "11010010001101100" => rgb <= "000000";
					when "11010010001101101" => rgb <= "000000";
					when "11010010001101110" => rgb <= "101010";
					when "11010010001101111" => rgb <= "101010";
					when "11010010001110000" => rgb <= "101010";
					when "11010010001110001" => rgb <= "111111";
					when "11010010001110010" => rgb <= "111111";
					when "11010010001110011" => rgb <= "111111";
					when "11010010001110100" => rgb <= "111111";
					when "11010010001110101" => rgb <= "111111";
					when "11010010001110110" => rgb <= "111111";
					when "11010010001110111" => rgb <= "111111";
					when "11010010001111000" => rgb <= "111111";
					when "11010010001111001" => rgb <= "111111";
					when "11010010001111010" => rgb <= "111111";
					when "11010010001111011" => rgb <= "111111";
					when "11010010001111100" => rgb <= "111111";
					when "11010010001111101" => rgb <= "111111";
					when "11010010001111110" => rgb <= "111111";
					when "11010010001111111" => rgb <= "111111";
					when "11010010010000000" => rgb <= "111111";
					when "11010010010000001" => rgb <= "111111";
					when "11010010010000010" => rgb <= "101010";
					when "11010010010000011" => rgb <= "101010";
					when "11010010010000100" => rgb <= "101010";
					when "11010010010000101" => rgb <= "000000";
					when "11010010010000110" => rgb <= "000000";
					when "11010010010000111" => rgb <= "000000";
					when "11010010010001000" => rgb <= "000000";
					when "11010010010001001" => rgb <= "000000";
					when "11010010010001010" => rgb <= "000000";
					when "11010010010001011" => rgb <= "000000";
					when "11010010010001100" => rgb <= "000000";
					when "11010010010001101" => rgb <= "000000";
					when "11010010010001110" => rgb <= "000000";
					when "11010010010001111" => rgb <= "000000";
					when "11010010010010000" => rgb <= "000000";
					when "11010010010010001" => rgb <= "000000";
					when "11010010010010010" => rgb <= "000000";
					when "11010010010010011" => rgb <= "000000";
					when "11010010010010100" => rgb <= "000000";
					when "11010010010010101" => rgb <= "000000";
					when "11010010010010110" => rgb <= "000000";
					when "11010010010010111" => rgb <= "000000";
					when "11010010010011000" => rgb <= "000000";
					when "11010010010011001" => rgb <= "000000";
					when "11010010010011010" => rgb <= "000000";
					when "11010010010011011" => rgb <= "000000";
					when "11010010010011100" => rgb <= "000000";
					when "11010010010011101" => rgb <= "000000";
					when "11010010010011110" => rgb <= "000000";
					when "11010010010011111" => rgb <= "000000";
					when "11010010010100000" => rgb <= "000000";
					when "11010010010100001" => rgb <= "000000";
					when "11010010010100010" => rgb <= "000000";
					when "11010010010100011" => rgb <= "000000";
					when "11010010010100100" => rgb <= "000000";
					when "11010010010100101" => rgb <= "000000";
					when "11010010010100110" => rgb <= "000000";
					when "11010010010100111" => rgb <= "000000";
					when "11010010010101000" => rgb <= "000000";
					when "11010010010101001" => rgb <= "000000";
					when "11010010010101010" => rgb <= "101010";
					when "11010010010101011" => rgb <= "101010";
					when "11010010010101100" => rgb <= "101010";
					when "11010010010101101" => rgb <= "101010";
					when "11010010010101110" => rgb <= "111111";
					when "11010010010101111" => rgb <= "101010";
					when "11010010010110000" => rgb <= "101010";
					when "11010010010110001" => rgb <= "101010";
					when "11010010010110010" => rgb <= "000000";
					when "11010010010110011" => rgb <= "000000";
					when "11010010010110100" => rgb <= "000000";
					when "11010010010110101" => rgb <= "000000";
					when "11010010010110110" => rgb <= "000000";
					when "11010010010110111" => rgb <= "000000";
					when "11010010010111000" => rgb <= "000000";
					when "11010010010111001" => rgb <= "101010";
					when "11010010010111010" => rgb <= "101010";
					when "11010010010111011" => rgb <= "101010";
					when "11010010010111100" => rgb <= "111111";
					when "11010010010111101" => rgb <= "101010";
					when "11010010010111110" => rgb <= "101010";
					when "11010010010111111" => rgb <= "111111";
					when "11010010011000000" => rgb <= "111111";
					when "11010010011000001" => rgb <= "111111";
					when "11010010011000010" => rgb <= "111111";
					when "11010010011000011" => rgb <= "111111";
					when "11010010011000100" => rgb <= "111111";
					when "11010010011000101" => rgb <= "111111";
					when "11010010011000110" => rgb <= "111111";
					when "11010010011000111" => rgb <= "111111";
					when "11010010011001000" => rgb <= "000000";
					when "11010010011001001" => rgb <= "000000";
					when "11010010011001010" => rgb <= "000000";
					when "11010010011001011" => rgb <= "000000";
					when "11010010011001100" => rgb <= "000000";
					when "11010010011001101" => rgb <= "000000";
					when "11010010011001110" => rgb <= "000000";
					when "11010010011001111" => rgb <= "000000";
					when "11010010011010000" => rgb <= "000000";
					when "11010010011010001" => rgb <= "000000";
					when "11010010011010010" => rgb <= "000000";
					when "11010010011010011" => rgb <= "000000";
					when "11010010011010100" => rgb <= "000000";
					when "11010010011010101" => rgb <= "000000";
					when "11010010011010110" => rgb <= "000000";
					when "11010010011010111" => rgb <= "101010";
					when "11010010011011000" => rgb <= "111111";
					when "11010010011011001" => rgb <= "111111";
					when "11010010011011010" => rgb <= "111111";
					when "11010010011011011" => rgb <= "111111";
					when "11010010011011100" => rgb <= "111111";
					when "11010010011011101" => rgb <= "111111";
					when "11010010011011110" => rgb <= "111111";
					when "11010010011011111" => rgb <= "111111";
					when "11010010011100000" => rgb <= "101010";
					when "11010010011100001" => rgb <= "101010";
					when "11010010011100010" => rgb <= "111111";
					when "11010010011100011" => rgb <= "111111";
					when "11010010011100100" => rgb <= "101010";
					when "11010010011100101" => rgb <= "111111";
					when "11010010011100110" => rgb <= "000000";
					when "11010010011100111" => rgb <= "000000";
					when "11010010011101000" => rgb <= "000000";
					when "11010010011101001" => rgb <= "000000";
					when "11010010011101010" => rgb <= "000000";
					when "11010010011101011" => rgb <= "000000";
					when "11010010011101100" => rgb <= "000000";
					when "11010010011101101" => rgb <= "010101";
					when "11010010011101110" => rgb <= "111111";
					when "11010010011101111" => rgb <= "101010";
					when "11010010011110000" => rgb <= "111111";
					when "11010010011110001" => rgb <= "111111";
					when "11010010011110010" => rgb <= "111111";
					when "11010010011110011" => rgb <= "101010";
					when "11010010011110100" => rgb <= "101010";
					when "11010010011110101" => rgb <= "000000";
					when "11010010011110110" => rgb <= "000000";
					when "11010010011110111" => rgb <= "000000";
					when "11010010011111000" => rgb <= "000000";
					when "11010010011111001" => rgb <= "000000";
					when "11010010011111010" => rgb <= "000000";
					when "11010010011111011" => rgb <= "000000";
					when "11010010011111100" => rgb <= "000000";
					when "11010010011111101" => rgb <= "000000";
					when "11010010011111110" => rgb <= "000000";
					when "11010010011111111" => rgb <= "000000";
					when "11010010100000000" => rgb <= "000000";
					when "11010010100000001" => rgb <= "000000";
					when "11010010100000010" => rgb <= "000000";
					when "11010010100000011" => rgb <= "000000";
					when "11010010100000100" => rgb <= "000000";
					when "11010010100000101" => rgb <= "000000";
					when "11010010100000110" => rgb <= "000000";
					when "11010010100000111" => rgb <= "000000";
					when "11010010100001000" => rgb <= "000000";
					when "11010010100001001" => rgb <= "000000";
					when "11010010100001010" => rgb <= "000000";
					when "11010010100001011" => rgb <= "010101";
					when "11010010100001100" => rgb <= "111111";
					when "11010010100001101" => rgb <= "101010";
					when "11010010100001110" => rgb <= "111111";
					when "11010010100001111" => rgb <= "111111";
					when "11010010100010000" => rgb <= "111111";
					when "11010010100010001" => rgb <= "111111";
					when "11010010100010010" => rgb <= "111111";
					when "11010010100010011" => rgb <= "111111";
					when "11010010100010100" => rgb <= "111111";
					when "11010010100010101" => rgb <= "111111";
					when "11010010100010110" => rgb <= "111111";
					when "11010010100010111" => rgb <= "111111";
					when "11010010100011000" => rgb <= "101010";
					when "11010010100011001" => rgb <= "111111";
					when "11010010100011010" => rgb <= "101010";
					when "11010010100011011" => rgb <= "000000";
					when "11010010100011100" => rgb <= "000000";
					when "11010010100011101" => rgb <= "000000";
					when "11010010100011110" => rgb <= "000000";
					when "11010010100011111" => rgb <= "000000";
					when "11010010100100000" => rgb <= "000000";
					when "11010010100100001" => rgb <= "000000";
					when "11010010100100010" => rgb <= "101010";
					when "11010010100100011" => rgb <= "101010";
					when "11010010100100100" => rgb <= "101010";
					when "11010010100100101" => rgb <= "111111";
					when "11010010100100110" => rgb <= "111111";
					when "11010010100100111" => rgb <= "111111";
					when "11010010100101000" => rgb <= "111111";
					when "11010010100101001" => rgb <= "111111";
					when "11010010100101010" => rgb <= "111111";
					when "11010010100101011" => rgb <= "111111";
					when "11010010100101100" => rgb <= "111111";
					when "11010010100101101" => rgb <= "111111";
					when "11010010100101110" => rgb <= "101010";
					when "11010010100101111" => rgb <= "101010";
					when "11010010100110000" => rgb <= "111111";
					when "11010010100110001" => rgb <= "000000";
					when "11010010100110010" => rgb <= "000000";
					when "11010010100110011" => rgb <= "000000";
					when "11010010100110100" => rgb <= "000000";
					when "11010010100110101" => rgb <= "000000";
					when "11010010100110110" => rgb <= "000000";
					when "11010010100110111" => rgb <= "000000";
					when "11010010100111000" => rgb <= "000000";
					when "11010010100111001" => rgb <= "000000";
					when "11010010100111010" => rgb <= "000000";
					when "11010010100111011" => rgb <= "000000";
					when "11010010100111100" => rgb <= "000000";
					when "11010010100111101" => rgb <= "000000";
					when "11010010100111110" => rgb <= "000000";
					when "11010010100111111" => rgb <= "000000";
					when "11010011000000000" => rgb <= "000000";
					when "11010011000000001" => rgb <= "000000";
					when "11010011000000010" => rgb <= "000000";
					when "11010011000000011" => rgb <= "000000";
					when "11010011000000100" => rgb <= "000000";
					when "11010011000000101" => rgb <= "000000";
					when "11010011000000110" => rgb <= "000000";
					when "11010011000000111" => rgb <= "000000";
					when "11010011000001000" => rgb <= "000000";
					when "11010011000001001" => rgb <= "000000";
					when "11010011000001010" => rgb <= "000000";
					when "11010011000001011" => rgb <= "000000";
					when "11010011000001100" => rgb <= "000000";
					when "11010011000001101" => rgb <= "000000";
					when "11010011000001110" => rgb <= "000000";
					when "11010011000001111" => rgb <= "000000";
					when "11010011000010000" => rgb <= "000000";
					when "11010011000010001" => rgb <= "000000";
					when "11010011000010010" => rgb <= "000000";
					when "11010011000010011" => rgb <= "000000";
					when "11010011000010100" => rgb <= "101010";
					when "11010011000010101" => rgb <= "111111";
					when "11010011000010110" => rgb <= "101010";
					when "11010011000010111" => rgb <= "101010";
					when "11010011000011000" => rgb <= "101010";
					when "11010011000011001" => rgb <= "101010";
					when "11010011000011010" => rgb <= "101010";
					when "11010011000011011" => rgb <= "101010";
					when "11010011000011100" => rgb <= "101010";
					when "11010011000011101" => rgb <= "101010";
					when "11010011000011110" => rgb <= "101010";
					when "11010011000011111" => rgb <= "101010";
					when "11010011000100000" => rgb <= "101010";
					when "11010011000100001" => rgb <= "101010";
					when "11010011000100010" => rgb <= "111111";
					when "11010011000100011" => rgb <= "000000";
					when "11010011000100100" => rgb <= "000000";
					when "11010011000100101" => rgb <= "000000";
					when "11010011000100110" => rgb <= "000000";
					when "11010011000100111" => rgb <= "000000";
					when "11010011000101000" => rgb <= "000000";
					when "11010011000101001" => rgb <= "000000";
					when "11010011000101010" => rgb <= "000000";
					when "11010011000101011" => rgb <= "000000";
					when "11010011000101100" => rgb <= "000000";
					when "11010011000101101" => rgb <= "000000";
					when "11010011000101110" => rgb <= "000000";
					when "11010011000101111" => rgb <= "000000";
					when "11010011000110000" => rgb <= "000000";
					when "11010011000110001" => rgb <= "000000";
					when "11010011000110010" => rgb <= "000000";
					when "11010011000110011" => rgb <= "000000";
					when "11010011000110100" => rgb <= "000000";
					when "11010011000110101" => rgb <= "000000";
					when "11010011000110110" => rgb <= "000000";
					when "11010011000110111" => rgb <= "000000";
					when "11010011000111000" => rgb <= "000000";
					when "11010011000111001" => rgb <= "000000";
					when "11010011000111010" => rgb <= "000000";
					when "11010011000111011" => rgb <= "000000";
					when "11010011000111100" => rgb <= "000000";
					when "11010011000111101" => rgb <= "000000";
					when "11010011000111110" => rgb <= "000000";
					when "11010011000111111" => rgb <= "000000";
					when "11010011001000000" => rgb <= "000000";
					when "11010011001000001" => rgb <= "101010";
					when "11010011001000010" => rgb <= "101010";
					when "11010011001000011" => rgb <= "111111";
					when "11010011001000100" => rgb <= "101010";
					when "11010011001000101" => rgb <= "101010";
					when "11010011001000110" => rgb <= "101010";
					when "11010011001000111" => rgb <= "101010";
					when "11010011001001000" => rgb <= "101010";
					when "11010011001001001" => rgb <= "101010";
					when "11010011001001010" => rgb <= "101010";
					when "11010011001001011" => rgb <= "101010";
					when "11010011001001100" => rgb <= "101010";
					when "11010011001001101" => rgb <= "101010";
					when "11010011001001110" => rgb <= "101010";
					when "11010011001001111" => rgb <= "101010";
					when "11010011001010000" => rgb <= "101010";
					when "11010011001010001" => rgb <= "101010";
					when "11010011001010010" => rgb <= "101010";
					when "11010011001010011" => rgb <= "101010";
					when "11010011001010100" => rgb <= "101010";
					when "11010011001010101" => rgb <= "101010";
					when "11010011001010110" => rgb <= "111111";
					when "11010011001010111" => rgb <= "010101";
					when "11010011001011000" => rgb <= "000000";
					when "11010011001011001" => rgb <= "000000";
					when "11010011001011010" => rgb <= "000000";
					when "11010011001011011" => rgb <= "000000";
					when "11010011001011100" => rgb <= "000000";
					when "11010011001011101" => rgb <= "000000";
					when "11010011001011110" => rgb <= "000000";
					when "11010011001011111" => rgb <= "000000";
					when "11010011001100000" => rgb <= "000000";
					when "11010011001100001" => rgb <= "000000";
					when "11010011001100010" => rgb <= "000000";
					when "11010011001100011" => rgb <= "000000";
					when "11010011001100100" => rgb <= "000000";
					when "11010011001100101" => rgb <= "000000";
					when "11010011001100110" => rgb <= "000000";
					when "11010011001100111" => rgb <= "000000";
					when "11010011001101000" => rgb <= "000000";
					when "11010011001101001" => rgb <= "000000";
					when "11010011001101010" => rgb <= "000000";
					when "11010011001101011" => rgb <= "000000";
					when "11010011001101100" => rgb <= "000000";
					when "11010011001101101" => rgb <= "000000";
					when "11010011001101110" => rgb <= "101010";
					when "11010011001101111" => rgb <= "111111";
					when "11010011001110000" => rgb <= "101010";
					when "11010011001110001" => rgb <= "101010";
					when "11010011001110010" => rgb <= "101010";
					when "11010011001110011" => rgb <= "101010";
					when "11010011001110100" => rgb <= "101010";
					when "11010011001110101" => rgb <= "101010";
					when "11010011001110110" => rgb <= "101010";
					when "11010011001110111" => rgb <= "101010";
					when "11010011001111000" => rgb <= "101010";
					when "11010011001111001" => rgb <= "101010";
					when "11010011001111010" => rgb <= "101010";
					when "11010011001111011" => rgb <= "101010";
					when "11010011001111100" => rgb <= "101010";
					when "11010011001111101" => rgb <= "101010";
					when "11010011001111110" => rgb <= "101010";
					when "11010011001111111" => rgb <= "101010";
					when "11010011010000000" => rgb <= "101010";
					when "11010011010000001" => rgb <= "101010";
					when "11010011010000010" => rgb <= "101010";
					when "11010011010000011" => rgb <= "101010";
					when "11010011010000100" => rgb <= "101010";
					when "11010011010000101" => rgb <= "000000";
					when "11010011010000110" => rgb <= "000000";
					when "11010011010000111" => rgb <= "000000";
					when "11010011010001000" => rgb <= "000000";
					when "11010011010001001" => rgb <= "000000";
					when "11010011010001010" => rgb <= "000000";
					when "11010011010001011" => rgb <= "000000";
					when "11010011010001100" => rgb <= "000000";
					when "11010011010001101" => rgb <= "000000";
					when "11010011010001110" => rgb <= "000000";
					when "11010011010001111" => rgb <= "000000";
					when "11010011010010000" => rgb <= "000000";
					when "11010011010010001" => rgb <= "000000";
					when "11010011010010010" => rgb <= "000000";
					when "11010011010010011" => rgb <= "000000";
					when "11010011010010100" => rgb <= "000000";
					when "11010011010010101" => rgb <= "000000";
					when "11010011010010110" => rgb <= "000000";
					when "11010011010010111" => rgb <= "000000";
					when "11010011010011000" => rgb <= "000000";
					when "11010011010011001" => rgb <= "000000";
					when "11010011010011010" => rgb <= "000000";
					when "11010011010011011" => rgb <= "000000";
					when "11010011010011100" => rgb <= "000000";
					when "11010011010011101" => rgb <= "000000";
					when "11010011010011110" => rgb <= "000000";
					when "11010011010011111" => rgb <= "000000";
					when "11010011010100000" => rgb <= "000000";
					when "11010011010100001" => rgb <= "000000";
					when "11010011010100010" => rgb <= "000000";
					when "11010011010100011" => rgb <= "000000";
					when "11010011010100100" => rgb <= "000000";
					when "11010011010100101" => rgb <= "000000";
					when "11010011010100110" => rgb <= "000000";
					when "11010011010100111" => rgb <= "000000";
					when "11010011010101000" => rgb <= "000000";
					when "11010011010101001" => rgb <= "000000";
					when "11010011010101010" => rgb <= "101010";
					when "11010011010101011" => rgb <= "101010";
					when "11010011010101100" => rgb <= "101010";
					when "11010011010101101" => rgb <= "101010";
					when "11010011010101110" => rgb <= "111111";
					when "11010011010101111" => rgb <= "101010";
					when "11010011010110000" => rgb <= "111111";
					when "11010011010110001" => rgb <= "101010";
					when "11010011010110010" => rgb <= "000000";
					when "11010011010110011" => rgb <= "000000";
					when "11010011010110100" => rgb <= "000000";
					when "11010011010110101" => rgb <= "000000";
					when "11010011010110110" => rgb <= "000000";
					when "11010011010110111" => rgb <= "000000";
					when "11010011010111000" => rgb <= "000000";
					when "11010011010111001" => rgb <= "101010";
					when "11010011010111010" => rgb <= "101010";
					when "11010011010111011" => rgb <= "101010";
					when "11010011010111100" => rgb <= "101010";
					when "11010011010111101" => rgb <= "101010";
					when "11010011010111110" => rgb <= "101010";
					when "11010011010111111" => rgb <= "111111";
					when "11010011011000000" => rgb <= "101010";
					when "11010011011000001" => rgb <= "101010";
					when "11010011011000010" => rgb <= "101010";
					when "11010011011000011" => rgb <= "101010";
					when "11010011011000100" => rgb <= "101010";
					when "11010011011000101" => rgb <= "101010";
					when "11010011011000110" => rgb <= "101010";
					when "11010011011000111" => rgb <= "101010";
					when "11010011011001000" => rgb <= "000000";
					when "11010011011001001" => rgb <= "000000";
					when "11010011011001010" => rgb <= "000000";
					when "11010011011001011" => rgb <= "000000";
					when "11010011011001100" => rgb <= "000000";
					when "11010011011001101" => rgb <= "000000";
					when "11010011011001110" => rgb <= "000000";
					when "11010011011001111" => rgb <= "000000";
					when "11010011011010000" => rgb <= "000000";
					when "11010011011010001" => rgb <= "000000";
					when "11010011011010010" => rgb <= "000000";
					when "11010011011010011" => rgb <= "000000";
					when "11010011011010100" => rgb <= "000000";
					when "11010011011010101" => rgb <= "000000";
					when "11010011011010110" => rgb <= "000000";
					when "11010011011010111" => rgb <= "101010";
					when "11010011011011000" => rgb <= "101010";
					when "11010011011011001" => rgb <= "101010";
					when "11010011011011010" => rgb <= "101010";
					when "11010011011011011" => rgb <= "101010";
					when "11010011011011100" => rgb <= "101010";
					when "11010011011011101" => rgb <= "101010";
					when "11010011011011110" => rgb <= "101010";
					when "11010011011011111" => rgb <= "101010";
					when "11010011011100000" => rgb <= "111111";
					when "11010011011100001" => rgb <= "101010";
					when "11010011011100010" => rgb <= "101010";
					when "11010011011100011" => rgb <= "101010";
					when "11010011011100100" => rgb <= "101010";
					when "11010011011100101" => rgb <= "111111";
					when "11010011011100110" => rgb <= "000000";
					when "11010011011100111" => rgb <= "000000";
					when "11010011011101000" => rgb <= "000000";
					when "11010011011101001" => rgb <= "000000";
					when "11010011011101010" => rgb <= "000000";
					when "11010011011101011" => rgb <= "000000";
					when "11010011011101100" => rgb <= "000000";
					when "11010011011101101" => rgb <= "010101";
					when "11010011011101110" => rgb <= "111111";
					when "11010011011101111" => rgb <= "101010";
					when "11010011011110000" => rgb <= "101010";
					when "11010011011110001" => rgb <= "101010";
					when "11010011011110010" => rgb <= "101010";
					when "11010011011110011" => rgb <= "101010";
					when "11010011011110100" => rgb <= "101010";
					when "11010011011110101" => rgb <= "000000";
					when "11010011011110110" => rgb <= "000000";
					when "11010011011110111" => rgb <= "000000";
					when "11010011011111000" => rgb <= "000000";
					when "11010011011111001" => rgb <= "000000";
					when "11010011011111010" => rgb <= "000000";
					when "11010011011111011" => rgb <= "000000";
					when "11010011011111100" => rgb <= "000000";
					when "11010011011111101" => rgb <= "000000";
					when "11010011011111110" => rgb <= "000000";
					when "11010011011111111" => rgb <= "000000";
					when "11010011100000000" => rgb <= "000000";
					when "11010011100000001" => rgb <= "000000";
					when "11010011100000010" => rgb <= "000000";
					when "11010011100000011" => rgb <= "000000";
					when "11010011100000100" => rgb <= "000000";
					when "11010011100000101" => rgb <= "000000";
					when "11010011100000110" => rgb <= "000000";
					when "11010011100000111" => rgb <= "000000";
					when "11010011100001000" => rgb <= "000000";
					when "11010011100001001" => rgb <= "000000";
					when "11010011100001010" => rgb <= "000000";
					when "11010011100001011" => rgb <= "010101";
					when "11010011100001100" => rgb <= "111111";
					when "11010011100001101" => rgb <= "101010";
					when "11010011100001110" => rgb <= "101010";
					when "11010011100001111" => rgb <= "101010";
					when "11010011100010000" => rgb <= "101010";
					when "11010011100010001" => rgb <= "101010";
					when "11010011100010010" => rgb <= "101010";
					when "11010011100010011" => rgb <= "101010";
					when "11010011100010100" => rgb <= "101010";
					when "11010011100010101" => rgb <= "101010";
					when "11010011100010110" => rgb <= "101010";
					when "11010011100010111" => rgb <= "101010";
					when "11010011100011000" => rgb <= "101010";
					when "11010011100011001" => rgb <= "101010";
					when "11010011100011010" => rgb <= "101010";
					when "11010011100011011" => rgb <= "000000";
					when "11010011100011100" => rgb <= "000000";
					when "11010011100011101" => rgb <= "000000";
					when "11010011100011110" => rgb <= "000000";
					when "11010011100011111" => rgb <= "000000";
					when "11010011100100000" => rgb <= "000000";
					when "11010011100100001" => rgb <= "000000";
					when "11010011100100010" => rgb <= "101010";
					when "11010011100100011" => rgb <= "101010";
					when "11010011100100100" => rgb <= "101010";
					when "11010011100100101" => rgb <= "101010";
					when "11010011100100110" => rgb <= "101010";
					when "11010011100100111" => rgb <= "101010";
					when "11010011100101000" => rgb <= "101010";
					when "11010011100101001" => rgb <= "101010";
					when "11010011100101010" => rgb <= "101010";
					when "11010011100101011" => rgb <= "101010";
					when "11010011100101100" => rgb <= "101010";
					when "11010011100101101" => rgb <= "101010";
					when "11010011100101110" => rgb <= "101010";
					when "11010011100101111" => rgb <= "101010";
					when "11010011100110000" => rgb <= "111111";
					when "11010011100110001" => rgb <= "000000";
					when "11010011100110010" => rgb <= "000000";
					when "11010011100110011" => rgb <= "000000";
					when "11010011100110100" => rgb <= "000000";
					when "11010011100110101" => rgb <= "000000";
					when "11010011100110110" => rgb <= "000000";
					when "11010011100110111" => rgb <= "000000";
					when "11010011100111000" => rgb <= "000000";
					when "11010011100111001" => rgb <= "000000";
					when "11010011100111010" => rgb <= "000000";
					when "11010011100111011" => rgb <= "000000";
					when "11010011100111100" => rgb <= "000000";
					when "11010011100111101" => rgb <= "000000";
					when "11010011100111110" => rgb <= "000000";
					when "11010011100111111" => rgb <= "000000";
					when "11010100000000000" => rgb <= "000000";
					when "11010100000000001" => rgb <= "000000";
					when "11010100000000010" => rgb <= "000000";
					when "11010100000000011" => rgb <= "000000";
					when "11010100000000100" => rgb <= "000000";
					when "11010100000000101" => rgb <= "000000";
					when "11010100000000110" => rgb <= "000000";
					when "11010100000000111" => rgb <= "000000";
					when "11010100000001000" => rgb <= "000000";
					when "11010100000001001" => rgb <= "000000";
					when "11010100000001010" => rgb <= "000000";
					when "11010100000001011" => rgb <= "000000";
					when "11010100000001100" => rgb <= "000000";
					when "11010100000001101" => rgb <= "000000";
					when "11010100000001110" => rgb <= "000000";
					when "11010100000001111" => rgb <= "000000";
					when "11010100000010000" => rgb <= "000000";
					when "11010100000010001" => rgb <= "000000";
					when "11010100000010010" => rgb <= "000000";
					when "11010100000010011" => rgb <= "000000";
					when "11010100000010100" => rgb <= "101010";
					when "11010100000010101" => rgb <= "111111";
					when "11010100000010110" => rgb <= "111111";
					when "11010100000010111" => rgb <= "111111";
					when "11010100000011000" => rgb <= "111111";
					when "11010100000011001" => rgb <= "101010";
					when "11010100000011010" => rgb <= "111111";
					when "11010100000011011" => rgb <= "111111";
					when "11010100000011100" => rgb <= "111111";
					when "11010100000011101" => rgb <= "111111";
					when "11010100000011110" => rgb <= "111111";
					when "11010100000011111" => rgb <= "111111";
					when "11010100000100000" => rgb <= "111111";
					when "11010100000100001" => rgb <= "111111";
					when "11010100000100010" => rgb <= "111111";
					when "11010100000100011" => rgb <= "000000";
					when "11010100000100100" => rgb <= "000000";
					when "11010100000100101" => rgb <= "000000";
					when "11010100000100110" => rgb <= "000000";
					when "11010100000100111" => rgb <= "000000";
					when "11010100000101000" => rgb <= "000000";
					when "11010100000101001" => rgb <= "000000";
					when "11010100000101010" => rgb <= "000000";
					when "11010100000101011" => rgb <= "000000";
					when "11010100000101100" => rgb <= "000000";
					when "11010100000101101" => rgb <= "000000";
					when "11010100000101110" => rgb <= "000000";
					when "11010100000101111" => rgb <= "000000";
					when "11010100000110000" => rgb <= "000000";
					when "11010100000110001" => rgb <= "000000";
					when "11010100000110010" => rgb <= "000000";
					when "11010100000110011" => rgb <= "000000";
					when "11010100000110100" => rgb <= "000000";
					when "11010100000110101" => rgb <= "000000";
					when "11010100000110110" => rgb <= "000000";
					when "11010100000110111" => rgb <= "000000";
					when "11010100000111000" => rgb <= "000000";
					when "11010100000111001" => rgb <= "000000";
					when "11010100000111010" => rgb <= "000000";
					when "11010100000111011" => rgb <= "000000";
					when "11010100000111100" => rgb <= "000000";
					when "11010100000111101" => rgb <= "000000";
					when "11010100000111110" => rgb <= "000000";
					when "11010100000111111" => rgb <= "000000";
					when "11010100001000000" => rgb <= "000000";
					when "11010100001000001" => rgb <= "101010";
					when "11010100001000010" => rgb <= "111111";
					when "11010100001000011" => rgb <= "101010";
					when "11010100001000100" => rgb <= "111111";
					when "11010100001000101" => rgb <= "111111";
					when "11010100001000110" => rgb <= "101010";
					when "11010100001000111" => rgb <= "111111";
					when "11010100001001000" => rgb <= "111111";
					when "11010100001001001" => rgb <= "111111";
					when "11010100001001010" => rgb <= "111111";
					when "11010100001001011" => rgb <= "101010";
					when "11010100001001100" => rgb <= "111111";
					when "11010100001001101" => rgb <= "111111";
					when "11010100001001110" => rgb <= "111111";
					when "11010100001001111" => rgb <= "111111";
					when "11010100001010000" => rgb <= "111111";
					when "11010100001010001" => rgb <= "101010";
					when "11010100001010010" => rgb <= "111111";
					when "11010100001010011" => rgb <= "101010";
					when "11010100001010100" => rgb <= "111111";
					when "11010100001010101" => rgb <= "111111";
					when "11010100001010110" => rgb <= "111111";
					when "11010100001010111" => rgb <= "101010";
					when "11010100001011000" => rgb <= "000000";
					when "11010100001011001" => rgb <= "000000";
					when "11010100001011010" => rgb <= "000000";
					when "11010100001011011" => rgb <= "000000";
					when "11010100001011100" => rgb <= "000000";
					when "11010100001011101" => rgb <= "000000";
					when "11010100001011110" => rgb <= "000000";
					when "11010100001011111" => rgb <= "000000";
					when "11010100001100000" => rgb <= "000000";
					when "11010100001100001" => rgb <= "000000";
					when "11010100001100010" => rgb <= "000000";
					when "11010100001100011" => rgb <= "000000";
					when "11010100001100100" => rgb <= "000000";
					when "11010100001100101" => rgb <= "000000";
					when "11010100001100110" => rgb <= "000000";
					when "11010100001100111" => rgb <= "000000";
					when "11010100001101000" => rgb <= "000000";
					when "11010100001101001" => rgb <= "000000";
					when "11010100001101010" => rgb <= "000000";
					when "11010100001101011" => rgb <= "000000";
					when "11010100001101100" => rgb <= "000000";
					when "11010100001101101" => rgb <= "000000";
					when "11010100001101110" => rgb <= "101010";
					when "11010100001101111" => rgb <= "111111";
					when "11010100001110000" => rgb <= "111111";
					when "11010100001110001" => rgb <= "111111";
					when "11010100001110010" => rgb <= "111111";
					when "11010100001110011" => rgb <= "111111";
					when "11010100001110100" => rgb <= "111111";
					when "11010100001110101" => rgb <= "111111";
					when "11010100001110110" => rgb <= "111111";
					when "11010100001110111" => rgb <= "111111";
					when "11010100001111000" => rgb <= "111111";
					when "11010100001111001" => rgb <= "111111";
					when "11010100001111010" => rgb <= "111111";
					when "11010100001111011" => rgb <= "111111";
					when "11010100001111100" => rgb <= "111111";
					when "11010100001111101" => rgb <= "111111";
					when "11010100001111110" => rgb <= "111111";
					when "11010100001111111" => rgb <= "111111";
					when "11010100010000000" => rgb <= "111111";
					when "11010100010000001" => rgb <= "111111";
					when "11010100010000010" => rgb <= "111111";
					when "11010100010000011" => rgb <= "111111";
					when "11010100010000100" => rgb <= "101010";
					when "11010100010000101" => rgb <= "000000";
					when "11010100010000110" => rgb <= "000000";
					when "11010100010000111" => rgb <= "000000";
					when "11010100010001000" => rgb <= "000000";
					when "11010100010001001" => rgb <= "000000";
					when "11010100010001010" => rgb <= "000000";
					when "11010100010001011" => rgb <= "000000";
					when "11010100010001100" => rgb <= "000000";
					when "11010100010001101" => rgb <= "000000";
					when "11010100010001110" => rgb <= "000000";
					when "11010100010001111" => rgb <= "000000";
					when "11010100010010000" => rgb <= "000000";
					when "11010100010010001" => rgb <= "000000";
					when "11010100010010010" => rgb <= "000000";
					when "11010100010010011" => rgb <= "000000";
					when "11010100010010100" => rgb <= "000000";
					when "11010100010010101" => rgb <= "000000";
					when "11010100010010110" => rgb <= "000000";
					when "11010100010010111" => rgb <= "000000";
					when "11010100010011000" => rgb <= "000000";
					when "11010100010011001" => rgb <= "000000";
					when "11010100010011010" => rgb <= "000000";
					when "11010100010011011" => rgb <= "000000";
					when "11010100010011100" => rgb <= "000000";
					when "11010100010011101" => rgb <= "000000";
					when "11010100010011110" => rgb <= "000000";
					when "11010100010011111" => rgb <= "000000";
					when "11010100010100000" => rgb <= "000000";
					when "11010100010100001" => rgb <= "000000";
					when "11010100010100010" => rgb <= "000000";
					when "11010100010100011" => rgb <= "000000";
					when "11010100010100100" => rgb <= "000000";
					when "11010100010100101" => rgb <= "000000";
					when "11010100010100110" => rgb <= "000000";
					when "11010100010100111" => rgb <= "000000";
					when "11010100010101000" => rgb <= "000000";
					when "11010100010101001" => rgb <= "000000";
					when "11010100010101010" => rgb <= "101010";
					when "11010100010101011" => rgb <= "111111";
					when "11010100010101100" => rgb <= "111111";
					when "11010100010101101" => rgb <= "111111";
					when "11010100010101110" => rgb <= "101010";
					when "11010100010101111" => rgb <= "111111";
					when "11010100010110000" => rgb <= "101010";
					when "11010100010110001" => rgb <= "101010";
					when "11010100010110010" => rgb <= "000000";
					when "11010100010110011" => rgb <= "000000";
					when "11010100010110100" => rgb <= "000000";
					when "11010100010110101" => rgb <= "000000";
					when "11010100010110110" => rgb <= "000000";
					when "11010100010110111" => rgb <= "000000";
					when "11010100010111000" => rgb <= "000000";
					when "11010100010111001" => rgb <= "101010";
					when "11010100010111010" => rgb <= "111111";
					when "11010100010111011" => rgb <= "101010";
					when "11010100010111100" => rgb <= "111111";
					when "11010100010111101" => rgb <= "111111";
					when "11010100010111110" => rgb <= "101010";
					when "11010100010111111" => rgb <= "111111";
					when "11010100011000000" => rgb <= "111111";
					when "11010100011000001" => rgb <= "111111";
					when "11010100011000010" => rgb <= "111111";
					when "11010100011000011" => rgb <= "111111";
					when "11010100011000100" => rgb <= "111111";
					when "11010100011000101" => rgb <= "111111";
					when "11010100011000110" => rgb <= "111111";
					when "11010100011000111" => rgb <= "111111";
					when "11010100011001000" => rgb <= "000000";
					when "11010100011001001" => rgb <= "000000";
					when "11010100011001010" => rgb <= "000000";
					when "11010100011001011" => rgb <= "000000";
					when "11010100011001100" => rgb <= "000000";
					when "11010100011001101" => rgb <= "000000";
					when "11010100011001110" => rgb <= "000000";
					when "11010100011001111" => rgb <= "000000";
					when "11010100011010000" => rgb <= "000000";
					when "11010100011010001" => rgb <= "000000";
					when "11010100011010010" => rgb <= "000000";
					when "11010100011010011" => rgb <= "000000";
					when "11010100011010100" => rgb <= "000000";
					when "11010100011010101" => rgb <= "000000";
					when "11010100011010110" => rgb <= "000000";
					when "11010100011010111" => rgb <= "101010";
					when "11010100011011000" => rgb <= "111111";
					when "11010100011011001" => rgb <= "111111";
					when "11010100011011010" => rgb <= "101010";
					when "11010100011011011" => rgb <= "111111";
					when "11010100011011100" => rgb <= "111111";
					when "11010100011011101" => rgb <= "111111";
					when "11010100011011110" => rgb <= "111111";
					when "11010100011011111" => rgb <= "111111";
					when "11010100011100000" => rgb <= "111111";
					when "11010100011100001" => rgb <= "101010";
					when "11010100011100010" => rgb <= "101010";
					when "11010100011100011" => rgb <= "111111";
					when "11010100011100100" => rgb <= "111111";
					when "11010100011100101" => rgb <= "101010";
					when "11010100011100110" => rgb <= "000000";
					when "11010100011100111" => rgb <= "000000";
					when "11010100011101000" => rgb <= "000000";
					when "11010100011101001" => rgb <= "000000";
					when "11010100011101010" => rgb <= "000000";
					when "11010100011101011" => rgb <= "000000";
					when "11010100011101100" => rgb <= "000000";
					when "11010100011101101" => rgb <= "010101";
					when "11010100011101110" => rgb <= "111111";
					when "11010100011101111" => rgb <= "111111";
					when "11010100011110000" => rgb <= "111111";
					when "11010100011110001" => rgb <= "101010";
					when "11010100011110010" => rgb <= "111111";
					when "11010100011110011" => rgb <= "101010";
					when "11010100011110100" => rgb <= "101010";
					when "11010100011110101" => rgb <= "000000";
					when "11010100011110110" => rgb <= "000000";
					when "11010100011110111" => rgb <= "000000";
					when "11010100011111000" => rgb <= "000000";
					when "11010100011111001" => rgb <= "000000";
					when "11010100011111010" => rgb <= "000000";
					when "11010100011111011" => rgb <= "000000";
					when "11010100011111100" => rgb <= "000000";
					when "11010100011111101" => rgb <= "000000";
					when "11010100011111110" => rgb <= "000000";
					when "11010100011111111" => rgb <= "000000";
					when "11010100100000000" => rgb <= "000000";
					when "11010100100000001" => rgb <= "000000";
					when "11010100100000010" => rgb <= "000000";
					when "11010100100000011" => rgb <= "000000";
					when "11010100100000100" => rgb <= "000000";
					when "11010100100000101" => rgb <= "000000";
					when "11010100100000110" => rgb <= "000000";
					when "11010100100000111" => rgb <= "000000";
					when "11010100100001000" => rgb <= "000000";
					when "11010100100001001" => rgb <= "000000";
					when "11010100100001010" => rgb <= "000000";
					when "11010100100001011" => rgb <= "010101";
					when "11010100100001100" => rgb <= "101010";
					when "11010100100001101" => rgb <= "111111";
					when "11010100100001110" => rgb <= "111111";
					when "11010100100001111" => rgb <= "111111";
					when "11010100100010000" => rgb <= "111111";
					when "11010100100010001" => rgb <= "111111";
					when "11010100100010010" => rgb <= "111111";
					when "11010100100010011" => rgb <= "111111";
					when "11010100100010100" => rgb <= "111111";
					when "11010100100010101" => rgb <= "111111";
					when "11010100100010110" => rgb <= "111111";
					when "11010100100010111" => rgb <= "111111";
					when "11010100100011000" => rgb <= "111111";
					when "11010100100011001" => rgb <= "111111";
					when "11010100100011010" => rgb <= "101010";
					when "11010100100011011" => rgb <= "000000";
					when "11010100100011100" => rgb <= "000000";
					when "11010100100011101" => rgb <= "000000";
					when "11010100100011110" => rgb <= "000000";
					when "11010100100011111" => rgb <= "000000";
					when "11010100100100000" => rgb <= "000000";
					when "11010100100100001" => rgb <= "000000";
					when "11010100100100010" => rgb <= "101010";
					when "11010100100100011" => rgb <= "111111";
					when "11010100100100100" => rgb <= "111111";
					when "11010100100100101" => rgb <= "111111";
					when "11010100100100110" => rgb <= "111111";
					when "11010100100100111" => rgb <= "111111";
					when "11010100100101000" => rgb <= "111111";
					when "11010100100101001" => rgb <= "111111";
					when "11010100100101010" => rgb <= "111111";
					when "11010100100101011" => rgb <= "111111";
					when "11010100100101100" => rgb <= "111111";
					when "11010100100101101" => rgb <= "111111";
					when "11010100100101110" => rgb <= "111111";
					when "11010100100101111" => rgb <= "111111";
					when "11010100100110000" => rgb <= "101010";
					when "11010100100110001" => rgb <= "000000";
					when "11010100100110010" => rgb <= "000000";
					when "11010100100110011" => rgb <= "000000";
					when "11010100100110100" => rgb <= "000000";
					when "11010100100110101" => rgb <= "000000";
					when "11010100100110110" => rgb <= "000000";
					when "11010100100110111" => rgb <= "000000";
					when "11010100100111000" => rgb <= "000000";
					when "11010100100111001" => rgb <= "000000";
					when "11010100100111010" => rgb <= "000000";
					when "11010100100111011" => rgb <= "000000";
					when "11010100100111100" => rgb <= "000000";
					when "11010100100111101" => rgb <= "000000";
					when "11010100100111110" => rgb <= "000000";
					when "11010100100111111" => rgb <= "000000";
					when "11010101000000000" => rgb <= "000000";
					when "11010101000000001" => rgb <= "000000";
					when "11010101000000010" => rgb <= "000000";
					when "11010101000000011" => rgb <= "000000";
					when "11010101000000100" => rgb <= "000000";
					when "11010101000000101" => rgb <= "000000";
					when "11010101000000110" => rgb <= "000000";
					when "11010101000000111" => rgb <= "000000";
					when "11010101000001000" => rgb <= "000000";
					when "11010101000001001" => rgb <= "000000";
					when "11010101000001010" => rgb <= "000000";
					when "11010101000001011" => rgb <= "000000";
					when "11010101000001100" => rgb <= "000000";
					when "11010101000001101" => rgb <= "000000";
					when "11010101000001110" => rgb <= "000000";
					when "11010101000001111" => rgb <= "000000";
					when "11010101000010000" => rgb <= "000000";
					when "11010101000010001" => rgb <= "000000";
					when "11010101000010010" => rgb <= "000000";
					when "11010101000010011" => rgb <= "000000";
					when "11010101000010100" => rgb <= "010101";
					when "11010101000010101" => rgb <= "010101";
					when "11010101000010110" => rgb <= "010101";
					when "11010101000010111" => rgb <= "010101";
					when "11010101000011000" => rgb <= "010101";
					when "11010101000011001" => rgb <= "010101";
					when "11010101000011010" => rgb <= "010101";
					when "11010101000011011" => rgb <= "010101";
					when "11010101000011100" => rgb <= "010101";
					when "11010101000011101" => rgb <= "010101";
					when "11010101000011110" => rgb <= "010101";
					when "11010101000011111" => rgb <= "010101";
					when "11010101000100000" => rgb <= "010101";
					when "11010101000100001" => rgb <= "010101";
					when "11010101000100010" => rgb <= "010101";
					when "11010101000100011" => rgb <= "000000";
					when "11010101000100100" => rgb <= "000000";
					when "11010101000100101" => rgb <= "000000";
					when "11010101000100110" => rgb <= "000000";
					when "11010101000100111" => rgb <= "000000";
					when "11010101000101000" => rgb <= "000000";
					when "11010101000101001" => rgb <= "000000";
					when "11010101000101010" => rgb <= "000000";
					when "11010101000101011" => rgb <= "000000";
					when "11010101000101100" => rgb <= "000000";
					when "11010101000101101" => rgb <= "000000";
					when "11010101000101110" => rgb <= "000000";
					when "11010101000101111" => rgb <= "000000";
					when "11010101000110000" => rgb <= "000000";
					when "11010101000110001" => rgb <= "000000";
					when "11010101000110010" => rgb <= "000000";
					when "11010101000110011" => rgb <= "000000";
					when "11010101000110100" => rgb <= "000000";
					when "11010101000110101" => rgb <= "000000";
					when "11010101000110110" => rgb <= "000000";
					when "11010101000110111" => rgb <= "000000";
					when "11010101000111000" => rgb <= "000000";
					when "11010101000111001" => rgb <= "000000";
					when "11010101000111010" => rgb <= "000000";
					when "11010101000111011" => rgb <= "000000";
					when "11010101000111100" => rgb <= "000000";
					when "11010101000111101" => rgb <= "000000";
					when "11010101000111110" => rgb <= "000000";
					when "11010101000111111" => rgb <= "000000";
					when "11010101001000000" => rgb <= "000000";
					when "11010101001000001" => rgb <= "010101";
					when "11010101001000010" => rgb <= "010101";
					when "11010101001000011" => rgb <= "010101";
					when "11010101001000100" => rgb <= "010101";
					when "11010101001000101" => rgb <= "010101";
					when "11010101001000110" => rgb <= "010101";
					when "11010101001000111" => rgb <= "010101";
					when "11010101001001000" => rgb <= "010101";
					when "11010101001001001" => rgb <= "010101";
					when "11010101001001010" => rgb <= "010101";
					when "11010101001001011" => rgb <= "010101";
					when "11010101001001100" => rgb <= "010101";
					when "11010101001001101" => rgb <= "010101";
					when "11010101001001110" => rgb <= "010101";
					when "11010101001001111" => rgb <= "010101";
					when "11010101001010000" => rgb <= "010101";
					when "11010101001010001" => rgb <= "010101";
					when "11010101001010010" => rgb <= "010101";
					when "11010101001010011" => rgb <= "010101";
					when "11010101001010100" => rgb <= "010101";
					when "11010101001010101" => rgb <= "010101";
					when "11010101001010110" => rgb <= "010101";
					when "11010101001010111" => rgb <= "010101";
					when "11010101001011000" => rgb <= "000000";
					when "11010101001011001" => rgb <= "000000";
					when "11010101001011010" => rgb <= "000000";
					when "11010101001011011" => rgb <= "000000";
					when "11010101001011100" => rgb <= "000000";
					when "11010101001011101" => rgb <= "000000";
					when "11010101001011110" => rgb <= "000000";
					when "11010101001011111" => rgb <= "000000";
					when "11010101001100000" => rgb <= "000000";
					when "11010101001100001" => rgb <= "000000";
					when "11010101001100010" => rgb <= "000000";
					when "11010101001100011" => rgb <= "000000";
					when "11010101001100100" => rgb <= "000000";
					when "11010101001100101" => rgb <= "000000";
					when "11010101001100110" => rgb <= "000000";
					when "11010101001100111" => rgb <= "000000";
					when "11010101001101000" => rgb <= "000000";
					when "11010101001101001" => rgb <= "000000";
					when "11010101001101010" => rgb <= "000000";
					when "11010101001101011" => rgb <= "000000";
					when "11010101001101100" => rgb <= "000000";
					when "11010101001101101" => rgb <= "000000";
					when "11010101001101110" => rgb <= "010101";
					when "11010101001101111" => rgb <= "010101";
					when "11010101001110000" => rgb <= "010101";
					when "11010101001110001" => rgb <= "010101";
					when "11010101001110010" => rgb <= "010101";
					when "11010101001110011" => rgb <= "010101";
					when "11010101001110100" => rgb <= "010101";
					when "11010101001110101" => rgb <= "010101";
					when "11010101001110110" => rgb <= "010101";
					when "11010101001110111" => rgb <= "010101";
					when "11010101001111000" => rgb <= "010101";
					when "11010101001111001" => rgb <= "010101";
					when "11010101001111010" => rgb <= "010101";
					when "11010101001111011" => rgb <= "010101";
					when "11010101001111100" => rgb <= "010101";
					when "11010101001111101" => rgb <= "010101";
					when "11010101001111110" => rgb <= "010101";
					when "11010101001111111" => rgb <= "010101";
					when "11010101010000000" => rgb <= "010101";
					when "11010101010000001" => rgb <= "010101";
					when "11010101010000010" => rgb <= "010101";
					when "11010101010000011" => rgb <= "010101";
					when "11010101010000100" => rgb <= "010101";
					when "11010101010000101" => rgb <= "000000";
					when "11010101010000110" => rgb <= "000000";
					when "11010101010000111" => rgb <= "000000";
					when "11010101010001000" => rgb <= "000000";
					when "11010101010001001" => rgb <= "000000";
					when "11010101010001010" => rgb <= "000000";
					when "11010101010001011" => rgb <= "000000";
					when "11010101010001100" => rgb <= "000000";
					when "11010101010001101" => rgb <= "000000";
					when "11010101010001110" => rgb <= "000000";
					when "11010101010001111" => rgb <= "000000";
					when "11010101010010000" => rgb <= "000000";
					when "11010101010010001" => rgb <= "000000";
					when "11010101010010010" => rgb <= "000000";
					when "11010101010010011" => rgb <= "000000";
					when "11010101010010100" => rgb <= "000000";
					when "11010101010010101" => rgb <= "000000";
					when "11010101010010110" => rgb <= "000000";
					when "11010101010010111" => rgb <= "000000";
					when "11010101010011000" => rgb <= "000000";
					when "11010101010011001" => rgb <= "000000";
					when "11010101010011010" => rgb <= "000000";
					when "11010101010011011" => rgb <= "000000";
					when "11010101010011100" => rgb <= "000000";
					when "11010101010011101" => rgb <= "000000";
					when "11010101010011110" => rgb <= "000000";
					when "11010101010011111" => rgb <= "000000";
					when "11010101010100000" => rgb <= "000000";
					when "11010101010100001" => rgb <= "000000";
					when "11010101010100010" => rgb <= "000000";
					when "11010101010100011" => rgb <= "000000";
					when "11010101010100100" => rgb <= "000000";
					when "11010101010100101" => rgb <= "000000";
					when "11010101010100110" => rgb <= "000000";
					when "11010101010100111" => rgb <= "000000";
					when "11010101010101000" => rgb <= "000000";
					when "11010101010101001" => rgb <= "000000";
					when "11010101010101010" => rgb <= "010101";
					when "11010101010101011" => rgb <= "010101";
					when "11010101010101100" => rgb <= "010101";
					when "11010101010101101" => rgb <= "010101";
					when "11010101010101110" => rgb <= "010101";
					when "11010101010101111" => rgb <= "010101";
					when "11010101010110000" => rgb <= "010101";
					when "11010101010110001" => rgb <= "010101";
					when "11010101010110010" => rgb <= "000000";
					when "11010101010110011" => rgb <= "000000";
					when "11010101010110100" => rgb <= "000000";
					when "11010101010110101" => rgb <= "000000";
					when "11010101010110110" => rgb <= "000000";
					when "11010101010110111" => rgb <= "000000";
					when "11010101010111000" => rgb <= "000000";
					when "11010101010111001" => rgb <= "010101";
					when "11010101010111010" => rgb <= "010101";
					when "11010101010111011" => rgb <= "010101";
					when "11010101010111100" => rgb <= "010101";
					when "11010101010111101" => rgb <= "010101";
					when "11010101010111110" => rgb <= "010101";
					when "11010101010111111" => rgb <= "010101";
					when "11010101011000000" => rgb <= "010101";
					when "11010101011000001" => rgb <= "010101";
					when "11010101011000010" => rgb <= "010101";
					when "11010101011000011" => rgb <= "010101";
					when "11010101011000100" => rgb <= "010101";
					when "11010101011000101" => rgb <= "010101";
					when "11010101011000110" => rgb <= "010101";
					when "11010101011000111" => rgb <= "010101";
					when "11010101011001000" => rgb <= "000000";
					when "11010101011001001" => rgb <= "000000";
					when "11010101011001010" => rgb <= "000000";
					when "11010101011001011" => rgb <= "000000";
					when "11010101011001100" => rgb <= "000000";
					when "11010101011001101" => rgb <= "000000";
					when "11010101011001110" => rgb <= "000000";
					when "11010101011001111" => rgb <= "000000";
					when "11010101011010000" => rgb <= "000000";
					when "11010101011010001" => rgb <= "000000";
					when "11010101011010010" => rgb <= "000000";
					when "11010101011010011" => rgb <= "000000";
					when "11010101011010100" => rgb <= "000000";
					when "11010101011010101" => rgb <= "000000";
					when "11010101011010110" => rgb <= "000000";
					when "11010101011010111" => rgb <= "010101";
					when "11010101011011000" => rgb <= "010101";
					when "11010101011011001" => rgb <= "010101";
					when "11010101011011010" => rgb <= "010101";
					when "11010101011011011" => rgb <= "010101";
					when "11010101011011100" => rgb <= "010101";
					when "11010101011011101" => rgb <= "010101";
					when "11010101011011110" => rgb <= "010101";
					when "11010101011011111" => rgb <= "010101";
					when "11010101011100000" => rgb <= "010101";
					when "11010101011100001" => rgb <= "010101";
					when "11010101011100010" => rgb <= "010101";
					when "11010101011100011" => rgb <= "010101";
					when "11010101011100100" => rgb <= "010101";
					when "11010101011100101" => rgb <= "010101";
					when "11010101011100110" => rgb <= "000000";
					when "11010101011100111" => rgb <= "000000";
					when "11010101011101000" => rgb <= "000000";
					when "11010101011101001" => rgb <= "000000";
					when "11010101011101010" => rgb <= "000000";
					when "11010101011101011" => rgb <= "000000";
					when "11010101011101100" => rgb <= "000000";
					when "11010101011101101" => rgb <= "000000";
					when "11010101011101110" => rgb <= "010101";
					when "11010101011101111" => rgb <= "010101";
					when "11010101011110000" => rgb <= "010101";
					when "11010101011110001" => rgb <= "010101";
					when "11010101011110010" => rgb <= "010101";
					when "11010101011110011" => rgb <= "010101";
					when "11010101011110100" => rgb <= "010101";
					when "11010101011110101" => rgb <= "000000";
					when "11010101011110110" => rgb <= "000000";
					when "11010101011110111" => rgb <= "000000";
					when "11010101011111000" => rgb <= "000000";
					when "11010101011111001" => rgb <= "000000";
					when "11010101011111010" => rgb <= "000000";
					when "11010101011111011" => rgb <= "000000";
					when "11010101011111100" => rgb <= "000000";
					when "11010101011111101" => rgb <= "000000";
					when "11010101011111110" => rgb <= "000000";
					when "11010101011111111" => rgb <= "000000";
					when "11010101100000000" => rgb <= "000000";
					when "11010101100000001" => rgb <= "000000";
					when "11010101100000010" => rgb <= "000000";
					when "11010101100000011" => rgb <= "000000";
					when "11010101100000100" => rgb <= "000000";
					when "11010101100000101" => rgb <= "000000";
					when "11010101100000110" => rgb <= "000000";
					when "11010101100000111" => rgb <= "000000";
					when "11010101100001000" => rgb <= "000000";
					when "11010101100001001" => rgb <= "000000";
					when "11010101100001010" => rgb <= "000000";
					when "11010101100001011" => rgb <= "000000";
					when "11010101100001100" => rgb <= "010101";
					when "11010101100001101" => rgb <= "010101";
					when "11010101100001110" => rgb <= "010101";
					when "11010101100001111" => rgb <= "010101";
					when "11010101100010000" => rgb <= "010101";
					when "11010101100010001" => rgb <= "010101";
					when "11010101100010010" => rgb <= "010101";
					when "11010101100010011" => rgb <= "010101";
					when "11010101100010100" => rgb <= "010101";
					when "11010101100010101" => rgb <= "010101";
					when "11010101100010110" => rgb <= "010101";
					when "11010101100010111" => rgb <= "010101";
					when "11010101100011000" => rgb <= "010101";
					when "11010101100011001" => rgb <= "010101";
					when "11010101100011010" => rgb <= "010101";
					when "11010101100011011" => rgb <= "000000";
					when "11010101100011100" => rgb <= "000000";
					when "11010101100011101" => rgb <= "000000";
					when "11010101100011110" => rgb <= "000000";
					when "11010101100011111" => rgb <= "000000";
					when "11010101100100000" => rgb <= "000000";
					when "11010101100100001" => rgb <= "000000";
					when "11010101100100010" => rgb <= "010101";
					when "11010101100100011" => rgb <= "010101";
					when "11010101100100100" => rgb <= "010101";
					when "11010101100100101" => rgb <= "010101";
					when "11010101100100110" => rgb <= "010101";
					when "11010101100100111" => rgb <= "010101";
					when "11010101100101000" => rgb <= "010101";
					when "11010101100101001" => rgb <= "010101";
					when "11010101100101010" => rgb <= "010101";
					when "11010101100101011" => rgb <= "010101";
					when "11010101100101100" => rgb <= "010101";
					when "11010101100101101" => rgb <= "010101";
					when "11010101100101110" => rgb <= "010101";
					when "11010101100101111" => rgb <= "010101";
					when "11010101100110000" => rgb <= "010101";
					when "11010101100110001" => rgb <= "000000";
					when "11010101100110010" => rgb <= "000000";
					when "11010101100110011" => rgb <= "000000";
					when "11010101100110100" => rgb <= "000000";
					when "11010101100110101" => rgb <= "000000";
					when "11010101100110110" => rgb <= "000000";
					when "11010101100110111" => rgb <= "000000";
					when "11010101100111000" => rgb <= "000000";
					when "11010101100111001" => rgb <= "000000";
					when "11010101100111010" => rgb <= "000000";
					when "11010101100111011" => rgb <= "000000";
					when "11010101100111100" => rgb <= "000000";
					when "11010101100111101" => rgb <= "000000";
					when "11010101100111110" => rgb <= "000000";
					when "11010101100111111" => rgb <= "000000";
					when "11010110000000000" => rgb <= "000000";
					when "11010110000000001" => rgb <= "000000";
					when "11010110000000010" => rgb <= "000000";
					when "11010110000000011" => rgb <= "000000";
					when "11010110000000100" => rgb <= "000000";
					when "11010110000000101" => rgb <= "000000";
					when "11010110000000110" => rgb <= "000000";
					when "11010110000000111" => rgb <= "000000";
					when "11010110000001000" => rgb <= "000000";
					when "11010110000001001" => rgb <= "000000";
					when "11010110000001010" => rgb <= "000000";
					when "11010110000001011" => rgb <= "000000";
					when "11010110000001100" => rgb <= "000000";
					when "11010110000001101" => rgb <= "000000";
					when "11010110000001110" => rgb <= "000000";
					when "11010110000001111" => rgb <= "000000";
					when "11010110000010000" => rgb <= "000000";
					when "11010110000010001" => rgb <= "000000";
					when "11010110000010010" => rgb <= "000000";
					when "11010110000010011" => rgb <= "000000";
					when "11010110000010100" => rgb <= "000000";
					when "11010110000010101" => rgb <= "000000";
					when "11010110000010110" => rgb <= "000000";
					when "11010110000010111" => rgb <= "000000";
					when "11010110000011000" => rgb <= "000000";
					when "11010110000011001" => rgb <= "000000";
					when "11010110000011010" => rgb <= "000000";
					when "11010110000011011" => rgb <= "000000";
					when "11010110000011100" => rgb <= "000000";
					when "11010110000011101" => rgb <= "000000";
					when "11010110000011110" => rgb <= "000000";
					when "11010110000011111" => rgb <= "000000";
					when "11010110000100000" => rgb <= "000000";
					when "11010110000100001" => rgb <= "000000";
					when "11010110000100010" => rgb <= "000000";
					when "11010110000100011" => rgb <= "000000";
					when "11010110000100100" => rgb <= "000000";
					when "11010110000100101" => rgb <= "000000";
					when "11010110000100110" => rgb <= "000000";
					when "11010110000100111" => rgb <= "000000";
					when "11010110000101000" => rgb <= "000000";
					when "11010110000101001" => rgb <= "000000";
					when "11010110000101010" => rgb <= "000000";
					when "11010110000101011" => rgb <= "000000";
					when "11010110000101100" => rgb <= "000000";
					when "11010110000101101" => rgb <= "000000";
					when "11010110000101110" => rgb <= "000000";
					when "11010110000101111" => rgb <= "000000";
					when "11010110000110000" => rgb <= "000000";
					when "11010110000110001" => rgb <= "000000";
					when "11010110000110010" => rgb <= "000000";
					when "11010110000110011" => rgb <= "000000";
					when "11010110000110100" => rgb <= "000000";
					when "11010110000110101" => rgb <= "000000";
					when "11010110000110110" => rgb <= "000000";
					when "11010110000110111" => rgb <= "000000";
					when "11010110000111000" => rgb <= "000000";
					when "11010110000111001" => rgb <= "000000";
					when "11010110000111010" => rgb <= "000000";
					when "11010110000111011" => rgb <= "000000";
					when "11010110000111100" => rgb <= "000000";
					when "11010110000111101" => rgb <= "000000";
					when "11010110000111110" => rgb <= "000000";
					when "11010110000111111" => rgb <= "000000";
					when "11010110001000000" => rgb <= "000000";
					when "11010110001000001" => rgb <= "000000";
					when "11010110001000010" => rgb <= "000000";
					when "11010110001000011" => rgb <= "000000";
					when "11010110001000100" => rgb <= "000000";
					when "11010110001000101" => rgb <= "000000";
					when "11010110001000110" => rgb <= "000000";
					when "11010110001000111" => rgb <= "000000";
					when "11010110001001000" => rgb <= "000000";
					when "11010110001001001" => rgb <= "000000";
					when "11010110001001010" => rgb <= "000000";
					when "11010110001001011" => rgb <= "000000";
					when "11010110001001100" => rgb <= "000000";
					when "11010110001001101" => rgb <= "000000";
					when "11010110001001110" => rgb <= "000000";
					when "11010110001001111" => rgb <= "000000";
					when "11010110001010000" => rgb <= "000000";
					when "11010110001010001" => rgb <= "000000";
					when "11010110001010010" => rgb <= "000000";
					when "11010110001010011" => rgb <= "000000";
					when "11010110001010100" => rgb <= "000000";
					when "11010110001010101" => rgb <= "000000";
					when "11010110001010110" => rgb <= "000000";
					when "11010110001010111" => rgb <= "000000";
					when "11010110001011000" => rgb <= "000000";
					when "11010110001011001" => rgb <= "000000";
					when "11010110001011010" => rgb <= "000000";
					when "11010110001011011" => rgb <= "000000";
					when "11010110001011100" => rgb <= "000000";
					when "11010110001011101" => rgb <= "000000";
					when "11010110001011110" => rgb <= "000000";
					when "11010110001011111" => rgb <= "000000";
					when "11010110001100000" => rgb <= "000000";
					when "11010110001100001" => rgb <= "000000";
					when "11010110001100010" => rgb <= "000000";
					when "11010110001100011" => rgb <= "000000";
					when "11010110001100100" => rgb <= "000000";
					when "11010110001100101" => rgb <= "000000";
					when "11010110001100110" => rgb <= "000000";
					when "11010110001100111" => rgb <= "000000";
					when "11010110001101000" => rgb <= "000000";
					when "11010110001101001" => rgb <= "000000";
					when "11010110001101010" => rgb <= "000000";
					when "11010110001101011" => rgb <= "000000";
					when "11010110001101100" => rgb <= "000000";
					when "11010110001101101" => rgb <= "000000";
					when "11010110001101110" => rgb <= "000000";
					when "11010110001101111" => rgb <= "000000";
					when "11010110001110000" => rgb <= "000000";
					when "11010110001110001" => rgb <= "000000";
					when "11010110001110010" => rgb <= "000000";
					when "11010110001110011" => rgb <= "000000";
					when "11010110001110100" => rgb <= "000000";
					when "11010110001110101" => rgb <= "000000";
					when "11010110001110110" => rgb <= "000000";
					when "11010110001110111" => rgb <= "000000";
					when "11010110001111000" => rgb <= "000000";
					when "11010110001111001" => rgb <= "000000";
					when "11010110001111010" => rgb <= "000000";
					when "11010110001111011" => rgb <= "000000";
					when "11010110001111100" => rgb <= "000000";
					when "11010110001111101" => rgb <= "000000";
					when "11010110001111110" => rgb <= "000000";
					when "11010110001111111" => rgb <= "000000";
					when "11010110010000000" => rgb <= "000000";
					when "11010110010000001" => rgb <= "000000";
					when "11010110010000010" => rgb <= "000000";
					when "11010110010000011" => rgb <= "000000";
					when "11010110010000100" => rgb <= "000000";
					when "11010110010000101" => rgb <= "000000";
					when "11010110010000110" => rgb <= "000000";
					when "11010110010000111" => rgb <= "000000";
					when "11010110010001000" => rgb <= "000000";
					when "11010110010001001" => rgb <= "000000";
					when "11010110010001010" => rgb <= "000000";
					when "11010110010001011" => rgb <= "000000";
					when "11010110010001100" => rgb <= "000000";
					when "11010110010001101" => rgb <= "000000";
					when "11010110010001110" => rgb <= "000000";
					when "11010110010001111" => rgb <= "000000";
					when "11010110010010000" => rgb <= "000000";
					when "11010110010010001" => rgb <= "000000";
					when "11010110010010010" => rgb <= "000000";
					when "11010110010010011" => rgb <= "000000";
					when "11010110010010100" => rgb <= "000000";
					when "11010110010010101" => rgb <= "000000";
					when "11010110010010110" => rgb <= "000000";
					when "11010110010010111" => rgb <= "000000";
					when "11010110010011000" => rgb <= "000000";
					when "11010110010011001" => rgb <= "000000";
					when "11010110010011010" => rgb <= "000000";
					when "11010110010011011" => rgb <= "000000";
					when "11010110010011100" => rgb <= "000000";
					when "11010110010011101" => rgb <= "000000";
					when "11010110010011110" => rgb <= "000000";
					when "11010110010011111" => rgb <= "000000";
					when "11010110010100000" => rgb <= "000000";
					when "11010110010100001" => rgb <= "000000";
					when "11010110010100010" => rgb <= "000000";
					when "11010110010100011" => rgb <= "000000";
					when "11010110010100100" => rgb <= "000000";
					when "11010110010100101" => rgb <= "000000";
					when "11010110010100110" => rgb <= "000000";
					when "11010110010100111" => rgb <= "000000";
					when "11010110010101000" => rgb <= "000000";
					when "11010110010101001" => rgb <= "000000";
					when "11010110010101010" => rgb <= "000000";
					when "11010110010101011" => rgb <= "000000";
					when "11010110010101100" => rgb <= "000000";
					when "11010110010101101" => rgb <= "000000";
					when "11010110010101110" => rgb <= "000000";
					when "11010110010101111" => rgb <= "000000";
					when "11010110010110000" => rgb <= "000000";
					when "11010110010110001" => rgb <= "000000";
					when "11010110010110010" => rgb <= "000000";
					when "11010110010110011" => rgb <= "000000";
					when "11010110010110100" => rgb <= "000000";
					when "11010110010110101" => rgb <= "000000";
					when "11010110010110110" => rgb <= "000000";
					when "11010110010110111" => rgb <= "000000";
					when "11010110010111000" => rgb <= "000000";
					when "11010110010111001" => rgb <= "000000";
					when "11010110010111010" => rgb <= "000000";
					when "11010110010111011" => rgb <= "000000";
					when "11010110010111100" => rgb <= "000000";
					when "11010110010111101" => rgb <= "000000";
					when "11010110010111110" => rgb <= "000000";
					when "11010110010111111" => rgb <= "000000";
					when "11010110011000000" => rgb <= "000000";
					when "11010110011000001" => rgb <= "000000";
					when "11010110011000010" => rgb <= "000000";
					when "11010110011000011" => rgb <= "000000";
					when "11010110011000100" => rgb <= "000000";
					when "11010110011000101" => rgb <= "000000";
					when "11010110011000110" => rgb <= "000000";
					when "11010110011000111" => rgb <= "000000";
					when "11010110011001000" => rgb <= "000000";
					when "11010110011001001" => rgb <= "000000";
					when "11010110011001010" => rgb <= "000000";
					when "11010110011001011" => rgb <= "000000";
					when "11010110011001100" => rgb <= "000000";
					when "11010110011001101" => rgb <= "000000";
					when "11010110011001110" => rgb <= "000000";
					when "11010110011001111" => rgb <= "000000";
					when "11010110011010000" => rgb <= "000000";
					when "11010110011010001" => rgb <= "000000";
					when "11010110011010010" => rgb <= "000000";
					when "11010110011010011" => rgb <= "000000";
					when "11010110011010100" => rgb <= "000000";
					when "11010110011010101" => rgb <= "000000";
					when "11010110011010110" => rgb <= "000000";
					when "11010110011010111" => rgb <= "000000";
					when "11010110011011000" => rgb <= "000000";
					when "11010110011011001" => rgb <= "000000";
					when "11010110011011010" => rgb <= "000000";
					when "11010110011011011" => rgb <= "000000";
					when "11010110011011100" => rgb <= "000000";
					when "11010110011011101" => rgb <= "000000";
					when "11010110011011110" => rgb <= "000000";
					when "11010110011011111" => rgb <= "000000";
					when "11010110011100000" => rgb <= "000000";
					when "11010110011100001" => rgb <= "000000";
					when "11010110011100010" => rgb <= "000000";
					when "11010110011100011" => rgb <= "000000";
					when "11010110011100100" => rgb <= "000000";
					when "11010110011100101" => rgb <= "000000";
					when "11010110011100110" => rgb <= "000000";
					when "11010110011100111" => rgb <= "000000";
					when "11010110011101000" => rgb <= "000000";
					when "11010110011101001" => rgb <= "000000";
					when "11010110011101010" => rgb <= "000000";
					when "11010110011101011" => rgb <= "000000";
					when "11010110011101100" => rgb <= "000000";
					when "11010110011101101" => rgb <= "000000";
					when "11010110011101110" => rgb <= "000000";
					when "11010110011101111" => rgb <= "000000";
					when "11010110011110000" => rgb <= "000000";
					when "11010110011110001" => rgb <= "000000";
					when "11010110011110010" => rgb <= "000000";
					when "11010110011110011" => rgb <= "000000";
					when "11010110011110100" => rgb <= "000000";
					when "11010110011110101" => rgb <= "000000";
					when "11010110011110110" => rgb <= "000000";
					when "11010110011110111" => rgb <= "000000";
					when "11010110011111000" => rgb <= "000000";
					when "11010110011111001" => rgb <= "000000";
					when "11010110011111010" => rgb <= "000000";
					when "11010110011111011" => rgb <= "000000";
					when "11010110011111100" => rgb <= "000000";
					when "11010110011111101" => rgb <= "000000";
					when "11010110011111110" => rgb <= "000000";
					when "11010110011111111" => rgb <= "000000";
					when "11010110100000000" => rgb <= "000000";
					when "11010110100000001" => rgb <= "000000";
					when "11010110100000010" => rgb <= "000000";
					when "11010110100000011" => rgb <= "000000";
					when "11010110100000100" => rgb <= "000000";
					when "11010110100000101" => rgb <= "000000";
					when "11010110100000110" => rgb <= "000000";
					when "11010110100000111" => rgb <= "000000";
					when "11010110100001000" => rgb <= "000000";
					when "11010110100001001" => rgb <= "000000";
					when "11010110100001010" => rgb <= "000000";
					when "11010110100001011" => rgb <= "000000";
					when "11010110100001100" => rgb <= "000000";
					when "11010110100001101" => rgb <= "000000";
					when "11010110100001110" => rgb <= "000000";
					when "11010110100001111" => rgb <= "000000";
					when "11010110100010000" => rgb <= "000000";
					when "11010110100010001" => rgb <= "000000";
					when "11010110100010010" => rgb <= "000000";
					when "11010110100010011" => rgb <= "000000";
					when "11010110100010100" => rgb <= "000000";
					when "11010110100010101" => rgb <= "000000";
					when "11010110100010110" => rgb <= "000000";
					when "11010110100010111" => rgb <= "000000";
					when "11010110100011000" => rgb <= "000000";
					when "11010110100011001" => rgb <= "000000";
					when "11010110100011010" => rgb <= "000000";
					when "11010110100011011" => rgb <= "000000";
					when "11010110100011100" => rgb <= "000000";
					when "11010110100011101" => rgb <= "000000";
					when "11010110100011110" => rgb <= "000000";
					when "11010110100011111" => rgb <= "000000";
					when "11010110100100000" => rgb <= "000000";
					when "11010110100100001" => rgb <= "000000";
					when "11010110100100010" => rgb <= "000000";
					when "11010110100100011" => rgb <= "000000";
					when "11010110100100100" => rgb <= "000000";
					when "11010110100100101" => rgb <= "000000";
					when "11010110100100110" => rgb <= "000000";
					when "11010110100100111" => rgb <= "000000";
					when "11010110100101000" => rgb <= "000000";
					when "11010110100101001" => rgb <= "000000";
					when "11010110100101010" => rgb <= "000000";
					when "11010110100101011" => rgb <= "000000";
					when "11010110100101100" => rgb <= "000000";
					when "11010110100101101" => rgb <= "000000";
					when "11010110100101110" => rgb <= "000000";
					when "11010110100101111" => rgb <= "000000";
					when "11010110100110000" => rgb <= "000000";
					when "11010110100110001" => rgb <= "000000";
					when "11010110100110010" => rgb <= "000000";
					when "11010110100110011" => rgb <= "000000";
					when "11010110100110100" => rgb <= "000000";
					when "11010110100110101" => rgb <= "000000";
					when "11010110100110110" => rgb <= "000000";
					when "11010110100110111" => rgb <= "000000";
					when "11010110100111000" => rgb <= "000000";
					when "11010110100111001" => rgb <= "000000";
					when "11010110100111010" => rgb <= "000000";
					when "11010110100111011" => rgb <= "000000";
					when "11010110100111100" => rgb <= "000000";
					when "11010110100111101" => rgb <= "000000";
					when "11010110100111110" => rgb <= "000000";
					when "11010110100111111" => rgb <= "000000";
					when "11010111000000000" => rgb <= "000000";
					when "11010111000000001" => rgb <= "000000";
					when "11010111000000010" => rgb <= "000000";
					when "11010111000000011" => rgb <= "000000";
					when "11010111000000100" => rgb <= "000000";
					when "11010111000000101" => rgb <= "000000";
					when "11010111000000110" => rgb <= "000000";
					when "11010111000000111" => rgb <= "000000";
					when "11010111000001000" => rgb <= "000000";
					when "11010111000001001" => rgb <= "000000";
					when "11010111000001010" => rgb <= "000000";
					when "11010111000001011" => rgb <= "000000";
					when "11010111000001100" => rgb <= "000000";
					when "11010111000001101" => rgb <= "000000";
					when "11010111000001110" => rgb <= "000000";
					when "11010111000001111" => rgb <= "000000";
					when "11010111000010000" => rgb <= "000000";
					when "11010111000010001" => rgb <= "000000";
					when "11010111000010010" => rgb <= "000000";
					when "11010111000010011" => rgb <= "000000";
					when "11010111000010100" => rgb <= "000000";
					when "11010111000010101" => rgb <= "000000";
					when "11010111000010110" => rgb <= "000000";
					when "11010111000010111" => rgb <= "000000";
					when "11010111000011000" => rgb <= "000000";
					when "11010111000011001" => rgb <= "000000";
					when "11010111000011010" => rgb <= "000000";
					when "11010111000011011" => rgb <= "000000";
					when "11010111000011100" => rgb <= "000000";
					when "11010111000011101" => rgb <= "000000";
					when "11010111000011110" => rgb <= "000000";
					when "11010111000011111" => rgb <= "000000";
					when "11010111000100000" => rgb <= "000000";
					when "11010111000100001" => rgb <= "000000";
					when "11010111000100010" => rgb <= "000000";
					when "11010111000100011" => rgb <= "000000";
					when "11010111000100100" => rgb <= "000000";
					when "11010111000100101" => rgb <= "000000";
					when "11010111000100110" => rgb <= "000000";
					when "11010111000100111" => rgb <= "000000";
					when "11010111000101000" => rgb <= "000000";
					when "11010111000101001" => rgb <= "000000";
					when "11010111000101010" => rgb <= "000000";
					when "11010111000101011" => rgb <= "000000";
					when "11010111000101100" => rgb <= "000000";
					when "11010111000101101" => rgb <= "000000";
					when "11010111000101110" => rgb <= "000000";
					when "11010111000101111" => rgb <= "000000";
					when "11010111000110000" => rgb <= "000000";
					when "11010111000110001" => rgb <= "000000";
					when "11010111000110010" => rgb <= "000000";
					when "11010111000110011" => rgb <= "000000";
					when "11010111000110100" => rgb <= "000000";
					when "11010111000110101" => rgb <= "000000";
					when "11010111000110110" => rgb <= "000000";
					when "11010111000110111" => rgb <= "000000";
					when "11010111000111000" => rgb <= "000000";
					when "11010111000111001" => rgb <= "000000";
					when "11010111000111010" => rgb <= "000000";
					when "11010111000111011" => rgb <= "000000";
					when "11010111000111100" => rgb <= "000000";
					when "11010111000111101" => rgb <= "000000";
					when "11010111000111110" => rgb <= "000000";
					when "11010111000111111" => rgb <= "000000";
					when "11010111001000000" => rgb <= "000000";
					when "11010111001000001" => rgb <= "000000";
					when "11010111001000010" => rgb <= "000000";
					when "11010111001000011" => rgb <= "000000";
					when "11010111001000100" => rgb <= "000000";
					when "11010111001000101" => rgb <= "000000";
					when "11010111001000110" => rgb <= "000000";
					when "11010111001000111" => rgb <= "000000";
					when "11010111001001000" => rgb <= "000000";
					when "11010111001001001" => rgb <= "000000";
					when "11010111001001010" => rgb <= "000000";
					when "11010111001001011" => rgb <= "000000";
					when "11010111001001100" => rgb <= "000000";
					when "11010111001001101" => rgb <= "000000";
					when "11010111001001110" => rgb <= "000000";
					when "11010111001001111" => rgb <= "000000";
					when "11010111001010000" => rgb <= "000000";
					when "11010111001010001" => rgb <= "000000";
					when "11010111001010010" => rgb <= "000000";
					when "11010111001010011" => rgb <= "000000";
					when "11010111001010100" => rgb <= "000000";
					when "11010111001010101" => rgb <= "000000";
					when "11010111001010110" => rgb <= "000000";
					when "11010111001010111" => rgb <= "000000";
					when "11010111001011000" => rgb <= "000000";
					when "11010111001011001" => rgb <= "000000";
					when "11010111001011010" => rgb <= "000000";
					when "11010111001011011" => rgb <= "000000";
					when "11010111001011100" => rgb <= "000000";
					when "11010111001011101" => rgb <= "000000";
					when "11010111001011110" => rgb <= "000000";
					when "11010111001011111" => rgb <= "000000";
					when "11010111001100000" => rgb <= "000000";
					when "11010111001100001" => rgb <= "000000";
					when "11010111001100010" => rgb <= "000000";
					when "11010111001100011" => rgb <= "000000";
					when "11010111001100100" => rgb <= "000000";
					when "11010111001100101" => rgb <= "000000";
					when "11010111001100110" => rgb <= "000000";
					when "11010111001100111" => rgb <= "000000";
					when "11010111001101000" => rgb <= "000000";
					when "11010111001101001" => rgb <= "000000";
					when "11010111001101010" => rgb <= "000000";
					when "11010111001101011" => rgb <= "000000";
					when "11010111001101100" => rgb <= "000000";
					when "11010111001101101" => rgb <= "000000";
					when "11010111001101110" => rgb <= "000000";
					when "11010111001101111" => rgb <= "000000";
					when "11010111001110000" => rgb <= "000000";
					when "11010111001110001" => rgb <= "000000";
					when "11010111001110010" => rgb <= "000000";
					when "11010111001110011" => rgb <= "000000";
					when "11010111001110100" => rgb <= "000000";
					when "11010111001110101" => rgb <= "000000";
					when "11010111001110110" => rgb <= "000000";
					when "11010111001110111" => rgb <= "000000";
					when "11010111001111000" => rgb <= "000000";
					when "11010111001111001" => rgb <= "000000";
					when "11010111001111010" => rgb <= "000000";
					when "11010111001111011" => rgb <= "000000";
					when "11010111001111100" => rgb <= "000000";
					when "11010111001111101" => rgb <= "000000";
					when "11010111001111110" => rgb <= "000000";
					when "11010111001111111" => rgb <= "000000";
					when "11010111010000000" => rgb <= "000000";
					when "11010111010000001" => rgb <= "000000";
					when "11010111010000010" => rgb <= "000000";
					when "11010111010000011" => rgb <= "000000";
					when "11010111010000100" => rgb <= "000000";
					when "11010111010000101" => rgb <= "000000";
					when "11010111010000110" => rgb <= "000000";
					when "11010111010000111" => rgb <= "000000";
					when "11010111010001000" => rgb <= "000000";
					when "11010111010001001" => rgb <= "000000";
					when "11010111010001010" => rgb <= "000000";
					when "11010111010001011" => rgb <= "000000";
					when "11010111010001100" => rgb <= "000000";
					when "11010111010001101" => rgb <= "000000";
					when "11010111010001110" => rgb <= "000000";
					when "11010111010001111" => rgb <= "000000";
					when "11010111010010000" => rgb <= "000000";
					when "11010111010010001" => rgb <= "000000";
					when "11010111010010010" => rgb <= "000000";
					when "11010111010010011" => rgb <= "000000";
					when "11010111010010100" => rgb <= "000000";
					when "11010111010010101" => rgb <= "000000";
					when "11010111010010110" => rgb <= "000000";
					when "11010111010010111" => rgb <= "000000";
					when "11010111010011000" => rgb <= "000000";
					when "11010111010011001" => rgb <= "000000";
					when "11010111010011010" => rgb <= "000000";
					when "11010111010011011" => rgb <= "000000";
					when "11010111010011100" => rgb <= "000000";
					when "11010111010011101" => rgb <= "000000";
					when "11010111010011110" => rgb <= "000000";
					when "11010111010011111" => rgb <= "000000";
					when "11010111010100000" => rgb <= "000000";
					when "11010111010100001" => rgb <= "000000";
					when "11010111010100010" => rgb <= "000000";
					when "11010111010100011" => rgb <= "000000";
					when "11010111010100100" => rgb <= "000000";
					when "11010111010100101" => rgb <= "000000";
					when "11010111010100110" => rgb <= "000000";
					when "11010111010100111" => rgb <= "000000";
					when "11010111010101000" => rgb <= "000000";
					when "11010111010101001" => rgb <= "000000";
					when "11010111010101010" => rgb <= "000000";
					when "11010111010101011" => rgb <= "000000";
					when "11010111010101100" => rgb <= "000000";
					when "11010111010101101" => rgb <= "000000";
					when "11010111010101110" => rgb <= "000000";
					when "11010111010101111" => rgb <= "000000";
					when "11010111010110000" => rgb <= "000000";
					when "11010111010110001" => rgb <= "000000";
					when "11010111010110010" => rgb <= "000000";
					when "11010111010110011" => rgb <= "000000";
					when "11010111010110100" => rgb <= "000000";
					when "11010111010110101" => rgb <= "000000";
					when "11010111010110110" => rgb <= "000000";
					when "11010111010110111" => rgb <= "000000";
					when "11010111010111000" => rgb <= "000000";
					when "11010111010111001" => rgb <= "000000";
					when "11010111010111010" => rgb <= "000000";
					when "11010111010111011" => rgb <= "000000";
					when "11010111010111100" => rgb <= "000000";
					when "11010111010111101" => rgb <= "000000";
					when "11010111010111110" => rgb <= "000000";
					when "11010111010111111" => rgb <= "000000";
					when "11010111011000000" => rgb <= "000000";
					when "11010111011000001" => rgb <= "000000";
					when "11010111011000010" => rgb <= "000000";
					when "11010111011000011" => rgb <= "000000";
					when "11010111011000100" => rgb <= "000000";
					when "11010111011000101" => rgb <= "000000";
					when "11010111011000110" => rgb <= "000000";
					when "11010111011000111" => rgb <= "000000";
					when "11010111011001000" => rgb <= "000000";
					when "11010111011001001" => rgb <= "000000";
					when "11010111011001010" => rgb <= "000000";
					when "11010111011001011" => rgb <= "000000";
					when "11010111011001100" => rgb <= "000000";
					when "11010111011001101" => rgb <= "000000";
					when "11010111011001110" => rgb <= "000000";
					when "11010111011001111" => rgb <= "000000";
					when "11010111011010000" => rgb <= "000000";
					when "11010111011010001" => rgb <= "000000";
					when "11010111011010010" => rgb <= "000000";
					when "11010111011010011" => rgb <= "000000";
					when "11010111011010100" => rgb <= "000000";
					when "11010111011010101" => rgb <= "000000";
					when "11010111011010110" => rgb <= "000000";
					when "11010111011010111" => rgb <= "000000";
					when "11010111011011000" => rgb <= "000000";
					when "11010111011011001" => rgb <= "000000";
					when "11010111011011010" => rgb <= "000000";
					when "11010111011011011" => rgb <= "000000";
					when "11010111011011100" => rgb <= "000000";
					when "11010111011011101" => rgb <= "000000";
					when "11010111011011110" => rgb <= "000000";
					when "11010111011011111" => rgb <= "000000";
					when "11010111011100000" => rgb <= "000000";
					when "11010111011100001" => rgb <= "000000";
					when "11010111011100010" => rgb <= "000000";
					when "11010111011100011" => rgb <= "000000";
					when "11010111011100100" => rgb <= "000000";
					when "11010111011100101" => rgb <= "000000";
					when "11010111011100110" => rgb <= "000000";
					when "11010111011100111" => rgb <= "000000";
					when "11010111011101000" => rgb <= "000000";
					when "11010111011101001" => rgb <= "000000";
					when "11010111011101010" => rgb <= "000000";
					when "11010111011101011" => rgb <= "000000";
					when "11010111011101100" => rgb <= "000000";
					when "11010111011101101" => rgb <= "000000";
					when "11010111011101110" => rgb <= "000000";
					when "11010111011101111" => rgb <= "000000";
					when "11010111011110000" => rgb <= "000000";
					when "11010111011110001" => rgb <= "000000";
					when "11010111011110010" => rgb <= "000000";
					when "11010111011110011" => rgb <= "000000";
					when "11010111011110100" => rgb <= "000000";
					when "11010111011110101" => rgb <= "000000";
					when "11010111011110110" => rgb <= "000000";
					when "11010111011110111" => rgb <= "000000";
					when "11010111011111000" => rgb <= "000000";
					when "11010111011111001" => rgb <= "000000";
					when "11010111011111010" => rgb <= "000000";
					when "11010111011111011" => rgb <= "000000";
					when "11010111011111100" => rgb <= "000000";
					when "11010111011111101" => rgb <= "000000";
					when "11010111011111110" => rgb <= "000000";
					when "11010111011111111" => rgb <= "000000";
					when "11010111100000000" => rgb <= "000000";
					when "11010111100000001" => rgb <= "000000";
					when "11010111100000010" => rgb <= "000000";
					when "11010111100000011" => rgb <= "000000";
					when "11010111100000100" => rgb <= "000000";
					when "11010111100000101" => rgb <= "000000";
					when "11010111100000110" => rgb <= "000000";
					when "11010111100000111" => rgb <= "000000";
					when "11010111100001000" => rgb <= "000000";
					when "11010111100001001" => rgb <= "000000";
					when "11010111100001010" => rgb <= "000000";
					when "11010111100001011" => rgb <= "000000";
					when "11010111100001100" => rgb <= "000000";
					when "11010111100001101" => rgb <= "000000";
					when "11010111100001110" => rgb <= "000000";
					when "11010111100001111" => rgb <= "000000";
					when "11010111100010000" => rgb <= "000000";
					when "11010111100010001" => rgb <= "000000";
					when "11010111100010010" => rgb <= "000000";
					when "11010111100010011" => rgb <= "000000";
					when "11010111100010100" => rgb <= "000000";
					when "11010111100010101" => rgb <= "000000";
					when "11010111100010110" => rgb <= "000000";
					when "11010111100010111" => rgb <= "000000";
					when "11010111100011000" => rgb <= "000000";
					when "11010111100011001" => rgb <= "000000";
					when "11010111100011010" => rgb <= "000000";
					when "11010111100011011" => rgb <= "000000";
					when "11010111100011100" => rgb <= "000000";
					when "11010111100011101" => rgb <= "000000";
					when "11010111100011110" => rgb <= "000000";
					when "11010111100011111" => rgb <= "000000";
					when "11010111100100000" => rgb <= "000000";
					when "11010111100100001" => rgb <= "000000";
					when "11010111100100010" => rgb <= "000000";
					when "11010111100100011" => rgb <= "000000";
					when "11010111100100100" => rgb <= "000000";
					when "11010111100100101" => rgb <= "000000";
					when "11010111100100110" => rgb <= "000000";
					when "11010111100100111" => rgb <= "000000";
					when "11010111100101000" => rgb <= "000000";
					when "11010111100101001" => rgb <= "000000";
					when "11010111100101010" => rgb <= "000000";
					when "11010111100101011" => rgb <= "000000";
					when "11010111100101100" => rgb <= "000000";
					when "11010111100101101" => rgb <= "000000";
					when "11010111100101110" => rgb <= "000000";
					when "11010111100101111" => rgb <= "000000";
					when "11010111100110000" => rgb <= "000000";
					when "11010111100110001" => rgb <= "000000";
					when "11010111100110010" => rgb <= "000000";
					when "11010111100110011" => rgb <= "000000";
					when "11010111100110100" => rgb <= "000000";
					when "11010111100110101" => rgb <= "000000";
					when "11010111100110110" => rgb <= "000000";
					when "11010111100110111" => rgb <= "000000";
					when "11010111100111000" => rgb <= "000000";
					when "11010111100111001" => rgb <= "000000";
					when "11010111100111010" => rgb <= "000000";
					when "11010111100111011" => rgb <= "000000";
					when "11010111100111100" => rgb <= "000000";
					when "11010111100111101" => rgb <= "000000";
					when "11010111100111110" => rgb <= "000000";
					when "11010111100111111" => rgb <= "000000";
					when "11011000000000000" => rgb <= "000000";
					when "11011000000000001" => rgb <= "000000";
					when "11011000000000010" => rgb <= "000000";
					when "11011000000000011" => rgb <= "000000";
					when "11011000000000100" => rgb <= "000000";
					when "11011000000000101" => rgb <= "000000";
					when "11011000000000110" => rgb <= "000000";
					when "11011000000000111" => rgb <= "000000";
					when "11011000000001000" => rgb <= "000000";
					when "11011000000001001" => rgb <= "000000";
					when "11011000000001010" => rgb <= "000000";
					when "11011000000001011" => rgb <= "000000";
					when "11011000000001100" => rgb <= "000000";
					when "11011000000001101" => rgb <= "000000";
					when "11011000000001110" => rgb <= "000000";
					when "11011000000001111" => rgb <= "000000";
					when "11011000000010000" => rgb <= "000000";
					when "11011000000010001" => rgb <= "000000";
					when "11011000000010010" => rgb <= "000000";
					when "11011000000010011" => rgb <= "000000";
					when "11011000000010100" => rgb <= "000000";
					when "11011000000010101" => rgb <= "000000";
					when "11011000000010110" => rgb <= "000000";
					when "11011000000010111" => rgb <= "000000";
					when "11011000000011000" => rgb <= "000000";
					when "11011000000011001" => rgb <= "000000";
					when "11011000000011010" => rgb <= "000000";
					when "11011000000011011" => rgb <= "000000";
					when "11011000000011100" => rgb <= "000000";
					when "11011000000011101" => rgb <= "000000";
					when "11011000000011110" => rgb <= "000000";
					when "11011000000011111" => rgb <= "000000";
					when "11011000000100000" => rgb <= "000000";
					when "11011000000100001" => rgb <= "000000";
					when "11011000000100010" => rgb <= "000000";
					when "11011000000100011" => rgb <= "000000";
					when "11011000000100100" => rgb <= "000000";
					when "11011000000100101" => rgb <= "000000";
					when "11011000000100110" => rgb <= "000000";
					when "11011000000100111" => rgb <= "000000";
					when "11011000000101000" => rgb <= "000000";
					when "11011000000101001" => rgb <= "000000";
					when "11011000000101010" => rgb <= "000000";
					when "11011000000101011" => rgb <= "000000";
					when "11011000000101100" => rgb <= "000000";
					when "11011000000101101" => rgb <= "000000";
					when "11011000000101110" => rgb <= "000000";
					when "11011000000101111" => rgb <= "000000";
					when "11011000000110000" => rgb <= "000000";
					when "11011000000110001" => rgb <= "000000";
					when "11011000000110010" => rgb <= "000000";
					when "11011000000110011" => rgb <= "000000";
					when "11011000000110100" => rgb <= "000000";
					when "11011000000110101" => rgb <= "000000";
					when "11011000000110110" => rgb <= "000000";
					when "11011000000110111" => rgb <= "000000";
					when "11011000000111000" => rgb <= "000000";
					when "11011000000111001" => rgb <= "000000";
					when "11011000000111010" => rgb <= "000000";
					when "11011000000111011" => rgb <= "000000";
					when "11011000000111100" => rgb <= "000000";
					when "11011000000111101" => rgb <= "000000";
					when "11011000000111110" => rgb <= "000000";
					when "11011000000111111" => rgb <= "000000";
					when "11011000001000000" => rgb <= "000000";
					when "11011000001000001" => rgb <= "000000";
					when "11011000001000010" => rgb <= "000000";
					when "11011000001000011" => rgb <= "000000";
					when "11011000001000100" => rgb <= "000000";
					when "11011000001000101" => rgb <= "000000";
					when "11011000001000110" => rgb <= "000000";
					when "11011000001000111" => rgb <= "000000";
					when "11011000001001000" => rgb <= "000000";
					when "11011000001001001" => rgb <= "000000";
					when "11011000001001010" => rgb <= "000000";
					when "11011000001001011" => rgb <= "000000";
					when "11011000001001100" => rgb <= "000000";
					when "11011000001001101" => rgb <= "000000";
					when "11011000001001110" => rgb <= "000000";
					when "11011000001001111" => rgb <= "000000";
					when "11011000001010000" => rgb <= "000000";
					when "11011000001010001" => rgb <= "000000";
					when "11011000001010010" => rgb <= "000000";
					when "11011000001010011" => rgb <= "000000";
					when "11011000001010100" => rgb <= "000000";
					when "11011000001010101" => rgb <= "000000";
					when "11011000001010110" => rgb <= "000000";
					when "11011000001010111" => rgb <= "000000";
					when "11011000001011000" => rgb <= "000000";
					when "11011000001011001" => rgb <= "000000";
					when "11011000001011010" => rgb <= "000000";
					when "11011000001011011" => rgb <= "000000";
					when "11011000001011100" => rgb <= "000000";
					when "11011000001011101" => rgb <= "000000";
					when "11011000001011110" => rgb <= "000000";
					when "11011000001011111" => rgb <= "000000";
					when "11011000001100000" => rgb <= "000000";
					when "11011000001100001" => rgb <= "000000";
					when "11011000001100010" => rgb <= "000000";
					when "11011000001100011" => rgb <= "000000";
					when "11011000001100100" => rgb <= "000000";
					when "11011000001100101" => rgb <= "000000";
					when "11011000001100110" => rgb <= "000000";
					when "11011000001100111" => rgb <= "000000";
					when "11011000001101000" => rgb <= "000000";
					when "11011000001101001" => rgb <= "000000";
					when "11011000001101010" => rgb <= "000000";
					when "11011000001101011" => rgb <= "000000";
					when "11011000001101100" => rgb <= "000000";
					when "11011000001101101" => rgb <= "000000";
					when "11011000001101110" => rgb <= "000000";
					when "11011000001101111" => rgb <= "000000";
					when "11011000001110000" => rgb <= "000000";
					when "11011000001110001" => rgb <= "000000";
					when "11011000001110010" => rgb <= "000000";
					when "11011000001110011" => rgb <= "000000";
					when "11011000001110100" => rgb <= "000000";
					when "11011000001110101" => rgb <= "000000";
					when "11011000001110110" => rgb <= "000000";
					when "11011000001110111" => rgb <= "000000";
					when "11011000001111000" => rgb <= "000000";
					when "11011000001111001" => rgb <= "000000";
					when "11011000001111010" => rgb <= "000000";
					when "11011000001111011" => rgb <= "000000";
					when "11011000001111100" => rgb <= "000000";
					when "11011000001111101" => rgb <= "000000";
					when "11011000001111110" => rgb <= "000000";
					when "11011000001111111" => rgb <= "000000";
					when "11011000010000000" => rgb <= "000000";
					when "11011000010000001" => rgb <= "000000";
					when "11011000010000010" => rgb <= "000000";
					when "11011000010000011" => rgb <= "000000";
					when "11011000010000100" => rgb <= "000000";
					when "11011000010000101" => rgb <= "000000";
					when "11011000010000110" => rgb <= "000000";
					when "11011000010000111" => rgb <= "000000";
					when "11011000010001000" => rgb <= "000000";
					when "11011000010001001" => rgb <= "000000";
					when "11011000010001010" => rgb <= "000000";
					when "11011000010001011" => rgb <= "000000";
					when "11011000010001100" => rgb <= "000000";
					when "11011000010001101" => rgb <= "000000";
					when "11011000010001110" => rgb <= "000000";
					when "11011000010001111" => rgb <= "000000";
					when "11011000010010000" => rgb <= "000000";
					when "11011000010010001" => rgb <= "000000";
					when "11011000010010010" => rgb <= "000000";
					when "11011000010010011" => rgb <= "000000";
					when "11011000010010100" => rgb <= "000000";
					when "11011000010010101" => rgb <= "000000";
					when "11011000010010110" => rgb <= "000000";
					when "11011000010010111" => rgb <= "000000";
					when "11011000010011000" => rgb <= "000000";
					when "11011000010011001" => rgb <= "000000";
					when "11011000010011010" => rgb <= "000000";
					when "11011000010011011" => rgb <= "000000";
					when "11011000010011100" => rgb <= "000000";
					when "11011000010011101" => rgb <= "000000";
					when "11011000010011110" => rgb <= "000000";
					when "11011000010011111" => rgb <= "000000";
					when "11011000010100000" => rgb <= "000000";
					when "11011000010100001" => rgb <= "000000";
					when "11011000010100010" => rgb <= "000000";
					when "11011000010100011" => rgb <= "000000";
					when "11011000010100100" => rgb <= "000000";
					when "11011000010100101" => rgb <= "000000";
					when "11011000010100110" => rgb <= "000000";
					when "11011000010100111" => rgb <= "000000";
					when "11011000010101000" => rgb <= "000000";
					when "11011000010101001" => rgb <= "000000";
					when "11011000010101010" => rgb <= "000000";
					when "11011000010101011" => rgb <= "000000";
					when "11011000010101100" => rgb <= "000000";
					when "11011000010101101" => rgb <= "000000";
					when "11011000010101110" => rgb <= "000000";
					when "11011000010101111" => rgb <= "000000";
					when "11011000010110000" => rgb <= "000000";
					when "11011000010110001" => rgb <= "000000";
					when "11011000010110010" => rgb <= "000000";
					when "11011000010110011" => rgb <= "000000";
					when "11011000010110100" => rgb <= "000000";
					when "11011000010110101" => rgb <= "000000";
					when "11011000010110110" => rgb <= "000000";
					when "11011000010110111" => rgb <= "000000";
					when "11011000010111000" => rgb <= "000000";
					when "11011000010111001" => rgb <= "000000";
					when "11011000010111010" => rgb <= "000000";
					when "11011000010111011" => rgb <= "000000";
					when "11011000010111100" => rgb <= "000000";
					when "11011000010111101" => rgb <= "000000";
					when "11011000010111110" => rgb <= "000000";
					when "11011000010111111" => rgb <= "000000";
					when "11011000011000000" => rgb <= "000000";
					when "11011000011000001" => rgb <= "000000";
					when "11011000011000010" => rgb <= "000000";
					when "11011000011000011" => rgb <= "000000";
					when "11011000011000100" => rgb <= "000000";
					when "11011000011000101" => rgb <= "000000";
					when "11011000011000110" => rgb <= "000000";
					when "11011000011000111" => rgb <= "000000";
					when "11011000011001000" => rgb <= "000000";
					when "11011000011001001" => rgb <= "000000";
					when "11011000011001010" => rgb <= "000000";
					when "11011000011001011" => rgb <= "000000";
					when "11011000011001100" => rgb <= "000000";
					when "11011000011001101" => rgb <= "000000";
					when "11011000011001110" => rgb <= "000000";
					when "11011000011001111" => rgb <= "000000";
					when "11011000011010000" => rgb <= "000000";
					when "11011000011010001" => rgb <= "000000";
					when "11011000011010010" => rgb <= "000000";
					when "11011000011010011" => rgb <= "000000";
					when "11011000011010100" => rgb <= "000000";
					when "11011000011010101" => rgb <= "000000";
					when "11011000011010110" => rgb <= "000000";
					when "11011000011010111" => rgb <= "000000";
					when "11011000011011000" => rgb <= "000000";
					when "11011000011011001" => rgb <= "000000";
					when "11011000011011010" => rgb <= "000000";
					when "11011000011011011" => rgb <= "000000";
					when "11011000011011100" => rgb <= "000000";
					when "11011000011011101" => rgb <= "000000";
					when "11011000011011110" => rgb <= "000000";
					when "11011000011011111" => rgb <= "000000";
					when "11011000011100000" => rgb <= "000000";
					when "11011000011100001" => rgb <= "000000";
					when "11011000011100010" => rgb <= "000000";
					when "11011000011100011" => rgb <= "000000";
					when "11011000011100100" => rgb <= "000000";
					when "11011000011100101" => rgb <= "000000";
					when "11011000011100110" => rgb <= "000000";
					when "11011000011100111" => rgb <= "000000";
					when "11011000011101000" => rgb <= "000000";
					when "11011000011101001" => rgb <= "000000";
					when "11011000011101010" => rgb <= "000000";
					when "11011000011101011" => rgb <= "000000";
					when "11011000011101100" => rgb <= "000000";
					when "11011000011101101" => rgb <= "000000";
					when "11011000011101110" => rgb <= "000000";
					when "11011000011101111" => rgb <= "000000";
					when "11011000011110000" => rgb <= "000000";
					when "11011000011110001" => rgb <= "000000";
					when "11011000011110010" => rgb <= "000000";
					when "11011000011110011" => rgb <= "000000";
					when "11011000011110100" => rgb <= "000000";
					when "11011000011110101" => rgb <= "000000";
					when "11011000011110110" => rgb <= "000000";
					when "11011000011110111" => rgb <= "000000";
					when "11011000011111000" => rgb <= "000000";
					when "11011000011111001" => rgb <= "000000";
					when "11011000011111010" => rgb <= "000000";
					when "11011000011111011" => rgb <= "000000";
					when "11011000011111100" => rgb <= "000000";
					when "11011000011111101" => rgb <= "000000";
					when "11011000011111110" => rgb <= "000000";
					when "11011000011111111" => rgb <= "000000";
					when "11011000100000000" => rgb <= "000000";
					when "11011000100000001" => rgb <= "000000";
					when "11011000100000010" => rgb <= "000000";
					when "11011000100000011" => rgb <= "000000";
					when "11011000100000100" => rgb <= "000000";
					when "11011000100000101" => rgb <= "000000";
					when "11011000100000110" => rgb <= "000000";
					when "11011000100000111" => rgb <= "000000";
					when "11011000100001000" => rgb <= "000000";
					when "11011000100001001" => rgb <= "000000";
					when "11011000100001010" => rgb <= "000000";
					when "11011000100001011" => rgb <= "000000";
					when "11011000100001100" => rgb <= "000000";
					when "11011000100001101" => rgb <= "000000";
					when "11011000100001110" => rgb <= "000000";
					when "11011000100001111" => rgb <= "000000";
					when "11011000100010000" => rgb <= "000000";
					when "11011000100010001" => rgb <= "000000";
					when "11011000100010010" => rgb <= "000000";
					when "11011000100010011" => rgb <= "000000";
					when "11011000100010100" => rgb <= "000000";
					when "11011000100010101" => rgb <= "000000";
					when "11011000100010110" => rgb <= "000000";
					when "11011000100010111" => rgb <= "000000";
					when "11011000100011000" => rgb <= "000000";
					when "11011000100011001" => rgb <= "000000";
					when "11011000100011010" => rgb <= "000000";
					when "11011000100011011" => rgb <= "000000";
					when "11011000100011100" => rgb <= "000000";
					when "11011000100011101" => rgb <= "000000";
					when "11011000100011110" => rgb <= "000000";
					when "11011000100011111" => rgb <= "000000";
					when "11011000100100000" => rgb <= "000000";
					when "11011000100100001" => rgb <= "000000";
					when "11011000100100010" => rgb <= "000000";
					when "11011000100100011" => rgb <= "000000";
					when "11011000100100100" => rgb <= "000000";
					when "11011000100100101" => rgb <= "000000";
					when "11011000100100110" => rgb <= "000000";
					when "11011000100100111" => rgb <= "000000";
					when "11011000100101000" => rgb <= "000000";
					when "11011000100101001" => rgb <= "000000";
					when "11011000100101010" => rgb <= "000000";
					when "11011000100101011" => rgb <= "000000";
					when "11011000100101100" => rgb <= "000000";
					when "11011000100101101" => rgb <= "000000";
					when "11011000100101110" => rgb <= "000000";
					when "11011000100101111" => rgb <= "000000";
					when "11011000100110000" => rgb <= "000000";
					when "11011000100110001" => rgb <= "000000";
					when "11011000100110010" => rgb <= "000000";
					when "11011000100110011" => rgb <= "000000";
					when "11011000100110100" => rgb <= "000000";
					when "11011000100110101" => rgb <= "000000";
					when "11011000100110110" => rgb <= "000000";
					when "11011000100110111" => rgb <= "000000";
					when "11011000100111000" => rgb <= "000000";
					when "11011000100111001" => rgb <= "000000";
					when "11011000100111010" => rgb <= "000000";
					when "11011000100111011" => rgb <= "000000";
					when "11011000100111100" => rgb <= "000000";
					when "11011000100111101" => rgb <= "000000";
					when "11011000100111110" => rgb <= "000000";
					when "11011000100111111" => rgb <= "000000";
					when "11011001000000000" => rgb <= "000000";
					when "11011001000000001" => rgb <= "000000";
					when "11011001000000010" => rgb <= "000000";
					when "11011001000000011" => rgb <= "000000";
					when "11011001000000100" => rgb <= "000000";
					when "11011001000000101" => rgb <= "000000";
					when "11011001000000110" => rgb <= "000000";
					when "11011001000000111" => rgb <= "000000";
					when "11011001000001000" => rgb <= "000000";
					when "11011001000001001" => rgb <= "000000";
					when "11011001000001010" => rgb <= "000000";
					when "11011001000001011" => rgb <= "000000";
					when "11011001000001100" => rgb <= "000000";
					when "11011001000001101" => rgb <= "000000";
					when "11011001000001110" => rgb <= "000000";
					when "11011001000001111" => rgb <= "000000";
					when "11011001000010000" => rgb <= "000000";
					when "11011001000010001" => rgb <= "000000";
					when "11011001000010010" => rgb <= "000000";
					when "11011001000010011" => rgb <= "000000";
					when "11011001000010100" => rgb <= "000000";
					when "11011001000010101" => rgb <= "000000";
					when "11011001000010110" => rgb <= "000000";
					when "11011001000010111" => rgb <= "000000";
					when "11011001000011000" => rgb <= "000000";
					when "11011001000011001" => rgb <= "000000";
					when "11011001000011010" => rgb <= "000000";
					when "11011001000011011" => rgb <= "000000";
					when "11011001000011100" => rgb <= "000000";
					when "11011001000011101" => rgb <= "000000";
					when "11011001000011110" => rgb <= "000000";
					when "11011001000011111" => rgb <= "000000";
					when "11011001000100000" => rgb <= "000000";
					when "11011001000100001" => rgb <= "000000";
					when "11011001000100010" => rgb <= "000000";
					when "11011001000100011" => rgb <= "000000";
					when "11011001000100100" => rgb <= "000000";
					when "11011001000100101" => rgb <= "000000";
					when "11011001000100110" => rgb <= "000000";
					when "11011001000100111" => rgb <= "000000";
					when "11011001000101000" => rgb <= "000000";
					when "11011001000101001" => rgb <= "000000";
					when "11011001000101010" => rgb <= "000000";
					when "11011001000101011" => rgb <= "000000";
					when "11011001000101100" => rgb <= "000000";
					when "11011001000101101" => rgb <= "000000";
					when "11011001000101110" => rgb <= "000000";
					when "11011001000101111" => rgb <= "000000";
					when "11011001000110000" => rgb <= "000000";
					when "11011001000110001" => rgb <= "000000";
					when "11011001000110010" => rgb <= "000000";
					when "11011001000110011" => rgb <= "000000";
					when "11011001000110100" => rgb <= "000000";
					when "11011001000110101" => rgb <= "000000";
					when "11011001000110110" => rgb <= "000000";
					when "11011001000110111" => rgb <= "000000";
					when "11011001000111000" => rgb <= "000000";
					when "11011001000111001" => rgb <= "000000";
					when "11011001000111010" => rgb <= "000000";
					when "11011001000111011" => rgb <= "000000";
					when "11011001000111100" => rgb <= "000000";
					when "11011001000111101" => rgb <= "000000";
					when "11011001000111110" => rgb <= "000000";
					when "11011001000111111" => rgb <= "000000";
					when "11011001001000000" => rgb <= "000000";
					when "11011001001000001" => rgb <= "000000";
					when "11011001001000010" => rgb <= "000000";
					when "11011001001000011" => rgb <= "000000";
					when "11011001001000100" => rgb <= "000000";
					when "11011001001000101" => rgb <= "000000";
					when "11011001001000110" => rgb <= "000000";
					when "11011001001000111" => rgb <= "000000";
					when "11011001001001000" => rgb <= "000000";
					when "11011001001001001" => rgb <= "000000";
					when "11011001001001010" => rgb <= "000000";
					when "11011001001001011" => rgb <= "000000";
					when "11011001001001100" => rgb <= "000000";
					when "11011001001001101" => rgb <= "000000";
					when "11011001001001110" => rgb <= "000000";
					when "11011001001001111" => rgb <= "000000";
					when "11011001001010000" => rgb <= "000000";
					when "11011001001010001" => rgb <= "000000";
					when "11011001001010010" => rgb <= "000000";
					when "11011001001010011" => rgb <= "000000";
					when "11011001001010100" => rgb <= "000000";
					when "11011001001010101" => rgb <= "000000";
					when "11011001001010110" => rgb <= "000000";
					when "11011001001010111" => rgb <= "000000";
					when "11011001001011000" => rgb <= "000000";
					when "11011001001011001" => rgb <= "000000";
					when "11011001001011010" => rgb <= "000000";
					when "11011001001011011" => rgb <= "000000";
					when "11011001001011100" => rgb <= "000000";
					when "11011001001011101" => rgb <= "000000";
					when "11011001001011110" => rgb <= "000000";
					when "11011001001011111" => rgb <= "000000";
					when "11011001001100000" => rgb <= "000000";
					when "11011001001100001" => rgb <= "000000";
					when "11011001001100010" => rgb <= "000000";
					when "11011001001100011" => rgb <= "000000";
					when "11011001001100100" => rgb <= "000000";
					when "11011001001100101" => rgb <= "000000";
					when "11011001001100110" => rgb <= "000000";
					when "11011001001100111" => rgb <= "000000";
					when "11011001001101000" => rgb <= "000000";
					when "11011001001101001" => rgb <= "000000";
					when "11011001001101010" => rgb <= "000000";
					when "11011001001101011" => rgb <= "000000";
					when "11011001001101100" => rgb <= "000000";
					when "11011001001101101" => rgb <= "000000";
					when "11011001001101110" => rgb <= "000000";
					when "11011001001101111" => rgb <= "000000";
					when "11011001001110000" => rgb <= "000000";
					when "11011001001110001" => rgb <= "000000";
					when "11011001001110010" => rgb <= "000000";
					when "11011001001110011" => rgb <= "000000";
					when "11011001001110100" => rgb <= "000000";
					when "11011001001110101" => rgb <= "000000";
					when "11011001001110110" => rgb <= "000000";
					when "11011001001110111" => rgb <= "000000";
					when "11011001001111000" => rgb <= "000000";
					when "11011001001111001" => rgb <= "000000";
					when "11011001001111010" => rgb <= "000000";
					when "11011001001111011" => rgb <= "000000";
					when "11011001001111100" => rgb <= "000000";
					when "11011001001111101" => rgb <= "000000";
					when "11011001001111110" => rgb <= "000000";
					when "11011001001111111" => rgb <= "000000";
					when "11011001010000000" => rgb <= "000000";
					when "11011001010000001" => rgb <= "000000";
					when "11011001010000010" => rgb <= "000000";
					when "11011001010000011" => rgb <= "000000";
					when "11011001010000100" => rgb <= "000000";
					when "11011001010000101" => rgb <= "000000";
					when "11011001010000110" => rgb <= "000000";
					when "11011001010000111" => rgb <= "000000";
					when "11011001010001000" => rgb <= "000000";
					when "11011001010001001" => rgb <= "000000";
					when "11011001010001010" => rgb <= "000000";
					when "11011001010001011" => rgb <= "000000";
					when "11011001010001100" => rgb <= "000000";
					when "11011001010001101" => rgb <= "000000";
					when "11011001010001110" => rgb <= "000000";
					when "11011001010001111" => rgb <= "000000";
					when "11011001010010000" => rgb <= "000000";
					when "11011001010010001" => rgb <= "000000";
					when "11011001010010010" => rgb <= "000000";
					when "11011001010010011" => rgb <= "000000";
					when "11011001010010100" => rgb <= "000000";
					when "11011001010010101" => rgb <= "000000";
					when "11011001010010110" => rgb <= "000000";
					when "11011001010010111" => rgb <= "000000";
					when "11011001010011000" => rgb <= "000000";
					when "11011001010011001" => rgb <= "000000";
					when "11011001010011010" => rgb <= "000000";
					when "11011001010011011" => rgb <= "000000";
					when "11011001010011100" => rgb <= "000000";
					when "11011001010011101" => rgb <= "000000";
					when "11011001010011110" => rgb <= "000000";
					when "11011001010011111" => rgb <= "000000";
					when "11011001010100000" => rgb <= "000000";
					when "11011001010100001" => rgb <= "000000";
					when "11011001010100010" => rgb <= "000000";
					when "11011001010100011" => rgb <= "000000";
					when "11011001010100100" => rgb <= "000000";
					when "11011001010100101" => rgb <= "000000";
					when "11011001010100110" => rgb <= "000000";
					when "11011001010100111" => rgb <= "000000";
					when "11011001010101000" => rgb <= "000000";
					when "11011001010101001" => rgb <= "000000";
					when "11011001010101010" => rgb <= "000000";
					when "11011001010101011" => rgb <= "000000";
					when "11011001010101100" => rgb <= "000000";
					when "11011001010101101" => rgb <= "000000";
					when "11011001010101110" => rgb <= "000000";
					when "11011001010101111" => rgb <= "000000";
					when "11011001010110000" => rgb <= "000000";
					when "11011001010110001" => rgb <= "000000";
					when "11011001010110010" => rgb <= "000000";
					when "11011001010110011" => rgb <= "000000";
					when "11011001010110100" => rgb <= "000000";
					when "11011001010110101" => rgb <= "000000";
					when "11011001010110110" => rgb <= "000000";
					when "11011001010110111" => rgb <= "000000";
					when "11011001010111000" => rgb <= "000000";
					when "11011001010111001" => rgb <= "000000";
					when "11011001010111010" => rgb <= "000000";
					when "11011001010111011" => rgb <= "000000";
					when "11011001010111100" => rgb <= "000000";
					when "11011001010111101" => rgb <= "000000";
					when "11011001010111110" => rgb <= "000000";
					when "11011001010111111" => rgb <= "000000";
					when "11011001011000000" => rgb <= "000000";
					when "11011001011000001" => rgb <= "000000";
					when "11011001011000010" => rgb <= "000000";
					when "11011001011000011" => rgb <= "000000";
					when "11011001011000100" => rgb <= "000000";
					when "11011001011000101" => rgb <= "000000";
					when "11011001011000110" => rgb <= "000000";
					when "11011001011000111" => rgb <= "000000";
					when "11011001011001000" => rgb <= "000000";
					when "11011001011001001" => rgb <= "000000";
					when "11011001011001010" => rgb <= "000000";
					when "11011001011001011" => rgb <= "000000";
					when "11011001011001100" => rgb <= "000000";
					when "11011001011001101" => rgb <= "000000";
					when "11011001011001110" => rgb <= "000000";
					when "11011001011001111" => rgb <= "000000";
					when "11011001011010000" => rgb <= "000000";
					when "11011001011010001" => rgb <= "000000";
					when "11011001011010010" => rgb <= "000000";
					when "11011001011010011" => rgb <= "000000";
					when "11011001011010100" => rgb <= "000000";
					when "11011001011010101" => rgb <= "000000";
					when "11011001011010110" => rgb <= "000000";
					when "11011001011010111" => rgb <= "000000";
					when "11011001011011000" => rgb <= "000000";
					when "11011001011011001" => rgb <= "000000";
					when "11011001011011010" => rgb <= "000000";
					when "11011001011011011" => rgb <= "000000";
					when "11011001011011100" => rgb <= "000000";
					when "11011001011011101" => rgb <= "000000";
					when "11011001011011110" => rgb <= "000000";
					when "11011001011011111" => rgb <= "000000";
					when "11011001011100000" => rgb <= "000000";
					when "11011001011100001" => rgb <= "000000";
					when "11011001011100010" => rgb <= "000000";
					when "11011001011100011" => rgb <= "000000";
					when "11011001011100100" => rgb <= "000000";
					when "11011001011100101" => rgb <= "000000";
					when "11011001011100110" => rgb <= "000000";
					when "11011001011100111" => rgb <= "000000";
					when "11011001011101000" => rgb <= "000000";
					when "11011001011101001" => rgb <= "000000";
					when "11011001011101010" => rgb <= "000000";
					when "11011001011101011" => rgb <= "000000";
					when "11011001011101100" => rgb <= "000000";
					when "11011001011101101" => rgb <= "000000";
					when "11011001011101110" => rgb <= "000000";
					when "11011001011101111" => rgb <= "000000";
					when "11011001011110000" => rgb <= "000000";
					when "11011001011110001" => rgb <= "000000";
					when "11011001011110010" => rgb <= "000000";
					when "11011001011110011" => rgb <= "000000";
					when "11011001011110100" => rgb <= "000000";
					when "11011001011110101" => rgb <= "000000";
					when "11011001011110110" => rgb <= "000000";
					when "11011001011110111" => rgb <= "000000";
					when "11011001011111000" => rgb <= "000000";
					when "11011001011111001" => rgb <= "000000";
					when "11011001011111010" => rgb <= "000000";
					when "11011001011111011" => rgb <= "000000";
					when "11011001011111100" => rgb <= "000000";
					when "11011001011111101" => rgb <= "000000";
					when "11011001011111110" => rgb <= "000000";
					when "11011001011111111" => rgb <= "000000";
					when "11011001100000000" => rgb <= "000000";
					when "11011001100000001" => rgb <= "000000";
					when "11011001100000010" => rgb <= "000000";
					when "11011001100000011" => rgb <= "000000";
					when "11011001100000100" => rgb <= "000000";
					when "11011001100000101" => rgb <= "000000";
					when "11011001100000110" => rgb <= "000000";
					when "11011001100000111" => rgb <= "000000";
					when "11011001100001000" => rgb <= "000000";
					when "11011001100001001" => rgb <= "000000";
					when "11011001100001010" => rgb <= "000000";
					when "11011001100001011" => rgb <= "000000";
					when "11011001100001100" => rgb <= "000000";
					when "11011001100001101" => rgb <= "000000";
					when "11011001100001110" => rgb <= "000000";
					when "11011001100001111" => rgb <= "000000";
					when "11011001100010000" => rgb <= "000000";
					when "11011001100010001" => rgb <= "000000";
					when "11011001100010010" => rgb <= "000000";
					when "11011001100010011" => rgb <= "000000";
					when "11011001100010100" => rgb <= "000000";
					when "11011001100010101" => rgb <= "000000";
					when "11011001100010110" => rgb <= "000000";
					when "11011001100010111" => rgb <= "000000";
					when "11011001100011000" => rgb <= "000000";
					when "11011001100011001" => rgb <= "000000";
					when "11011001100011010" => rgb <= "000000";
					when "11011001100011011" => rgb <= "000000";
					when "11011001100011100" => rgb <= "000000";
					when "11011001100011101" => rgb <= "000000";
					when "11011001100011110" => rgb <= "000000";
					when "11011001100011111" => rgb <= "000000";
					when "11011001100100000" => rgb <= "000000";
					when "11011001100100001" => rgb <= "000000";
					when "11011001100100010" => rgb <= "000000";
					when "11011001100100011" => rgb <= "000000";
					when "11011001100100100" => rgb <= "000000";
					when "11011001100100101" => rgb <= "000000";
					when "11011001100100110" => rgb <= "000000";
					when "11011001100100111" => rgb <= "000000";
					when "11011001100101000" => rgb <= "000000";
					when "11011001100101001" => rgb <= "000000";
					when "11011001100101010" => rgb <= "000000";
					when "11011001100101011" => rgb <= "000000";
					when "11011001100101100" => rgb <= "000000";
					when "11011001100101101" => rgb <= "000000";
					when "11011001100101110" => rgb <= "000000";
					when "11011001100101111" => rgb <= "000000";
					when "11011001100110000" => rgb <= "000000";
					when "11011001100110001" => rgb <= "000000";
					when "11011001100110010" => rgb <= "000000";
					when "11011001100110011" => rgb <= "000000";
					when "11011001100110100" => rgb <= "000000";
					when "11011001100110101" => rgb <= "000000";
					when "11011001100110110" => rgb <= "000000";
					when "11011001100110111" => rgb <= "000000";
					when "11011001100111000" => rgb <= "000000";
					when "11011001100111001" => rgb <= "000000";
					when "11011001100111010" => rgb <= "000000";
					when "11011001100111011" => rgb <= "000000";
					when "11011001100111100" => rgb <= "000000";
					when "11011001100111101" => rgb <= "000000";
					when "11011001100111110" => rgb <= "000000";
					when "11011001100111111" => rgb <= "000000";
					when "11011010000000000" => rgb <= "000000";
					when "11011010000000001" => rgb <= "000000";
					when "11011010000000010" => rgb <= "000000";
					when "11011010000000011" => rgb <= "000000";
					when "11011010000000100" => rgb <= "000000";
					when "11011010000000101" => rgb <= "000000";
					when "11011010000000110" => rgb <= "000000";
					when "11011010000000111" => rgb <= "000000";
					when "11011010000001000" => rgb <= "000000";
					when "11011010000001001" => rgb <= "000000";
					when "11011010000001010" => rgb <= "000000";
					when "11011010000001011" => rgb <= "000000";
					when "11011010000001100" => rgb <= "000000";
					when "11011010000001101" => rgb <= "000000";
					when "11011010000001110" => rgb <= "000000";
					when "11011010000001111" => rgb <= "000000";
					when "11011010000010000" => rgb <= "000000";
					when "11011010000010001" => rgb <= "000000";
					when "11011010000010010" => rgb <= "000000";
					when "11011010000010011" => rgb <= "000000";
					when "11011010000010100" => rgb <= "000000";
					when "11011010000010101" => rgb <= "000000";
					when "11011010000010110" => rgb <= "000000";
					when "11011010000010111" => rgb <= "000000";
					when "11011010000011000" => rgb <= "000000";
					when "11011010000011001" => rgb <= "000000";
					when "11011010000011010" => rgb <= "000000";
					when "11011010000011011" => rgb <= "000000";
					when "11011010000011100" => rgb <= "000000";
					when "11011010000011101" => rgb <= "000000";
					when "11011010000011110" => rgb <= "000000";
					when "11011010000011111" => rgb <= "000000";
					when "11011010000100000" => rgb <= "000000";
					when "11011010000100001" => rgb <= "000000";
					when "11011010000100010" => rgb <= "000000";
					when "11011010000100011" => rgb <= "000000";
					when "11011010000100100" => rgb <= "000000";
					when "11011010000100101" => rgb <= "000000";
					when "11011010000100110" => rgb <= "000000";
					when "11011010000100111" => rgb <= "000000";
					when "11011010000101000" => rgb <= "000000";
					when "11011010000101001" => rgb <= "000000";
					when "11011010000101010" => rgb <= "000000";
					when "11011010000101011" => rgb <= "000000";
					when "11011010000101100" => rgb <= "000000";
					when "11011010000101101" => rgb <= "000000";
					when "11011010000101110" => rgb <= "000000";
					when "11011010000101111" => rgb <= "000000";
					when "11011010000110000" => rgb <= "000000";
					when "11011010000110001" => rgb <= "000000";
					when "11011010000110010" => rgb <= "000000";
					when "11011010000110011" => rgb <= "000000";
					when "11011010000110100" => rgb <= "000000";
					when "11011010000110101" => rgb <= "000000";
					when "11011010000110110" => rgb <= "000000";
					when "11011010000110111" => rgb <= "000000";
					when "11011010000111000" => rgb <= "000000";
					when "11011010000111001" => rgb <= "000000";
					when "11011010000111010" => rgb <= "000000";
					when "11011010000111011" => rgb <= "000000";
					when "11011010000111100" => rgb <= "000000";
					when "11011010000111101" => rgb <= "000000";
					when "11011010000111110" => rgb <= "000000";
					when "11011010000111111" => rgb <= "000000";
					when "11011010001000000" => rgb <= "000000";
					when "11011010001000001" => rgb <= "000000";
					when "11011010001000010" => rgb <= "000000";
					when "11011010001000011" => rgb <= "000000";
					when "11011010001000100" => rgb <= "000000";
					when "11011010001000101" => rgb <= "000000";
					when "11011010001000110" => rgb <= "000000";
					when "11011010001000111" => rgb <= "000000";
					when "11011010001001000" => rgb <= "000000";
					when "11011010001001001" => rgb <= "000000";
					when "11011010001001010" => rgb <= "000000";
					when "11011010001001011" => rgb <= "000000";
					when "11011010001001100" => rgb <= "000000";
					when "11011010001001101" => rgb <= "000000";
					when "11011010001001110" => rgb <= "000000";
					when "11011010001001111" => rgb <= "000000";
					when "11011010001010000" => rgb <= "000000";
					when "11011010001010001" => rgb <= "000000";
					when "11011010001010010" => rgb <= "000000";
					when "11011010001010011" => rgb <= "000000";
					when "11011010001010100" => rgb <= "000000";
					when "11011010001010101" => rgb <= "000000";
					when "11011010001010110" => rgb <= "000000";
					when "11011010001010111" => rgb <= "000000";
					when "11011010001011000" => rgb <= "000000";
					when "11011010001011001" => rgb <= "000000";
					when "11011010001011010" => rgb <= "000000";
					when "11011010001011011" => rgb <= "000000";
					when "11011010001011100" => rgb <= "000000";
					when "11011010001011101" => rgb <= "000000";
					when "11011010001011110" => rgb <= "000000";
					when "11011010001011111" => rgb <= "000000";
					when "11011010001100000" => rgb <= "000000";
					when "11011010001100001" => rgb <= "000000";
					when "11011010001100010" => rgb <= "000000";
					when "11011010001100011" => rgb <= "000000";
					when "11011010001100100" => rgb <= "000000";
					when "11011010001100101" => rgb <= "000000";
					when "11011010001100110" => rgb <= "000000";
					when "11011010001100111" => rgb <= "000000";
					when "11011010001101000" => rgb <= "000000";
					when "11011010001101001" => rgb <= "000000";
					when "11011010001101010" => rgb <= "000000";
					when "11011010001101011" => rgb <= "000000";
					when "11011010001101100" => rgb <= "000000";
					when "11011010001101101" => rgb <= "000000";
					when "11011010001101110" => rgb <= "000000";
					when "11011010001101111" => rgb <= "000000";
					when "11011010001110000" => rgb <= "000000";
					when "11011010001110001" => rgb <= "000000";
					when "11011010001110010" => rgb <= "000000";
					when "11011010001110011" => rgb <= "000000";
					when "11011010001110100" => rgb <= "000000";
					when "11011010001110101" => rgb <= "000000";
					when "11011010001110110" => rgb <= "000000";
					when "11011010001110111" => rgb <= "000000";
					when "11011010001111000" => rgb <= "000000";
					when "11011010001111001" => rgb <= "000000";
					when "11011010001111010" => rgb <= "000000";
					when "11011010001111011" => rgb <= "000000";
					when "11011010001111100" => rgb <= "000000";
					when "11011010001111101" => rgb <= "000000";
					when "11011010001111110" => rgb <= "000000";
					when "11011010001111111" => rgb <= "000000";
					when "11011010010000000" => rgb <= "000000";
					when "11011010010000001" => rgb <= "000000";
					when "11011010010000010" => rgb <= "000000";
					when "11011010010000011" => rgb <= "000000";
					when "11011010010000100" => rgb <= "000000";
					when "11011010010000101" => rgb <= "000000";
					when "11011010010000110" => rgb <= "000000";
					when "11011010010000111" => rgb <= "000000";
					when "11011010010001000" => rgb <= "000000";
					when "11011010010001001" => rgb <= "000000";
					when "11011010010001010" => rgb <= "000000";
					when "11011010010001011" => rgb <= "000000";
					when "11011010010001100" => rgb <= "000000";
					when "11011010010001101" => rgb <= "000000";
					when "11011010010001110" => rgb <= "000000";
					when "11011010010001111" => rgb <= "000000";
					when "11011010010010000" => rgb <= "000000";
					when "11011010010010001" => rgb <= "000000";
					when "11011010010010010" => rgb <= "000000";
					when "11011010010010011" => rgb <= "000000";
					when "11011010010010100" => rgb <= "000000";
					when "11011010010010101" => rgb <= "000000";
					when "11011010010010110" => rgb <= "000000";
					when "11011010010010111" => rgb <= "000000";
					when "11011010010011000" => rgb <= "000000";
					when "11011010010011001" => rgb <= "000000";
					when "11011010010011010" => rgb <= "000000";
					when "11011010010011011" => rgb <= "000000";
					when "11011010010011100" => rgb <= "000000";
					when "11011010010011101" => rgb <= "000000";
					when "11011010010011110" => rgb <= "000000";
					when "11011010010011111" => rgb <= "000000";
					when "11011010010100000" => rgb <= "000000";
					when "11011010010100001" => rgb <= "000000";
					when "11011010010100010" => rgb <= "000000";
					when "11011010010100011" => rgb <= "000000";
					when "11011010010100100" => rgb <= "000000";
					when "11011010010100101" => rgb <= "000000";
					when "11011010010100110" => rgb <= "000000";
					when "11011010010100111" => rgb <= "000000";
					when "11011010010101000" => rgb <= "000000";
					when "11011010010101001" => rgb <= "000000";
					when "11011010010101010" => rgb <= "000000";
					when "11011010010101011" => rgb <= "000000";
					when "11011010010101100" => rgb <= "000000";
					when "11011010010101101" => rgb <= "000000";
					when "11011010010101110" => rgb <= "000000";
					when "11011010010101111" => rgb <= "000000";
					when "11011010010110000" => rgb <= "000000";
					when "11011010010110001" => rgb <= "000000";
					when "11011010010110010" => rgb <= "000000";
					when "11011010010110011" => rgb <= "000000";
					when "11011010010110100" => rgb <= "000000";
					when "11011010010110101" => rgb <= "000000";
					when "11011010010110110" => rgb <= "000000";
					when "11011010010110111" => rgb <= "000000";
					when "11011010010111000" => rgb <= "000000";
					when "11011010010111001" => rgb <= "000000";
					when "11011010010111010" => rgb <= "000000";
					when "11011010010111011" => rgb <= "000000";
					when "11011010010111100" => rgb <= "000000";
					when "11011010010111101" => rgb <= "000000";
					when "11011010010111110" => rgb <= "000000";
					when "11011010010111111" => rgb <= "000000";
					when "11011010011000000" => rgb <= "000000";
					when "11011010011000001" => rgb <= "000000";
					when "11011010011000010" => rgb <= "000000";
					when "11011010011000011" => rgb <= "000000";
					when "11011010011000100" => rgb <= "000000";
					when "11011010011000101" => rgb <= "000000";
					when "11011010011000110" => rgb <= "000000";
					when "11011010011000111" => rgb <= "000000";
					when "11011010011001000" => rgb <= "000000";
					when "11011010011001001" => rgb <= "000000";
					when "11011010011001010" => rgb <= "000000";
					when "11011010011001011" => rgb <= "000000";
					when "11011010011001100" => rgb <= "000000";
					when "11011010011001101" => rgb <= "000000";
					when "11011010011001110" => rgb <= "000000";
					when "11011010011001111" => rgb <= "000000";
					when "11011010011010000" => rgb <= "000000";
					when "11011010011010001" => rgb <= "000000";
					when "11011010011010010" => rgb <= "000000";
					when "11011010011010011" => rgb <= "000000";
					when "11011010011010100" => rgb <= "000000";
					when "11011010011010101" => rgb <= "000000";
					when "11011010011010110" => rgb <= "000000";
					when "11011010011010111" => rgb <= "000000";
					when "11011010011011000" => rgb <= "000000";
					when "11011010011011001" => rgb <= "000000";
					when "11011010011011010" => rgb <= "000000";
					when "11011010011011011" => rgb <= "000000";
					when "11011010011011100" => rgb <= "000000";
					when "11011010011011101" => rgb <= "000000";
					when "11011010011011110" => rgb <= "000000";
					when "11011010011011111" => rgb <= "000000";
					when "11011010011100000" => rgb <= "000000";
					when "11011010011100001" => rgb <= "000000";
					when "11011010011100010" => rgb <= "000000";
					when "11011010011100011" => rgb <= "000000";
					when "11011010011100100" => rgb <= "000000";
					when "11011010011100101" => rgb <= "000000";
					when "11011010011100110" => rgb <= "000000";
					when "11011010011100111" => rgb <= "000000";
					when "11011010011101000" => rgb <= "000000";
					when "11011010011101001" => rgb <= "000000";
					when "11011010011101010" => rgb <= "000000";
					when "11011010011101011" => rgb <= "000000";
					when "11011010011101100" => rgb <= "000000";
					when "11011010011101101" => rgb <= "000000";
					when "11011010011101110" => rgb <= "000000";
					when "11011010011101111" => rgb <= "000000";
					when "11011010011110000" => rgb <= "000000";
					when "11011010011110001" => rgb <= "000000";
					when "11011010011110010" => rgb <= "000000";
					when "11011010011110011" => rgb <= "000000";
					when "11011010011110100" => rgb <= "000000";
					when "11011010011110101" => rgb <= "000000";
					when "11011010011110110" => rgb <= "000000";
					when "11011010011110111" => rgb <= "000000";
					when "11011010011111000" => rgb <= "000000";
					when "11011010011111001" => rgb <= "000000";
					when "11011010011111010" => rgb <= "000000";
					when "11011010011111011" => rgb <= "000000";
					when "11011010011111100" => rgb <= "000000";
					when "11011010011111101" => rgb <= "000000";
					when "11011010011111110" => rgb <= "000000";
					when "11011010011111111" => rgb <= "000000";
					when "11011010100000000" => rgb <= "000000";
					when "11011010100000001" => rgb <= "000000";
					when "11011010100000010" => rgb <= "000000";
					when "11011010100000011" => rgb <= "000000";
					when "11011010100000100" => rgb <= "000000";
					when "11011010100000101" => rgb <= "000000";
					when "11011010100000110" => rgb <= "000000";
					when "11011010100000111" => rgb <= "000000";
					when "11011010100001000" => rgb <= "000000";
					when "11011010100001001" => rgb <= "000000";
					when "11011010100001010" => rgb <= "000000";
					when "11011010100001011" => rgb <= "000000";
					when "11011010100001100" => rgb <= "000000";
					when "11011010100001101" => rgb <= "000000";
					when "11011010100001110" => rgb <= "000000";
					when "11011010100001111" => rgb <= "000000";
					when "11011010100010000" => rgb <= "000000";
					when "11011010100010001" => rgb <= "000000";
					when "11011010100010010" => rgb <= "000000";
					when "11011010100010011" => rgb <= "000000";
					when "11011010100010100" => rgb <= "000000";
					when "11011010100010101" => rgb <= "000000";
					when "11011010100010110" => rgb <= "000000";
					when "11011010100010111" => rgb <= "000000";
					when "11011010100011000" => rgb <= "000000";
					when "11011010100011001" => rgb <= "000000";
					when "11011010100011010" => rgb <= "000000";
					when "11011010100011011" => rgb <= "000000";
					when "11011010100011100" => rgb <= "000000";
					when "11011010100011101" => rgb <= "000000";
					when "11011010100011110" => rgb <= "000000";
					when "11011010100011111" => rgb <= "000000";
					when "11011010100100000" => rgb <= "000000";
					when "11011010100100001" => rgb <= "000000";
					when "11011010100100010" => rgb <= "000000";
					when "11011010100100011" => rgb <= "000000";
					when "11011010100100100" => rgb <= "000000";
					when "11011010100100101" => rgb <= "000000";
					when "11011010100100110" => rgb <= "000000";
					when "11011010100100111" => rgb <= "000000";
					when "11011010100101000" => rgb <= "000000";
					when "11011010100101001" => rgb <= "000000";
					when "11011010100101010" => rgb <= "000000";
					when "11011010100101011" => rgb <= "000000";
					when "11011010100101100" => rgb <= "000000";
					when "11011010100101101" => rgb <= "000000";
					when "11011010100101110" => rgb <= "000000";
					when "11011010100101111" => rgb <= "000000";
					when "11011010100110000" => rgb <= "000000";
					when "11011010100110001" => rgb <= "000000";
					when "11011010100110010" => rgb <= "000000";
					when "11011010100110011" => rgb <= "000000";
					when "11011010100110100" => rgb <= "000000";
					when "11011010100110101" => rgb <= "000000";
					when "11011010100110110" => rgb <= "000000";
					when "11011010100110111" => rgb <= "000000";
					when "11011010100111000" => rgb <= "000000";
					when "11011010100111001" => rgb <= "000000";
					when "11011010100111010" => rgb <= "000000";
					when "11011010100111011" => rgb <= "000000";
					when "11011010100111100" => rgb <= "000000";
					when "11011010100111101" => rgb <= "000000";
					when "11011010100111110" => rgb <= "000000";
					when "11011010100111111" => rgb <= "000000";
					when "11011011000000000" => rgb <= "000000";
					when "11011011000000001" => rgb <= "000000";
					when "11011011000000010" => rgb <= "000000";
					when "11011011000000011" => rgb <= "000000";
					when "11011011000000100" => rgb <= "000000";
					when "11011011000000101" => rgb <= "000000";
					when "11011011000000110" => rgb <= "000000";
					when "11011011000000111" => rgb <= "000000";
					when "11011011000001000" => rgb <= "000000";
					when "11011011000001001" => rgb <= "000000";
					when "11011011000001010" => rgb <= "000000";
					when "11011011000001011" => rgb <= "000000";
					when "11011011000001100" => rgb <= "000000";
					when "11011011000001101" => rgb <= "000000";
					when "11011011000001110" => rgb <= "000000";
					when "11011011000001111" => rgb <= "000000";
					when "11011011000010000" => rgb <= "000000";
					when "11011011000010001" => rgb <= "000000";
					when "11011011000010010" => rgb <= "000000";
					when "11011011000010011" => rgb <= "000000";
					when "11011011000010100" => rgb <= "000000";
					when "11011011000010101" => rgb <= "000000";
					when "11011011000010110" => rgb <= "000000";
					when "11011011000010111" => rgb <= "000000";
					when "11011011000011000" => rgb <= "000000";
					when "11011011000011001" => rgb <= "000000";
					when "11011011000011010" => rgb <= "000000";
					when "11011011000011011" => rgb <= "000000";
					when "11011011000011100" => rgb <= "000000";
					when "11011011000011101" => rgb <= "000000";
					when "11011011000011110" => rgb <= "000000";
					when "11011011000011111" => rgb <= "000000";
					when "11011011000100000" => rgb <= "000000";
					when "11011011000100001" => rgb <= "000000";
					when "11011011000100010" => rgb <= "000000";
					when "11011011000100011" => rgb <= "000000";
					when "11011011000100100" => rgb <= "000000";
					when "11011011000100101" => rgb <= "000000";
					when "11011011000100110" => rgb <= "000000";
					when "11011011000100111" => rgb <= "000000";
					when "11011011000101000" => rgb <= "000000";
					when "11011011000101001" => rgb <= "000000";
					when "11011011000101010" => rgb <= "000000";
					when "11011011000101011" => rgb <= "000000";
					when "11011011000101100" => rgb <= "000000";
					when "11011011000101101" => rgb <= "000000";
					when "11011011000101110" => rgb <= "000000";
					when "11011011000101111" => rgb <= "000000";
					when "11011011000110000" => rgb <= "000000";
					when "11011011000110001" => rgb <= "000000";
					when "11011011000110010" => rgb <= "000000";
					when "11011011000110011" => rgb <= "000000";
					when "11011011000110100" => rgb <= "000000";
					when "11011011000110101" => rgb <= "000000";
					when "11011011000110110" => rgb <= "000000";
					when "11011011000110111" => rgb <= "000000";
					when "11011011000111000" => rgb <= "000000";
					when "11011011000111001" => rgb <= "000000";
					when "11011011000111010" => rgb <= "000000";
					when "11011011000111011" => rgb <= "000000";
					when "11011011000111100" => rgb <= "000000";
					when "11011011000111101" => rgb <= "000000";
					when "11011011000111110" => rgb <= "000000";
					when "11011011000111111" => rgb <= "000000";
					when "11011011001000000" => rgb <= "000000";
					when "11011011001000001" => rgb <= "000000";
					when "11011011001000010" => rgb <= "000000";
					when "11011011001000011" => rgb <= "000000";
					when "11011011001000100" => rgb <= "000000";
					when "11011011001000101" => rgb <= "000000";
					when "11011011001000110" => rgb <= "000000";
					when "11011011001000111" => rgb <= "000000";
					when "11011011001001000" => rgb <= "000000";
					when "11011011001001001" => rgb <= "000000";
					when "11011011001001010" => rgb <= "000000";
					when "11011011001001011" => rgb <= "000000";
					when "11011011001001100" => rgb <= "000000";
					when "11011011001001101" => rgb <= "000000";
					when "11011011001001110" => rgb <= "000000";
					when "11011011001001111" => rgb <= "000000";
					when "11011011001010000" => rgb <= "000000";
					when "11011011001010001" => rgb <= "000000";
					when "11011011001010010" => rgb <= "000000";
					when "11011011001010011" => rgb <= "000000";
					when "11011011001010100" => rgb <= "000000";
					when "11011011001010101" => rgb <= "000000";
					when "11011011001010110" => rgb <= "000000";
					when "11011011001010111" => rgb <= "000000";
					when "11011011001011000" => rgb <= "000000";
					when "11011011001011001" => rgb <= "000000";
					when "11011011001011010" => rgb <= "000000";
					when "11011011001011011" => rgb <= "000000";
					when "11011011001011100" => rgb <= "000000";
					when "11011011001011101" => rgb <= "000000";
					when "11011011001011110" => rgb <= "000000";
					when "11011011001011111" => rgb <= "000000";
					when "11011011001100000" => rgb <= "000000";
					when "11011011001100001" => rgb <= "000000";
					when "11011011001100010" => rgb <= "000000";
					when "11011011001100011" => rgb <= "000000";
					when "11011011001100100" => rgb <= "000000";
					when "11011011001100101" => rgb <= "000000";
					when "11011011001100110" => rgb <= "000000";
					when "11011011001100111" => rgb <= "000000";
					when "11011011001101000" => rgb <= "000000";
					when "11011011001101001" => rgb <= "000000";
					when "11011011001101010" => rgb <= "000000";
					when "11011011001101011" => rgb <= "000000";
					when "11011011001101100" => rgb <= "000000";
					when "11011011001101101" => rgb <= "000000";
					when "11011011001101110" => rgb <= "000000";
					when "11011011001101111" => rgb <= "000000";
					when "11011011001110000" => rgb <= "000000";
					when "11011011001110001" => rgb <= "000000";
					when "11011011001110010" => rgb <= "000000";
					when "11011011001110011" => rgb <= "000000";
					when "11011011001110100" => rgb <= "000000";
					when "11011011001110101" => rgb <= "000000";
					when "11011011001110110" => rgb <= "000000";
					when "11011011001110111" => rgb <= "000000";
					when "11011011001111000" => rgb <= "000000";
					when "11011011001111001" => rgb <= "000000";
					when "11011011001111010" => rgb <= "000000";
					when "11011011001111011" => rgb <= "000000";
					when "11011011001111100" => rgb <= "000000";
					when "11011011001111101" => rgb <= "000000";
					when "11011011001111110" => rgb <= "000000";
					when "11011011001111111" => rgb <= "000000";
					when "11011011010000000" => rgb <= "000000";
					when "11011011010000001" => rgb <= "000000";
					when "11011011010000010" => rgb <= "000000";
					when "11011011010000011" => rgb <= "000000";
					when "11011011010000100" => rgb <= "000000";
					when "11011011010000101" => rgb <= "000000";
					when "11011011010000110" => rgb <= "000000";
					when "11011011010000111" => rgb <= "000000";
					when "11011011010001000" => rgb <= "000000";
					when "11011011010001001" => rgb <= "000000";
					when "11011011010001010" => rgb <= "000000";
					when "11011011010001011" => rgb <= "000000";
					when "11011011010001100" => rgb <= "000000";
					when "11011011010001101" => rgb <= "000000";
					when "11011011010001110" => rgb <= "000000";
					when "11011011010001111" => rgb <= "000000";
					when "11011011010010000" => rgb <= "000000";
					when "11011011010010001" => rgb <= "000000";
					when "11011011010010010" => rgb <= "000000";
					when "11011011010010011" => rgb <= "000000";
					when "11011011010010100" => rgb <= "000000";
					when "11011011010010101" => rgb <= "000000";
					when "11011011010010110" => rgb <= "000000";
					when "11011011010010111" => rgb <= "000000";
					when "11011011010011000" => rgb <= "000000";
					when "11011011010011001" => rgb <= "000000";
					when "11011011010011010" => rgb <= "000000";
					when "11011011010011011" => rgb <= "000000";
					when "11011011010011100" => rgb <= "000000";
					when "11011011010011101" => rgb <= "000000";
					when "11011011010011110" => rgb <= "000000";
					when "11011011010011111" => rgb <= "000000";
					when "11011011010100000" => rgb <= "000000";
					when "11011011010100001" => rgb <= "000000";
					when "11011011010100010" => rgb <= "000000";
					when "11011011010100011" => rgb <= "000000";
					when "11011011010100100" => rgb <= "000000";
					when "11011011010100101" => rgb <= "000000";
					when "11011011010100110" => rgb <= "000000";
					when "11011011010100111" => rgb <= "000000";
					when "11011011010101000" => rgb <= "000000";
					when "11011011010101001" => rgb <= "000000";
					when "11011011010101010" => rgb <= "000000";
					when "11011011010101011" => rgb <= "000000";
					when "11011011010101100" => rgb <= "000000";
					when "11011011010101101" => rgb <= "000000";
					when "11011011010101110" => rgb <= "000000";
					when "11011011010101111" => rgb <= "000000";
					when "11011011010110000" => rgb <= "000000";
					when "11011011010110001" => rgb <= "000000";
					when "11011011010110010" => rgb <= "000000";
					when "11011011010110011" => rgb <= "000000";
					when "11011011010110100" => rgb <= "000000";
					when "11011011010110101" => rgb <= "000000";
					when "11011011010110110" => rgb <= "000000";
					when "11011011010110111" => rgb <= "000000";
					when "11011011010111000" => rgb <= "000000";
					when "11011011010111001" => rgb <= "000000";
					when "11011011010111010" => rgb <= "000000";
					when "11011011010111011" => rgb <= "000000";
					when "11011011010111100" => rgb <= "000000";
					when "11011011010111101" => rgb <= "000000";
					when "11011011010111110" => rgb <= "000000";
					when "11011011010111111" => rgb <= "000000";
					when "11011011011000000" => rgb <= "000000";
					when "11011011011000001" => rgb <= "000000";
					when "11011011011000010" => rgb <= "000000";
					when "11011011011000011" => rgb <= "000000";
					when "11011011011000100" => rgb <= "000000";
					when "11011011011000101" => rgb <= "000000";
					when "11011011011000110" => rgb <= "000000";
					when "11011011011000111" => rgb <= "000000";
					when "11011011011001000" => rgb <= "000000";
					when "11011011011001001" => rgb <= "000000";
					when "11011011011001010" => rgb <= "000000";
					when "11011011011001011" => rgb <= "000000";
					when "11011011011001100" => rgb <= "000000";
					when "11011011011001101" => rgb <= "000000";
					when "11011011011001110" => rgb <= "000000";
					when "11011011011001111" => rgb <= "000000";
					when "11011011011010000" => rgb <= "000000";
					when "11011011011010001" => rgb <= "000000";
					when "11011011011010010" => rgb <= "000000";
					when "11011011011010011" => rgb <= "000000";
					when "11011011011010100" => rgb <= "000000";
					when "11011011011010101" => rgb <= "000000";
					when "11011011011010110" => rgb <= "000000";
					when "11011011011010111" => rgb <= "000000";
					when "11011011011011000" => rgb <= "000000";
					when "11011011011011001" => rgb <= "000000";
					when "11011011011011010" => rgb <= "000000";
					when "11011011011011011" => rgb <= "000000";
					when "11011011011011100" => rgb <= "000000";
					when "11011011011011101" => rgb <= "000000";
					when "11011011011011110" => rgb <= "000000";
					when "11011011011011111" => rgb <= "000000";
					when "11011011011100000" => rgb <= "000000";
					when "11011011011100001" => rgb <= "000000";
					when "11011011011100010" => rgb <= "000000";
					when "11011011011100011" => rgb <= "000000";
					when "11011011011100100" => rgb <= "000000";
					when "11011011011100101" => rgb <= "000000";
					when "11011011011100110" => rgb <= "000000";
					when "11011011011100111" => rgb <= "000000";
					when "11011011011101000" => rgb <= "000000";
					when "11011011011101001" => rgb <= "000000";
					when "11011011011101010" => rgb <= "000000";
					when "11011011011101011" => rgb <= "000000";
					when "11011011011101100" => rgb <= "000000";
					when "11011011011101101" => rgb <= "000000";
					when "11011011011101110" => rgb <= "000000";
					when "11011011011101111" => rgb <= "000000";
					when "11011011011110000" => rgb <= "000000";
					when "11011011011110001" => rgb <= "000000";
					when "11011011011110010" => rgb <= "000000";
					when "11011011011110011" => rgb <= "000000";
					when "11011011011110100" => rgb <= "000000";
					when "11011011011110101" => rgb <= "000000";
					when "11011011011110110" => rgb <= "000000";
					when "11011011011110111" => rgb <= "000000";
					when "11011011011111000" => rgb <= "000000";
					when "11011011011111001" => rgb <= "000000";
					when "11011011011111010" => rgb <= "000000";
					when "11011011011111011" => rgb <= "000000";
					when "11011011011111100" => rgb <= "000000";
					when "11011011011111101" => rgb <= "000000";
					when "11011011011111110" => rgb <= "000000";
					when "11011011011111111" => rgb <= "000000";
					when "11011011100000000" => rgb <= "000000";
					when "11011011100000001" => rgb <= "000000";
					when "11011011100000010" => rgb <= "000000";
					when "11011011100000011" => rgb <= "000000";
					when "11011011100000100" => rgb <= "000000";
					when "11011011100000101" => rgb <= "000000";
					when "11011011100000110" => rgb <= "000000";
					when "11011011100000111" => rgb <= "000000";
					when "11011011100001000" => rgb <= "000000";
					when "11011011100001001" => rgb <= "000000";
					when "11011011100001010" => rgb <= "000000";
					when "11011011100001011" => rgb <= "000000";
					when "11011011100001100" => rgb <= "000000";
					when "11011011100001101" => rgb <= "000000";
					when "11011011100001110" => rgb <= "000000";
					when "11011011100001111" => rgb <= "000000";
					when "11011011100010000" => rgb <= "000000";
					when "11011011100010001" => rgb <= "000000";
					when "11011011100010010" => rgb <= "000000";
					when "11011011100010011" => rgb <= "000000";
					when "11011011100010100" => rgb <= "000000";
					when "11011011100010101" => rgb <= "000000";
					when "11011011100010110" => rgb <= "000000";
					when "11011011100010111" => rgb <= "000000";
					when "11011011100011000" => rgb <= "000000";
					when "11011011100011001" => rgb <= "000000";
					when "11011011100011010" => rgb <= "000000";
					when "11011011100011011" => rgb <= "000000";
					when "11011011100011100" => rgb <= "000000";
					when "11011011100011101" => rgb <= "000000";
					when "11011011100011110" => rgb <= "000000";
					when "11011011100011111" => rgb <= "000000";
					when "11011011100100000" => rgb <= "000000";
					when "11011011100100001" => rgb <= "000000";
					when "11011011100100010" => rgb <= "000000";
					when "11011011100100011" => rgb <= "000000";
					when "11011011100100100" => rgb <= "000000";
					when "11011011100100101" => rgb <= "000000";
					when "11011011100100110" => rgb <= "000000";
					when "11011011100100111" => rgb <= "000000";
					when "11011011100101000" => rgb <= "000000";
					when "11011011100101001" => rgb <= "000000";
					when "11011011100101010" => rgb <= "000000";
					when "11011011100101011" => rgb <= "000000";
					when "11011011100101100" => rgb <= "000000";
					when "11011011100101101" => rgb <= "000000";
					when "11011011100101110" => rgb <= "000000";
					when "11011011100101111" => rgb <= "000000";
					when "11011011100110000" => rgb <= "000000";
					when "11011011100110001" => rgb <= "000000";
					when "11011011100110010" => rgb <= "000000";
					when "11011011100110011" => rgb <= "000000";
					when "11011011100110100" => rgb <= "000000";
					when "11011011100110101" => rgb <= "000000";
					when "11011011100110110" => rgb <= "000000";
					when "11011011100110111" => rgb <= "000000";
					when "11011011100111000" => rgb <= "000000";
					when "11011011100111001" => rgb <= "000000";
					when "11011011100111010" => rgb <= "000000";
					when "11011011100111011" => rgb <= "000000";
					when "11011011100111100" => rgb <= "000000";
					when "11011011100111101" => rgb <= "000000";
					when "11011011100111110" => rgb <= "000000";
					when "11011011100111111" => rgb <= "000000";
					when "11011100000000000" => rgb <= "000000";
					when "11011100000000001" => rgb <= "000000";
					when "11011100000000010" => rgb <= "000000";
					when "11011100000000011" => rgb <= "000000";
					when "11011100000000100" => rgb <= "000000";
					when "11011100000000101" => rgb <= "000000";
					when "11011100000000110" => rgb <= "000000";
					when "11011100000000111" => rgb <= "000000";
					when "11011100000001000" => rgb <= "000000";
					when "11011100000001001" => rgb <= "000000";
					when "11011100000001010" => rgb <= "000000";
					when "11011100000001011" => rgb <= "000000";
					when "11011100000001100" => rgb <= "000000";
					when "11011100000001101" => rgb <= "000000";
					when "11011100000001110" => rgb <= "000000";
					when "11011100000001111" => rgb <= "000000";
					when "11011100000010000" => rgb <= "000000";
					when "11011100000010001" => rgb <= "000000";
					when "11011100000010010" => rgb <= "000000";
					when "11011100000010011" => rgb <= "000000";
					when "11011100000010100" => rgb <= "000000";
					when "11011100000010101" => rgb <= "000000";
					when "11011100000010110" => rgb <= "000000";
					when "11011100000010111" => rgb <= "000000";
					when "11011100000011000" => rgb <= "000000";
					when "11011100000011001" => rgb <= "000000";
					when "11011100000011010" => rgb <= "000000";
					when "11011100000011011" => rgb <= "000000";
					when "11011100000011100" => rgb <= "000000";
					when "11011100000011101" => rgb <= "000000";
					when "11011100000011110" => rgb <= "000000";
					when "11011100000011111" => rgb <= "000000";
					when "11011100000100000" => rgb <= "000000";
					when "11011100000100001" => rgb <= "000000";
					when "11011100000100010" => rgb <= "000000";
					when "11011100000100011" => rgb <= "000000";
					when "11011100000100100" => rgb <= "000000";
					when "11011100000100101" => rgb <= "000000";
					when "11011100000100110" => rgb <= "000000";
					when "11011100000100111" => rgb <= "000000";
					when "11011100000101000" => rgb <= "000000";
					when "11011100000101001" => rgb <= "000000";
					when "11011100000101010" => rgb <= "000000";
					when "11011100000101011" => rgb <= "000000";
					when "11011100000101100" => rgb <= "000000";
					when "11011100000101101" => rgb <= "000000";
					when "11011100000101110" => rgb <= "000000";
					when "11011100000101111" => rgb <= "000000";
					when "11011100000110000" => rgb <= "000000";
					when "11011100000110001" => rgb <= "000000";
					when "11011100000110010" => rgb <= "000000";
					when "11011100000110011" => rgb <= "000000";
					when "11011100000110100" => rgb <= "000000";
					when "11011100000110101" => rgb <= "000000";
					when "11011100000110110" => rgb <= "000000";
					when "11011100000110111" => rgb <= "000000";
					when "11011100000111000" => rgb <= "000000";
					when "11011100000111001" => rgb <= "000000";
					when "11011100000111010" => rgb <= "000000";
					when "11011100000111011" => rgb <= "000000";
					when "11011100000111100" => rgb <= "000000";
					when "11011100000111101" => rgb <= "000000";
					when "11011100000111110" => rgb <= "000000";
					when "11011100000111111" => rgb <= "000000";
					when "11011100001000000" => rgb <= "000000";
					when "11011100001000001" => rgb <= "000000";
					when "11011100001000010" => rgb <= "000000";
					when "11011100001000011" => rgb <= "000000";
					when "11011100001000100" => rgb <= "000000";
					when "11011100001000101" => rgb <= "000000";
					when "11011100001000110" => rgb <= "000000";
					when "11011100001000111" => rgb <= "000000";
					when "11011100001001000" => rgb <= "000000";
					when "11011100001001001" => rgb <= "000000";
					when "11011100001001010" => rgb <= "000000";
					when "11011100001001011" => rgb <= "000000";
					when "11011100001001100" => rgb <= "000000";
					when "11011100001001101" => rgb <= "000000";
					when "11011100001001110" => rgb <= "000000";
					when "11011100001001111" => rgb <= "000000";
					when "11011100001010000" => rgb <= "000000";
					when "11011100001010001" => rgb <= "000000";
					when "11011100001010010" => rgb <= "000000";
					when "11011100001010011" => rgb <= "000000";
					when "11011100001010100" => rgb <= "000000";
					when "11011100001010101" => rgb <= "000000";
					when "11011100001010110" => rgb <= "000000";
					when "11011100001010111" => rgb <= "000000";
					when "11011100001011000" => rgb <= "000000";
					when "11011100001011001" => rgb <= "000000";
					when "11011100001011010" => rgb <= "000000";
					when "11011100001011011" => rgb <= "000000";
					when "11011100001011100" => rgb <= "000000";
					when "11011100001011101" => rgb <= "000000";
					when "11011100001011110" => rgb <= "000000";
					when "11011100001011111" => rgb <= "000000";
					when "11011100001100000" => rgb <= "000000";
					when "11011100001100001" => rgb <= "000000";
					when "11011100001100010" => rgb <= "000000";
					when "11011100001100011" => rgb <= "000000";
					when "11011100001100100" => rgb <= "000000";
					when "11011100001100101" => rgb <= "000000";
					when "11011100001100110" => rgb <= "000000";
					when "11011100001100111" => rgb <= "000000";
					when "11011100001101000" => rgb <= "000000";
					when "11011100001101001" => rgb <= "000000";
					when "11011100001101010" => rgb <= "000000";
					when "11011100001101011" => rgb <= "000000";
					when "11011100001101100" => rgb <= "000000";
					when "11011100001101101" => rgb <= "000000";
					when "11011100001101110" => rgb <= "000000";
					when "11011100001101111" => rgb <= "000000";
					when "11011100001110000" => rgb <= "000000";
					when "11011100001110001" => rgb <= "000000";
					when "11011100001110010" => rgb <= "000000";
					when "11011100001110011" => rgb <= "000000";
					when "11011100001110100" => rgb <= "000000";
					when "11011100001110101" => rgb <= "000000";
					when "11011100001110110" => rgb <= "000000";
					when "11011100001110111" => rgb <= "000000";
					when "11011100001111000" => rgb <= "000000";
					when "11011100001111001" => rgb <= "000000";
					when "11011100001111010" => rgb <= "000000";
					when "11011100001111011" => rgb <= "000000";
					when "11011100001111100" => rgb <= "000000";
					when "11011100001111101" => rgb <= "000000";
					when "11011100001111110" => rgb <= "000000";
					when "11011100001111111" => rgb <= "000000";
					when "11011100010000000" => rgb <= "000000";
					when "11011100010000001" => rgb <= "000000";
					when "11011100010000010" => rgb <= "000000";
					when "11011100010000011" => rgb <= "000000";
					when "11011100010000100" => rgb <= "000000";
					when "11011100010000101" => rgb <= "000000";
					when "11011100010000110" => rgb <= "000000";
					when "11011100010000111" => rgb <= "000000";
					when "11011100010001000" => rgb <= "000000";
					when "11011100010001001" => rgb <= "000000";
					when "11011100010001010" => rgb <= "000000";
					when "11011100010001011" => rgb <= "000000";
					when "11011100010001100" => rgb <= "000000";
					when "11011100010001101" => rgb <= "000000";
					when "11011100010001110" => rgb <= "000000";
					when "11011100010001111" => rgb <= "000000";
					when "11011100010010000" => rgb <= "000000";
					when "11011100010010001" => rgb <= "000000";
					when "11011100010010010" => rgb <= "000000";
					when "11011100010010011" => rgb <= "000000";
					when "11011100010010100" => rgb <= "000000";
					when "11011100010010101" => rgb <= "000000";
					when "11011100010010110" => rgb <= "000000";
					when "11011100010010111" => rgb <= "000000";
					when "11011100010011000" => rgb <= "000000";
					when "11011100010011001" => rgb <= "000000";
					when "11011100010011010" => rgb <= "000000";
					when "11011100010011011" => rgb <= "000000";
					when "11011100010011100" => rgb <= "000000";
					when "11011100010011101" => rgb <= "000000";
					when "11011100010011110" => rgb <= "000000";
					when "11011100010011111" => rgb <= "000000";
					when "11011100010100000" => rgb <= "000000";
					when "11011100010100001" => rgb <= "000000";
					when "11011100010100010" => rgb <= "000000";
					when "11011100010100011" => rgb <= "000000";
					when "11011100010100100" => rgb <= "000000";
					when "11011100010100101" => rgb <= "000000";
					when "11011100010100110" => rgb <= "000000";
					when "11011100010100111" => rgb <= "000000";
					when "11011100010101000" => rgb <= "000000";
					when "11011100010101001" => rgb <= "000000";
					when "11011100010101010" => rgb <= "000000";
					when "11011100010101011" => rgb <= "000000";
					when "11011100010101100" => rgb <= "000000";
					when "11011100010101101" => rgb <= "000000";
					when "11011100010101110" => rgb <= "000000";
					when "11011100010101111" => rgb <= "000000";
					when "11011100010110000" => rgb <= "000000";
					when "11011100010110001" => rgb <= "000000";
					when "11011100010110010" => rgb <= "000000";
					when "11011100010110011" => rgb <= "000000";
					when "11011100010110100" => rgb <= "000000";
					when "11011100010110101" => rgb <= "000000";
					when "11011100010110110" => rgb <= "000000";
					when "11011100010110111" => rgb <= "000000";
					when "11011100010111000" => rgb <= "000000";
					when "11011100010111001" => rgb <= "000000";
					when "11011100010111010" => rgb <= "000000";
					when "11011100010111011" => rgb <= "000000";
					when "11011100010111100" => rgb <= "000000";
					when "11011100010111101" => rgb <= "000000";
					when "11011100010111110" => rgb <= "000000";
					when "11011100010111111" => rgb <= "000000";
					when "11011100011000000" => rgb <= "000000";
					when "11011100011000001" => rgb <= "000000";
					when "11011100011000010" => rgb <= "000000";
					when "11011100011000011" => rgb <= "000000";
					when "11011100011000100" => rgb <= "000000";
					when "11011100011000101" => rgb <= "000000";
					when "11011100011000110" => rgb <= "000000";
					when "11011100011000111" => rgb <= "000000";
					when "11011100011001000" => rgb <= "000000";
					when "11011100011001001" => rgb <= "000000";
					when "11011100011001010" => rgb <= "000000";
					when "11011100011001011" => rgb <= "000000";
					when "11011100011001100" => rgb <= "000000";
					when "11011100011001101" => rgb <= "000000";
					when "11011100011001110" => rgb <= "000000";
					when "11011100011001111" => rgb <= "000000";
					when "11011100011010000" => rgb <= "000000";
					when "11011100011010001" => rgb <= "000000";
					when "11011100011010010" => rgb <= "000000";
					when "11011100011010011" => rgb <= "000000";
					when "11011100011010100" => rgb <= "000000";
					when "11011100011010101" => rgb <= "000000";
					when "11011100011010110" => rgb <= "000000";
					when "11011100011010111" => rgb <= "000000";
					when "11011100011011000" => rgb <= "000000";
					when "11011100011011001" => rgb <= "000000";
					when "11011100011011010" => rgb <= "000000";
					when "11011100011011011" => rgb <= "000000";
					when "11011100011011100" => rgb <= "000000";
					when "11011100011011101" => rgb <= "000000";
					when "11011100011011110" => rgb <= "000000";
					when "11011100011011111" => rgb <= "000000";
					when "11011100011100000" => rgb <= "000000";
					when "11011100011100001" => rgb <= "000000";
					when "11011100011100010" => rgb <= "000000";
					when "11011100011100011" => rgb <= "000000";
					when "11011100011100100" => rgb <= "000000";
					when "11011100011100101" => rgb <= "000000";
					when "11011100011100110" => rgb <= "000000";
					when "11011100011100111" => rgb <= "000000";
					when "11011100011101000" => rgb <= "000000";
					when "11011100011101001" => rgb <= "000000";
					when "11011100011101010" => rgb <= "000000";
					when "11011100011101011" => rgb <= "000000";
					when "11011100011101100" => rgb <= "000000";
					when "11011100011101101" => rgb <= "000000";
					when "11011100011101110" => rgb <= "000000";
					when "11011100011101111" => rgb <= "000000";
					when "11011100011110000" => rgb <= "000000";
					when "11011100011110001" => rgb <= "000000";
					when "11011100011110010" => rgb <= "000000";
					when "11011100011110011" => rgb <= "000000";
					when "11011100011110100" => rgb <= "000000";
					when "11011100011110101" => rgb <= "000000";
					when "11011100011110110" => rgb <= "000000";
					when "11011100011110111" => rgb <= "000000";
					when "11011100011111000" => rgb <= "000000";
					when "11011100011111001" => rgb <= "000000";
					when "11011100011111010" => rgb <= "000000";
					when "11011100011111011" => rgb <= "000000";
					when "11011100011111100" => rgb <= "000000";
					when "11011100011111101" => rgb <= "000000";
					when "11011100011111110" => rgb <= "000000";
					when "11011100011111111" => rgb <= "000000";
					when "11011100100000000" => rgb <= "000000";
					when "11011100100000001" => rgb <= "000000";
					when "11011100100000010" => rgb <= "000000";
					when "11011100100000011" => rgb <= "000000";
					when "11011100100000100" => rgb <= "000000";
					when "11011100100000101" => rgb <= "000000";
					when "11011100100000110" => rgb <= "000000";
					when "11011100100000111" => rgb <= "000000";
					when "11011100100001000" => rgb <= "000000";
					when "11011100100001001" => rgb <= "000000";
					when "11011100100001010" => rgb <= "000000";
					when "11011100100001011" => rgb <= "000000";
					when "11011100100001100" => rgb <= "000000";
					when "11011100100001101" => rgb <= "000000";
					when "11011100100001110" => rgb <= "000000";
					when "11011100100001111" => rgb <= "000000";
					when "11011100100010000" => rgb <= "000000";
					when "11011100100010001" => rgb <= "000000";
					when "11011100100010010" => rgb <= "000000";
					when "11011100100010011" => rgb <= "000000";
					when "11011100100010100" => rgb <= "000000";
					when "11011100100010101" => rgb <= "000000";
					when "11011100100010110" => rgb <= "000000";
					when "11011100100010111" => rgb <= "000000";
					when "11011100100011000" => rgb <= "000000";
					when "11011100100011001" => rgb <= "000000";
					when "11011100100011010" => rgb <= "000000";
					when "11011100100011011" => rgb <= "000000";
					when "11011100100011100" => rgb <= "000000";
					when "11011100100011101" => rgb <= "000000";
					when "11011100100011110" => rgb <= "000000";
					when "11011100100011111" => rgb <= "000000";
					when "11011100100100000" => rgb <= "000000";
					when "11011100100100001" => rgb <= "000000";
					when "11011100100100010" => rgb <= "000000";
					when "11011100100100011" => rgb <= "000000";
					when "11011100100100100" => rgb <= "000000";
					when "11011100100100101" => rgb <= "000000";
					when "11011100100100110" => rgb <= "000000";
					when "11011100100100111" => rgb <= "000000";
					when "11011100100101000" => rgb <= "000000";
					when "11011100100101001" => rgb <= "000000";
					when "11011100100101010" => rgb <= "000000";
					when "11011100100101011" => rgb <= "000000";
					when "11011100100101100" => rgb <= "000000";
					when "11011100100101101" => rgb <= "000000";
					when "11011100100101110" => rgb <= "000000";
					when "11011100100101111" => rgb <= "000000";
					when "11011100100110000" => rgb <= "000000";
					when "11011100100110001" => rgb <= "000000";
					when "11011100100110010" => rgb <= "000000";
					when "11011100100110011" => rgb <= "000000";
					when "11011100100110100" => rgb <= "000000";
					when "11011100100110101" => rgb <= "000000";
					when "11011100100110110" => rgb <= "000000";
					when "11011100100110111" => rgb <= "000000";
					when "11011100100111000" => rgb <= "000000";
					when "11011100100111001" => rgb <= "000000";
					when "11011100100111010" => rgb <= "000000";
					when "11011100100111011" => rgb <= "000000";
					when "11011100100111100" => rgb <= "000000";
					when "11011100100111101" => rgb <= "000000";
					when "11011100100111110" => rgb <= "000000";
					when "11011100100111111" => rgb <= "000000";
					when "11011101000000000" => rgb <= "000000";
					when "11011101000000001" => rgb <= "000000";
					when "11011101000000010" => rgb <= "000000";
					when "11011101000000011" => rgb <= "000000";
					when "11011101000000100" => rgb <= "000000";
					when "11011101000000101" => rgb <= "000000";
					when "11011101000000110" => rgb <= "000000";
					when "11011101000000111" => rgb <= "000000";
					when "11011101000001000" => rgb <= "000000";
					when "11011101000001001" => rgb <= "000000";
					when "11011101000001010" => rgb <= "000000";
					when "11011101000001011" => rgb <= "000000";
					when "11011101000001100" => rgb <= "000000";
					when "11011101000001101" => rgb <= "000000";
					when "11011101000001110" => rgb <= "000000";
					when "11011101000001111" => rgb <= "000000";
					when "11011101000010000" => rgb <= "000000";
					when "11011101000010001" => rgb <= "000000";
					when "11011101000010010" => rgb <= "000000";
					when "11011101000010011" => rgb <= "000000";
					when "11011101000010100" => rgb <= "000000";
					when "11011101000010101" => rgb <= "000000";
					when "11011101000010110" => rgb <= "000000";
					when "11011101000010111" => rgb <= "000000";
					when "11011101000011000" => rgb <= "000000";
					when "11011101000011001" => rgb <= "000000";
					when "11011101000011010" => rgb <= "000000";
					when "11011101000011011" => rgb <= "000000";
					when "11011101000011100" => rgb <= "000000";
					when "11011101000011101" => rgb <= "000000";
					when "11011101000011110" => rgb <= "000000";
					when "11011101000011111" => rgb <= "000000";
					when "11011101000100000" => rgb <= "000000";
					when "11011101000100001" => rgb <= "000000";
					when "11011101000100010" => rgb <= "000000";
					when "11011101000100011" => rgb <= "000000";
					when "11011101000100100" => rgb <= "000000";
					when "11011101000100101" => rgb <= "000000";
					when "11011101000100110" => rgb <= "000000";
					when "11011101000100111" => rgb <= "000000";
					when "11011101000101000" => rgb <= "000000";
					when "11011101000101001" => rgb <= "000000";
					when "11011101000101010" => rgb <= "000000";
					when "11011101000101011" => rgb <= "000000";
					when "11011101000101100" => rgb <= "000000";
					when "11011101000101101" => rgb <= "000000";
					when "11011101000101110" => rgb <= "000000";
					when "11011101000101111" => rgb <= "000000";
					when "11011101000110000" => rgb <= "000000";
					when "11011101000110001" => rgb <= "000000";
					when "11011101000110010" => rgb <= "000000";
					when "11011101000110011" => rgb <= "000000";
					when "11011101000110100" => rgb <= "000000";
					when "11011101000110101" => rgb <= "000000";
					when "11011101000110110" => rgb <= "000000";
					when "11011101000110111" => rgb <= "000000";
					when "11011101000111000" => rgb <= "000000";
					when "11011101000111001" => rgb <= "000000";
					when "11011101000111010" => rgb <= "000000";
					when "11011101000111011" => rgb <= "000000";
					when "11011101000111100" => rgb <= "000000";
					when "11011101000111101" => rgb <= "000000";
					when "11011101000111110" => rgb <= "000000";
					when "11011101000111111" => rgb <= "000000";
					when "11011101001000000" => rgb <= "000000";
					when "11011101001000001" => rgb <= "000000";
					when "11011101001000010" => rgb <= "000000";
					when "11011101001000011" => rgb <= "000000";
					when "11011101001000100" => rgb <= "000000";
					when "11011101001000101" => rgb <= "000000";
					when "11011101001000110" => rgb <= "000000";
					when "11011101001000111" => rgb <= "000000";
					when "11011101001001000" => rgb <= "000000";
					when "11011101001001001" => rgb <= "000000";
					when "11011101001001010" => rgb <= "000000";
					when "11011101001001011" => rgb <= "000000";
					when "11011101001001100" => rgb <= "000000";
					when "11011101001001101" => rgb <= "000000";
					when "11011101001001110" => rgb <= "000000";
					when "11011101001001111" => rgb <= "000000";
					when "11011101001010000" => rgb <= "000000";
					when "11011101001010001" => rgb <= "000000";
					when "11011101001010010" => rgb <= "000000";
					when "11011101001010011" => rgb <= "000000";
					when "11011101001010100" => rgb <= "000000";
					when "11011101001010101" => rgb <= "000000";
					when "11011101001010110" => rgb <= "000000";
					when "11011101001010111" => rgb <= "000000";
					when "11011101001011000" => rgb <= "000000";
					when "11011101001011001" => rgb <= "000000";
					when "11011101001011010" => rgb <= "000000";
					when "11011101001011011" => rgb <= "000000";
					when "11011101001011100" => rgb <= "000000";
					when "11011101001011101" => rgb <= "000000";
					when "11011101001011110" => rgb <= "000000";
					when "11011101001011111" => rgb <= "000000";
					when "11011101001100000" => rgb <= "000000";
					when "11011101001100001" => rgb <= "000000";
					when "11011101001100010" => rgb <= "000000";
					when "11011101001100011" => rgb <= "000000";
					when "11011101001100100" => rgb <= "000000";
					when "11011101001100101" => rgb <= "000000";
					when "11011101001100110" => rgb <= "000000";
					when "11011101001100111" => rgb <= "000000";
					when "11011101001101000" => rgb <= "000000";
					when "11011101001101001" => rgb <= "000000";
					when "11011101001101010" => rgb <= "000000";
					when "11011101001101011" => rgb <= "000000";
					when "11011101001101100" => rgb <= "000000";
					when "11011101001101101" => rgb <= "000000";
					when "11011101001101110" => rgb <= "000000";
					when "11011101001101111" => rgb <= "000000";
					when "11011101001110000" => rgb <= "000000";
					when "11011101001110001" => rgb <= "000000";
					when "11011101001110010" => rgb <= "000000";
					when "11011101001110011" => rgb <= "000000";
					when "11011101001110100" => rgb <= "000000";
					when "11011101001110101" => rgb <= "000000";
					when "11011101001110110" => rgb <= "000000";
					when "11011101001110111" => rgb <= "000000";
					when "11011101001111000" => rgb <= "000000";
					when "11011101001111001" => rgb <= "000000";
					when "11011101001111010" => rgb <= "000000";
					when "11011101001111011" => rgb <= "000000";
					when "11011101001111100" => rgb <= "000000";
					when "11011101001111101" => rgb <= "000000";
					when "11011101001111110" => rgb <= "000000";
					when "11011101001111111" => rgb <= "000000";
					when "11011101010000000" => rgb <= "000000";
					when "11011101010000001" => rgb <= "000000";
					when "11011101010000010" => rgb <= "000000";
					when "11011101010000011" => rgb <= "000000";
					when "11011101010000100" => rgb <= "000000";
					when "11011101010000101" => rgb <= "000000";
					when "11011101010000110" => rgb <= "000000";
					when "11011101010000111" => rgb <= "000000";
					when "11011101010001000" => rgb <= "000000";
					when "11011101010001001" => rgb <= "000000";
					when "11011101010001010" => rgb <= "000000";
					when "11011101010001011" => rgb <= "000000";
					when "11011101010001100" => rgb <= "000000";
					when "11011101010001101" => rgb <= "000000";
					when "11011101010001110" => rgb <= "000000";
					when "11011101010001111" => rgb <= "000000";
					when "11011101010010000" => rgb <= "000000";
					when "11011101010010001" => rgb <= "000000";
					when "11011101010010010" => rgb <= "000000";
					when "11011101010010011" => rgb <= "000000";
					when "11011101010010100" => rgb <= "000000";
					when "11011101010010101" => rgb <= "000000";
					when "11011101010010110" => rgb <= "000000";
					when "11011101010010111" => rgb <= "000000";
					when "11011101010011000" => rgb <= "000000";
					when "11011101010011001" => rgb <= "000000";
					when "11011101010011010" => rgb <= "000000";
					when "11011101010011011" => rgb <= "000000";
					when "11011101010011100" => rgb <= "000000";
					when "11011101010011101" => rgb <= "000000";
					when "11011101010011110" => rgb <= "000000";
					when "11011101010011111" => rgb <= "000000";
					when "11011101010100000" => rgb <= "000000";
					when "11011101010100001" => rgb <= "000000";
					when "11011101010100010" => rgb <= "000000";
					when "11011101010100011" => rgb <= "000000";
					when "11011101010100100" => rgb <= "000000";
					when "11011101010100101" => rgb <= "000000";
					when "11011101010100110" => rgb <= "000000";
					when "11011101010100111" => rgb <= "000000";
					when "11011101010101000" => rgb <= "000000";
					when "11011101010101001" => rgb <= "000000";
					when "11011101010101010" => rgb <= "000000";
					when "11011101010101011" => rgb <= "000000";
					when "11011101010101100" => rgb <= "000000";
					when "11011101010101101" => rgb <= "000000";
					when "11011101010101110" => rgb <= "000000";
					when "11011101010101111" => rgb <= "000000";
					when "11011101010110000" => rgb <= "000000";
					when "11011101010110001" => rgb <= "000000";
					when "11011101010110010" => rgb <= "000000";
					when "11011101010110011" => rgb <= "000000";
					when "11011101010110100" => rgb <= "000000";
					when "11011101010110101" => rgb <= "000000";
					when "11011101010110110" => rgb <= "000000";
					when "11011101010110111" => rgb <= "000000";
					when "11011101010111000" => rgb <= "000000";
					when "11011101010111001" => rgb <= "000000";
					when "11011101010111010" => rgb <= "000000";
					when "11011101010111011" => rgb <= "000000";
					when "11011101010111100" => rgb <= "000000";
					when "11011101010111101" => rgb <= "000000";
					when "11011101010111110" => rgb <= "000000";
					when "11011101010111111" => rgb <= "000000";
					when "11011101011000000" => rgb <= "000000";
					when "11011101011000001" => rgb <= "000000";
					when "11011101011000010" => rgb <= "000000";
					when "11011101011000011" => rgb <= "000000";
					when "11011101011000100" => rgb <= "000000";
					when "11011101011000101" => rgb <= "000000";
					when "11011101011000110" => rgb <= "000000";
					when "11011101011000111" => rgb <= "000000";
					when "11011101011001000" => rgb <= "000000";
					when "11011101011001001" => rgb <= "000000";
					when "11011101011001010" => rgb <= "000000";
					when "11011101011001011" => rgb <= "000000";
					when "11011101011001100" => rgb <= "000000";
					when "11011101011001101" => rgb <= "000000";
					when "11011101011001110" => rgb <= "000000";
					when "11011101011001111" => rgb <= "000000";
					when "11011101011010000" => rgb <= "000000";
					when "11011101011010001" => rgb <= "000000";
					when "11011101011010010" => rgb <= "000000";
					when "11011101011010011" => rgb <= "000000";
					when "11011101011010100" => rgb <= "000000";
					when "11011101011010101" => rgb <= "000000";
					when "11011101011010110" => rgb <= "000000";
					when "11011101011010111" => rgb <= "000000";
					when "11011101011011000" => rgb <= "000000";
					when "11011101011011001" => rgb <= "000000";
					when "11011101011011010" => rgb <= "000000";
					when "11011101011011011" => rgb <= "000000";
					when "11011101011011100" => rgb <= "000000";
					when "11011101011011101" => rgb <= "000000";
					when "11011101011011110" => rgb <= "000000";
					when "11011101011011111" => rgb <= "000000";
					when "11011101011100000" => rgb <= "000000";
					when "11011101011100001" => rgb <= "000000";
					when "11011101011100010" => rgb <= "000000";
					when "11011101011100011" => rgb <= "000000";
					when "11011101011100100" => rgb <= "000000";
					when "11011101011100101" => rgb <= "000000";
					when "11011101011100110" => rgb <= "000000";
					when "11011101011100111" => rgb <= "000000";
					when "11011101011101000" => rgb <= "000000";
					when "11011101011101001" => rgb <= "000000";
					when "11011101011101010" => rgb <= "000000";
					when "11011101011101011" => rgb <= "000000";
					when "11011101011101100" => rgb <= "000000";
					when "11011101011101101" => rgb <= "000000";
					when "11011101011101110" => rgb <= "000000";
					when "11011101011101111" => rgb <= "000000";
					when "11011101011110000" => rgb <= "000000";
					when "11011101011110001" => rgb <= "000000";
					when "11011101011110010" => rgb <= "000000";
					when "11011101011110011" => rgb <= "000000";
					when "11011101011110100" => rgb <= "000000";
					when "11011101011110101" => rgb <= "000000";
					when "11011101011110110" => rgb <= "000000";
					when "11011101011110111" => rgb <= "000000";
					when "11011101011111000" => rgb <= "000000";
					when "11011101011111001" => rgb <= "000000";
					when "11011101011111010" => rgb <= "000000";
					when "11011101011111011" => rgb <= "000000";
					when "11011101011111100" => rgb <= "000000";
					when "11011101011111101" => rgb <= "000000";
					when "11011101011111110" => rgb <= "000000";
					when "11011101011111111" => rgb <= "000000";
					when "11011101100000000" => rgb <= "000000";
					when "11011101100000001" => rgb <= "000000";
					when "11011101100000010" => rgb <= "000000";
					when "11011101100000011" => rgb <= "000000";
					when "11011101100000100" => rgb <= "000000";
					when "11011101100000101" => rgb <= "000000";
					when "11011101100000110" => rgb <= "000000";
					when "11011101100000111" => rgb <= "000000";
					when "11011101100001000" => rgb <= "000000";
					when "11011101100001001" => rgb <= "000000";
					when "11011101100001010" => rgb <= "000000";
					when "11011101100001011" => rgb <= "000000";
					when "11011101100001100" => rgb <= "000000";
					when "11011101100001101" => rgb <= "000000";
					when "11011101100001110" => rgb <= "000000";
					when "11011101100001111" => rgb <= "000000";
					when "11011101100010000" => rgb <= "000000";
					when "11011101100010001" => rgb <= "000000";
					when "11011101100010010" => rgb <= "000000";
					when "11011101100010011" => rgb <= "000000";
					when "11011101100010100" => rgb <= "000000";
					when "11011101100010101" => rgb <= "000000";
					when "11011101100010110" => rgb <= "000000";
					when "11011101100010111" => rgb <= "000000";
					when "11011101100011000" => rgb <= "000000";
					when "11011101100011001" => rgb <= "000000";
					when "11011101100011010" => rgb <= "000000";
					when "11011101100011011" => rgb <= "000000";
					when "11011101100011100" => rgb <= "000000";
					when "11011101100011101" => rgb <= "000000";
					when "11011101100011110" => rgb <= "000000";
					when "11011101100011111" => rgb <= "000000";
					when "11011101100100000" => rgb <= "000000";
					when "11011101100100001" => rgb <= "000000";
					when "11011101100100010" => rgb <= "000000";
					when "11011101100100011" => rgb <= "000000";
					when "11011101100100100" => rgb <= "000000";
					when "11011101100100101" => rgb <= "000000";
					when "11011101100100110" => rgb <= "000000";
					when "11011101100100111" => rgb <= "000000";
					when "11011101100101000" => rgb <= "000000";
					when "11011101100101001" => rgb <= "000000";
					when "11011101100101010" => rgb <= "000000";
					when "11011101100101011" => rgb <= "000000";
					when "11011101100101100" => rgb <= "000000";
					when "11011101100101101" => rgb <= "000000";
					when "11011101100101110" => rgb <= "000000";
					when "11011101100101111" => rgb <= "000000";
					when "11011101100110000" => rgb <= "000000";
					when "11011101100110001" => rgb <= "000000";
					when "11011101100110010" => rgb <= "000000";
					when "11011101100110011" => rgb <= "000000";
					when "11011101100110100" => rgb <= "000000";
					when "11011101100110101" => rgb <= "000000";
					when "11011101100110110" => rgb <= "000000";
					when "11011101100110111" => rgb <= "000000";
					when "11011101100111000" => rgb <= "000000";
					when "11011101100111001" => rgb <= "000000";
					when "11011101100111010" => rgb <= "000000";
					when "11011101100111011" => rgb <= "000000";
					when "11011101100111100" => rgb <= "000000";
					when "11011101100111101" => rgb <= "000000";
					when "11011101100111110" => rgb <= "000000";
					when "11011101100111111" => rgb <= "000000";
					when "11011110000000000" => rgb <= "000000";
					when "11011110000000001" => rgb <= "000000";
					when "11011110000000010" => rgb <= "000000";
					when "11011110000000011" => rgb <= "000000";
					when "11011110000000100" => rgb <= "000000";
					when "11011110000000101" => rgb <= "000000";
					when "11011110000000110" => rgb <= "000000";
					when "11011110000000111" => rgb <= "000000";
					when "11011110000001000" => rgb <= "000000";
					when "11011110000001001" => rgb <= "000000";
					when "11011110000001010" => rgb <= "000000";
					when "11011110000001011" => rgb <= "000000";
					when "11011110000001100" => rgb <= "000000";
					when "11011110000001101" => rgb <= "000000";
					when "11011110000001110" => rgb <= "000000";
					when "11011110000001111" => rgb <= "000000";
					when "11011110000010000" => rgb <= "000000";
					when "11011110000010001" => rgb <= "000000";
					when "11011110000010010" => rgb <= "000000";
					when "11011110000010011" => rgb <= "000000";
					when "11011110000010100" => rgb <= "000000";
					when "11011110000010101" => rgb <= "000000";
					when "11011110000010110" => rgb <= "000000";
					when "11011110000010111" => rgb <= "000000";
					when "11011110000011000" => rgb <= "000000";
					when "11011110000011001" => rgb <= "000000";
					when "11011110000011010" => rgb <= "000000";
					when "11011110000011011" => rgb <= "000000";
					when "11011110000011100" => rgb <= "000000";
					when "11011110000011101" => rgb <= "000000";
					when "11011110000011110" => rgb <= "000000";
					when "11011110000011111" => rgb <= "000000";
					when "11011110000100000" => rgb <= "000000";
					when "11011110000100001" => rgb <= "000000";
					when "11011110000100010" => rgb <= "000000";
					when "11011110000100011" => rgb <= "000000";
					when "11011110000100100" => rgb <= "000000";
					when "11011110000100101" => rgb <= "000000";
					when "11011110000100110" => rgb <= "000000";
					when "11011110000100111" => rgb <= "000000";
					when "11011110000101000" => rgb <= "000000";
					when "11011110000101001" => rgb <= "000000";
					when "11011110000101010" => rgb <= "000000";
					when "11011110000101011" => rgb <= "000000";
					when "11011110000101100" => rgb <= "000000";
					when "11011110000101101" => rgb <= "000000";
					when "11011110000101110" => rgb <= "000000";
					when "11011110000101111" => rgb <= "000000";
					when "11011110000110000" => rgb <= "000000";
					when "11011110000110001" => rgb <= "000000";
					when "11011110000110010" => rgb <= "000000";
					when "11011110000110011" => rgb <= "000000";
					when "11011110000110100" => rgb <= "000000";
					when "11011110000110101" => rgb <= "000000";
					when "11011110000110110" => rgb <= "000000";
					when "11011110000110111" => rgb <= "000000";
					when "11011110000111000" => rgb <= "000000";
					when "11011110000111001" => rgb <= "000000";
					when "11011110000111010" => rgb <= "000000";
					when "11011110000111011" => rgb <= "000000";
					when "11011110000111100" => rgb <= "000000";
					when "11011110000111101" => rgb <= "000000";
					when "11011110000111110" => rgb <= "000000";
					when "11011110000111111" => rgb <= "000000";
					when "11011110001000000" => rgb <= "000000";
					when "11011110001000001" => rgb <= "000000";
					when "11011110001000010" => rgb <= "000000";
					when "11011110001000011" => rgb <= "000000";
					when "11011110001000100" => rgb <= "000000";
					when "11011110001000101" => rgb <= "000000";
					when "11011110001000110" => rgb <= "000000";
					when "11011110001000111" => rgb <= "000000";
					when "11011110001001000" => rgb <= "000000";
					when "11011110001001001" => rgb <= "000000";
					when "11011110001001010" => rgb <= "000000";
					when "11011110001001011" => rgb <= "000000";
					when "11011110001001100" => rgb <= "000000";
					when "11011110001001101" => rgb <= "000000";
					when "11011110001001110" => rgb <= "000000";
					when "11011110001001111" => rgb <= "000000";
					when "11011110001010000" => rgb <= "000000";
					when "11011110001010001" => rgb <= "000000";
					when "11011110001010010" => rgb <= "000000";
					when "11011110001010011" => rgb <= "000000";
					when "11011110001010100" => rgb <= "000000";
					when "11011110001010101" => rgb <= "000000";
					when "11011110001010110" => rgb <= "000000";
					when "11011110001010111" => rgb <= "000000";
					when "11011110001011000" => rgb <= "000000";
					when "11011110001011001" => rgb <= "000000";
					when "11011110001011010" => rgb <= "000000";
					when "11011110001011011" => rgb <= "000000";
					when "11011110001011100" => rgb <= "000000";
					when "11011110001011101" => rgb <= "000000";
					when "11011110001011110" => rgb <= "000000";
					when "11011110001011111" => rgb <= "000000";
					when "11011110001100000" => rgb <= "000000";
					when "11011110001100001" => rgb <= "000000";
					when "11011110001100010" => rgb <= "000000";
					when "11011110001100011" => rgb <= "000000";
					when "11011110001100100" => rgb <= "000000";
					when "11011110001100101" => rgb <= "000000";
					when "11011110001100110" => rgb <= "000000";
					when "11011110001100111" => rgb <= "000000";
					when "11011110001101000" => rgb <= "000000";
					when "11011110001101001" => rgb <= "000000";
					when "11011110001101010" => rgb <= "000000";
					when "11011110001101011" => rgb <= "000000";
					when "11011110001101100" => rgb <= "000000";
					when "11011110001101101" => rgb <= "000000";
					when "11011110001101110" => rgb <= "000000";
					when "11011110001101111" => rgb <= "000000";
					when "11011110001110000" => rgb <= "000000";
					when "11011110001110001" => rgb <= "000000";
					when "11011110001110010" => rgb <= "000000";
					when "11011110001110011" => rgb <= "000000";
					when "11011110001110100" => rgb <= "000000";
					when "11011110001110101" => rgb <= "000000";
					when "11011110001110110" => rgb <= "000000";
					when "11011110001110111" => rgb <= "000000";
					when "11011110001111000" => rgb <= "000000";
					when "11011110001111001" => rgb <= "000000";
					when "11011110001111010" => rgb <= "000000";
					when "11011110001111011" => rgb <= "000000";
					when "11011110001111100" => rgb <= "000000";
					when "11011110001111101" => rgb <= "000000";
					when "11011110001111110" => rgb <= "000000";
					when "11011110001111111" => rgb <= "000000";
					when "11011110010000000" => rgb <= "000000";
					when "11011110010000001" => rgb <= "000000";
					when "11011110010000010" => rgb <= "000000";
					when "11011110010000011" => rgb <= "000000";
					when "11011110010000100" => rgb <= "000000";
					when "11011110010000101" => rgb <= "000000";
					when "11011110010000110" => rgb <= "000000";
					when "11011110010000111" => rgb <= "000000";
					when "11011110010001000" => rgb <= "000000";
					when "11011110010001001" => rgb <= "000000";
					when "11011110010001010" => rgb <= "000000";
					when "11011110010001011" => rgb <= "000000";
					when "11011110010001100" => rgb <= "000000";
					when "11011110010001101" => rgb <= "000000";
					when "11011110010001110" => rgb <= "000000";
					when "11011110010001111" => rgb <= "000000";
					when "11011110010010000" => rgb <= "000000";
					when "11011110010010001" => rgb <= "000000";
					when "11011110010010010" => rgb <= "000000";
					when "11011110010010011" => rgb <= "000000";
					when "11011110010010100" => rgb <= "000000";
					when "11011110010010101" => rgb <= "000000";
					when "11011110010010110" => rgb <= "000000";
					when "11011110010010111" => rgb <= "000000";
					when "11011110010011000" => rgb <= "000000";
					when "11011110010011001" => rgb <= "000000";
					when "11011110010011010" => rgb <= "000000";
					when "11011110010011011" => rgb <= "000000";
					when "11011110010011100" => rgb <= "000000";
					when "11011110010011101" => rgb <= "000000";
					when "11011110010011110" => rgb <= "000000";
					when "11011110010011111" => rgb <= "000000";
					when "11011110010100000" => rgb <= "000000";
					when "11011110010100001" => rgb <= "000000";
					when "11011110010100010" => rgb <= "000000";
					when "11011110010100011" => rgb <= "000000";
					when "11011110010100100" => rgb <= "000000";
					when "11011110010100101" => rgb <= "000000";
					when "11011110010100110" => rgb <= "000000";
					when "11011110010100111" => rgb <= "000000";
					when "11011110010101000" => rgb <= "000000";
					when "11011110010101001" => rgb <= "000000";
					when "11011110010101010" => rgb <= "000000";
					when "11011110010101011" => rgb <= "000000";
					when "11011110010101100" => rgb <= "000000";
					when "11011110010101101" => rgb <= "000000";
					when "11011110010101110" => rgb <= "000000";
					when "11011110010101111" => rgb <= "000000";
					when "11011110010110000" => rgb <= "000000";
					when "11011110010110001" => rgb <= "000000";
					when "11011110010110010" => rgb <= "000000";
					when "11011110010110011" => rgb <= "000000";
					when "11011110010110100" => rgb <= "000000";
					when "11011110010110101" => rgb <= "000000";
					when "11011110010110110" => rgb <= "000000";
					when "11011110010110111" => rgb <= "000000";
					when "11011110010111000" => rgb <= "000000";
					when "11011110010111001" => rgb <= "000000";
					when "11011110010111010" => rgb <= "000000";
					when "11011110010111011" => rgb <= "000000";
					when "11011110010111100" => rgb <= "000000";
					when "11011110010111101" => rgb <= "000000";
					when "11011110010111110" => rgb <= "000000";
					when "11011110010111111" => rgb <= "000000";
					when "11011110011000000" => rgb <= "000000";
					when "11011110011000001" => rgb <= "000000";
					when "11011110011000010" => rgb <= "000000";
					when "11011110011000011" => rgb <= "000000";
					when "11011110011000100" => rgb <= "000000";
					when "11011110011000101" => rgb <= "000000";
					when "11011110011000110" => rgb <= "000000";
					when "11011110011000111" => rgb <= "000000";
					when "11011110011001000" => rgb <= "000000";
					when "11011110011001001" => rgb <= "000000";
					when "11011110011001010" => rgb <= "000000";
					when "11011110011001011" => rgb <= "000000";
					when "11011110011001100" => rgb <= "000000";
					when "11011110011001101" => rgb <= "000000";
					when "11011110011001110" => rgb <= "000000";
					when "11011110011001111" => rgb <= "000000";
					when "11011110011010000" => rgb <= "000000";
					when "11011110011010001" => rgb <= "000000";
					when "11011110011010010" => rgb <= "000000";
					when "11011110011010011" => rgb <= "000000";
					when "11011110011010100" => rgb <= "000000";
					when "11011110011010101" => rgb <= "000000";
					when "11011110011010110" => rgb <= "000000";
					when "11011110011010111" => rgb <= "000000";
					when "11011110011011000" => rgb <= "000000";
					when "11011110011011001" => rgb <= "000000";
					when "11011110011011010" => rgb <= "000000";
					when "11011110011011011" => rgb <= "000000";
					when "11011110011011100" => rgb <= "000000";
					when "11011110011011101" => rgb <= "000000";
					when "11011110011011110" => rgb <= "000000";
					when "11011110011011111" => rgb <= "000000";
					when "11011110011100000" => rgb <= "000000";
					when "11011110011100001" => rgb <= "000000";
					when "11011110011100010" => rgb <= "000000";
					when "11011110011100011" => rgb <= "000000";
					when "11011110011100100" => rgb <= "000000";
					when "11011110011100101" => rgb <= "000000";
					when "11011110011100110" => rgb <= "000000";
					when "11011110011100111" => rgb <= "000000";
					when "11011110011101000" => rgb <= "000000";
					when "11011110011101001" => rgb <= "000000";
					when "11011110011101010" => rgb <= "000000";
					when "11011110011101011" => rgb <= "000000";
					when "11011110011101100" => rgb <= "000000";
					when "11011110011101101" => rgb <= "000000";
					when "11011110011101110" => rgb <= "000000";
					when "11011110011101111" => rgb <= "000000";
					when "11011110011110000" => rgb <= "000000";
					when "11011110011110001" => rgb <= "000000";
					when "11011110011110010" => rgb <= "000000";
					when "11011110011110011" => rgb <= "000000";
					when "11011110011110100" => rgb <= "000000";
					when "11011110011110101" => rgb <= "000000";
					when "11011110011110110" => rgb <= "000000";
					when "11011110011110111" => rgb <= "000000";
					when "11011110011111000" => rgb <= "000000";
					when "11011110011111001" => rgb <= "000000";
					when "11011110011111010" => rgb <= "000000";
					when "11011110011111011" => rgb <= "000000";
					when "11011110011111100" => rgb <= "000000";
					when "11011110011111101" => rgb <= "000000";
					when "11011110011111110" => rgb <= "000000";
					when "11011110011111111" => rgb <= "000000";
					when "11011110100000000" => rgb <= "000000";
					when "11011110100000001" => rgb <= "000000";
					when "11011110100000010" => rgb <= "000000";
					when "11011110100000011" => rgb <= "000000";
					when "11011110100000100" => rgb <= "000000";
					when "11011110100000101" => rgb <= "000000";
					when "11011110100000110" => rgb <= "000000";
					when "11011110100000111" => rgb <= "000000";
					when "11011110100001000" => rgb <= "000000";
					when "11011110100001001" => rgb <= "000000";
					when "11011110100001010" => rgb <= "000000";
					when "11011110100001011" => rgb <= "000000";
					when "11011110100001100" => rgb <= "000000";
					when "11011110100001101" => rgb <= "000000";
					when "11011110100001110" => rgb <= "000000";
					when "11011110100001111" => rgb <= "000000";
					when "11011110100010000" => rgb <= "000000";
					when "11011110100010001" => rgb <= "000000";
					when "11011110100010010" => rgb <= "000000";
					when "11011110100010011" => rgb <= "000000";
					when "11011110100010100" => rgb <= "000000";
					when "11011110100010101" => rgb <= "000000";
					when "11011110100010110" => rgb <= "000000";
					when "11011110100010111" => rgb <= "000000";
					when "11011110100011000" => rgb <= "000000";
					when "11011110100011001" => rgb <= "000000";
					when "11011110100011010" => rgb <= "000000";
					when "11011110100011011" => rgb <= "000000";
					when "11011110100011100" => rgb <= "000000";
					when "11011110100011101" => rgb <= "000000";
					when "11011110100011110" => rgb <= "000000";
					when "11011110100011111" => rgb <= "000000";
					when "11011110100100000" => rgb <= "000000";
					when "11011110100100001" => rgb <= "000000";
					when "11011110100100010" => rgb <= "000000";
					when "11011110100100011" => rgb <= "000000";
					when "11011110100100100" => rgb <= "000000";
					when "11011110100100101" => rgb <= "000000";
					when "11011110100100110" => rgb <= "000000";
					when "11011110100100111" => rgb <= "000000";
					when "11011110100101000" => rgb <= "000000";
					when "11011110100101001" => rgb <= "000000";
					when "11011110100101010" => rgb <= "000000";
					when "11011110100101011" => rgb <= "000000";
					when "11011110100101100" => rgb <= "000000";
					when "11011110100101101" => rgb <= "000000";
					when "11011110100101110" => rgb <= "000000";
					when "11011110100101111" => rgb <= "000000";
					when "11011110100110000" => rgb <= "000000";
					when "11011110100110001" => rgb <= "000000";
					when "11011110100110010" => rgb <= "000000";
					when "11011110100110011" => rgb <= "000000";
					when "11011110100110100" => rgb <= "000000";
					when "11011110100110101" => rgb <= "000000";
					when "11011110100110110" => rgb <= "000000";
					when "11011110100110111" => rgb <= "000000";
					when "11011110100111000" => rgb <= "000000";
					when "11011110100111001" => rgb <= "000000";
					when "11011110100111010" => rgb <= "000000";
					when "11011110100111011" => rgb <= "000000";
					when "11011110100111100" => rgb <= "000000";
					when "11011110100111101" => rgb <= "000000";
					when "11011110100111110" => rgb <= "000000";
					when "11011110100111111" => rgb <= "000000";
					when "11011111000000000" => rgb <= "000000";
					when "11011111000000001" => rgb <= "000000";
					when "11011111000000010" => rgb <= "000000";
					when "11011111000000011" => rgb <= "000000";
					when "11011111000000100" => rgb <= "000000";
					when "11011111000000101" => rgb <= "000000";
					when "11011111000000110" => rgb <= "000000";
					when "11011111000000111" => rgb <= "000000";
					when "11011111000001000" => rgb <= "000000";
					when "11011111000001001" => rgb <= "000000";
					when "11011111000001010" => rgb <= "000000";
					when "11011111000001011" => rgb <= "000000";
					when "11011111000001100" => rgb <= "000000";
					when "11011111000001101" => rgb <= "000000";
					when "11011111000001110" => rgb <= "000000";
					when "11011111000001111" => rgb <= "000000";
					when "11011111000010000" => rgb <= "000000";
					when "11011111000010001" => rgb <= "000000";
					when "11011111000010010" => rgb <= "000000";
					when "11011111000010011" => rgb <= "000000";
					when "11011111000010100" => rgb <= "000000";
					when "11011111000010101" => rgb <= "000000";
					when "11011111000010110" => rgb <= "000000";
					when "11011111000010111" => rgb <= "000000";
					when "11011111000011000" => rgb <= "000000";
					when "11011111000011001" => rgb <= "000000";
					when "11011111000011010" => rgb <= "000000";
					when "11011111000011011" => rgb <= "000000";
					when "11011111000011100" => rgb <= "000000";
					when "11011111000011101" => rgb <= "000000";
					when "11011111000011110" => rgb <= "000000";
					when "11011111000011111" => rgb <= "000000";
					when "11011111000100000" => rgb <= "000000";
					when "11011111000100001" => rgb <= "000000";
					when "11011111000100010" => rgb <= "000000";
					when "11011111000100011" => rgb <= "000000";
					when "11011111000100100" => rgb <= "000000";
					when "11011111000100101" => rgb <= "000000";
					when "11011111000100110" => rgb <= "000000";
					when "11011111000100111" => rgb <= "000000";
					when "11011111000101000" => rgb <= "000000";
					when "11011111000101001" => rgb <= "000000";
					when "11011111000101010" => rgb <= "000000";
					when "11011111000101011" => rgb <= "000000";
					when "11011111000101100" => rgb <= "000000";
					when "11011111000101101" => rgb <= "000000";
					when "11011111000101110" => rgb <= "000000";
					when "11011111000101111" => rgb <= "000000";
					when "11011111000110000" => rgb <= "000000";
					when "11011111000110001" => rgb <= "000000";
					when "11011111000110010" => rgb <= "000000";
					when "11011111000110011" => rgb <= "000000";
					when "11011111000110100" => rgb <= "000000";
					when "11011111000110101" => rgb <= "000000";
					when "11011111000110110" => rgb <= "000000";
					when "11011111000110111" => rgb <= "000000";
					when "11011111000111000" => rgb <= "000000";
					when "11011111000111001" => rgb <= "000000";
					when "11011111000111010" => rgb <= "000000";
					when "11011111000111011" => rgb <= "000000";
					when "11011111000111100" => rgb <= "000000";
					when "11011111000111101" => rgb <= "000000";
					when "11011111000111110" => rgb <= "000000";
					when "11011111000111111" => rgb <= "000000";
					when "11011111001000000" => rgb <= "000000";
					when "11011111001000001" => rgb <= "000000";
					when "11011111001000010" => rgb <= "000000";
					when "11011111001000011" => rgb <= "000000";
					when "11011111001000100" => rgb <= "000000";
					when "11011111001000101" => rgb <= "000000";
					when "11011111001000110" => rgb <= "000000";
					when "11011111001000111" => rgb <= "000000";
					when "11011111001001000" => rgb <= "000000";
					when "11011111001001001" => rgb <= "000000";
					when "11011111001001010" => rgb <= "000000";
					when "11011111001001011" => rgb <= "000000";
					when "11011111001001100" => rgb <= "000000";
					when "11011111001001101" => rgb <= "000000";
					when "11011111001001110" => rgb <= "000000";
					when "11011111001001111" => rgb <= "000000";
					when "11011111001010000" => rgb <= "000000";
					when "11011111001010001" => rgb <= "000000";
					when "11011111001010010" => rgb <= "000000";
					when "11011111001010011" => rgb <= "000000";
					when "11011111001010100" => rgb <= "000000";
					when "11011111001010101" => rgb <= "000000";
					when "11011111001010110" => rgb <= "000000";
					when "11011111001010111" => rgb <= "000000";
					when "11011111001011000" => rgb <= "000000";
					when "11011111001011001" => rgb <= "000000";
					when "11011111001011010" => rgb <= "000000";
					when "11011111001011011" => rgb <= "000000";
					when "11011111001011100" => rgb <= "000000";
					when "11011111001011101" => rgb <= "000000";
					when "11011111001011110" => rgb <= "000000";
					when "11011111001011111" => rgb <= "000000";
					when "11011111001100000" => rgb <= "000000";
					when "11011111001100001" => rgb <= "000000";
					when "11011111001100010" => rgb <= "000000";
					when "11011111001100011" => rgb <= "000000";
					when "11011111001100100" => rgb <= "000000";
					when "11011111001100101" => rgb <= "000000";
					when "11011111001100110" => rgb <= "000000";
					when "11011111001100111" => rgb <= "000000";
					when "11011111001101000" => rgb <= "000000";
					when "11011111001101001" => rgb <= "000000";
					when "11011111001101010" => rgb <= "000000";
					when "11011111001101011" => rgb <= "000000";
					when "11011111001101100" => rgb <= "000000";
					when "11011111001101101" => rgb <= "000000";
					when "11011111001101110" => rgb <= "000000";
					when "11011111001101111" => rgb <= "000000";
					when "11011111001110000" => rgb <= "000000";
					when "11011111001110001" => rgb <= "000000";
					when "11011111001110010" => rgb <= "000000";
					when "11011111001110011" => rgb <= "000000";
					when "11011111001110100" => rgb <= "000000";
					when "11011111001110101" => rgb <= "000000";
					when "11011111001110110" => rgb <= "000000";
					when "11011111001110111" => rgb <= "000000";
					when "11011111001111000" => rgb <= "000000";
					when "11011111001111001" => rgb <= "000000";
					when "11011111001111010" => rgb <= "000000";
					when "11011111001111011" => rgb <= "000000";
					when "11011111001111100" => rgb <= "000000";
					when "11011111001111101" => rgb <= "000000";
					when "11011111001111110" => rgb <= "000000";
					when "11011111001111111" => rgb <= "000000";
					when "11011111010000000" => rgb <= "000000";
					when "11011111010000001" => rgb <= "000000";
					when "11011111010000010" => rgb <= "000000";
					when "11011111010000011" => rgb <= "000000";
					when "11011111010000100" => rgb <= "000000";
					when "11011111010000101" => rgb <= "000000";
					when "11011111010000110" => rgb <= "000000";
					when "11011111010000111" => rgb <= "000000";
					when "11011111010001000" => rgb <= "000000";
					when "11011111010001001" => rgb <= "000000";
					when "11011111010001010" => rgb <= "000000";
					when "11011111010001011" => rgb <= "000000";
					when "11011111010001100" => rgb <= "000000";
					when "11011111010001101" => rgb <= "000000";
					when "11011111010001110" => rgb <= "000000";
					when "11011111010001111" => rgb <= "000000";
					when "11011111010010000" => rgb <= "000000";
					when "11011111010010001" => rgb <= "000000";
					when "11011111010010010" => rgb <= "000000";
					when "11011111010010011" => rgb <= "000000";
					when "11011111010010100" => rgb <= "000000";
					when "11011111010010101" => rgb <= "000000";
					when "11011111010010110" => rgb <= "000000";
					when "11011111010010111" => rgb <= "000000";
					when "11011111010011000" => rgb <= "000000";
					when "11011111010011001" => rgb <= "000000";
					when "11011111010011010" => rgb <= "000000";
					when "11011111010011011" => rgb <= "000000";
					when "11011111010011100" => rgb <= "000000";
					when "11011111010011101" => rgb <= "000000";
					when "11011111010011110" => rgb <= "000000";
					when "11011111010011111" => rgb <= "000000";
					when "11011111010100000" => rgb <= "000000";
					when "11011111010100001" => rgb <= "000000";
					when "11011111010100010" => rgb <= "000000";
					when "11011111010100011" => rgb <= "000000";
					when "11011111010100100" => rgb <= "000000";
					when "11011111010100101" => rgb <= "000000";
					when "11011111010100110" => rgb <= "000000";
					when "11011111010100111" => rgb <= "000000";
					when "11011111010101000" => rgb <= "000000";
					when "11011111010101001" => rgb <= "000000";
					when "11011111010101010" => rgb <= "000000";
					when "11011111010101011" => rgb <= "000000";
					when "11011111010101100" => rgb <= "000000";
					when "11011111010101101" => rgb <= "000000";
					when "11011111010101110" => rgb <= "000000";
					when "11011111010101111" => rgb <= "000000";
					when "11011111010110000" => rgb <= "000000";
					when "11011111010110001" => rgb <= "000000";
					when "11011111010110010" => rgb <= "000000";
					when "11011111010110011" => rgb <= "000000";
					when "11011111010110100" => rgb <= "000000";
					when "11011111010110101" => rgb <= "000000";
					when "11011111010110110" => rgb <= "000000";
					when "11011111010110111" => rgb <= "000000";
					when "11011111010111000" => rgb <= "000000";
					when "11011111010111001" => rgb <= "000000";
					when "11011111010111010" => rgb <= "000000";
					when "11011111010111011" => rgb <= "000000";
					when "11011111010111100" => rgb <= "000000";
					when "11011111010111101" => rgb <= "000000";
					when "11011111010111110" => rgb <= "000000";
					when "11011111010111111" => rgb <= "000000";
					when "11011111011000000" => rgb <= "000000";
					when "11011111011000001" => rgb <= "000000";
					when "11011111011000010" => rgb <= "000000";
					when "11011111011000011" => rgb <= "000000";
					when "11011111011000100" => rgb <= "000000";
					when "11011111011000101" => rgb <= "000000";
					when "11011111011000110" => rgb <= "000000";
					when "11011111011000111" => rgb <= "000000";
					when "11011111011001000" => rgb <= "000000";
					when "11011111011001001" => rgb <= "000000";
					when "11011111011001010" => rgb <= "000000";
					when "11011111011001011" => rgb <= "000000";
					when "11011111011001100" => rgb <= "000000";
					when "11011111011001101" => rgb <= "000000";
					when "11011111011001110" => rgb <= "000000";
					when "11011111011001111" => rgb <= "000000";
					when "11011111011010000" => rgb <= "000000";
					when "11011111011010001" => rgb <= "000000";
					when "11011111011010010" => rgb <= "000000";
					when "11011111011010011" => rgb <= "000000";
					when "11011111011010100" => rgb <= "000000";
					when "11011111011010101" => rgb <= "000000";
					when "11011111011010110" => rgb <= "000000";
					when "11011111011010111" => rgb <= "000000";
					when "11011111011011000" => rgb <= "000000";
					when "11011111011011001" => rgb <= "000000";
					when "11011111011011010" => rgb <= "000000";
					when "11011111011011011" => rgb <= "000000";
					when "11011111011011100" => rgb <= "000000";
					when "11011111011011101" => rgb <= "000000";
					when "11011111011011110" => rgb <= "000000";
					when "11011111011011111" => rgb <= "000000";
					when "11011111011100000" => rgb <= "000000";
					when "11011111011100001" => rgb <= "000000";
					when "11011111011100010" => rgb <= "000000";
					when "11011111011100011" => rgb <= "000000";
					when "11011111011100100" => rgb <= "000000";
					when "11011111011100101" => rgb <= "000000";
					when "11011111011100110" => rgb <= "000000";
					when "11011111011100111" => rgb <= "000000";
					when "11011111011101000" => rgb <= "000000";
					when "11011111011101001" => rgb <= "000000";
					when "11011111011101010" => rgb <= "000000";
					when "11011111011101011" => rgb <= "000000";
					when "11011111011101100" => rgb <= "000000";
					when "11011111011101101" => rgb <= "000000";
					when "11011111011101110" => rgb <= "000000";
					when "11011111011101111" => rgb <= "000000";
					when "11011111011110000" => rgb <= "000000";
					when "11011111011110001" => rgb <= "000000";
					when "11011111011110010" => rgb <= "000000";
					when "11011111011110011" => rgb <= "000000";
					when "11011111011110100" => rgb <= "000000";
					when "11011111011110101" => rgb <= "000000";
					when "11011111011110110" => rgb <= "000000";
					when "11011111011110111" => rgb <= "000000";
					when "11011111011111000" => rgb <= "000000";
					when "11011111011111001" => rgb <= "000000";
					when "11011111011111010" => rgb <= "000000";
					when "11011111011111011" => rgb <= "000000";
					when "11011111011111100" => rgb <= "000000";
					when "11011111011111101" => rgb <= "000000";
					when "11011111011111110" => rgb <= "000000";
					when "11011111011111111" => rgb <= "000000";
					when "11011111100000000" => rgb <= "000000";
					when "11011111100000001" => rgb <= "000000";
					when "11011111100000010" => rgb <= "000000";
					when "11011111100000011" => rgb <= "000000";
					when "11011111100000100" => rgb <= "000000";
					when "11011111100000101" => rgb <= "000000";
					when "11011111100000110" => rgb <= "000000";
					when "11011111100000111" => rgb <= "000000";
					when "11011111100001000" => rgb <= "000000";
					when "11011111100001001" => rgb <= "000000";
					when "11011111100001010" => rgb <= "000000";
					when "11011111100001011" => rgb <= "000000";
					when "11011111100001100" => rgb <= "000000";
					when "11011111100001101" => rgb <= "000000";
					when "11011111100001110" => rgb <= "000000";
					when "11011111100001111" => rgb <= "000000";
					when "11011111100010000" => rgb <= "000000";
					when "11011111100010001" => rgb <= "000000";
					when "11011111100010010" => rgb <= "000000";
					when "11011111100010011" => rgb <= "000000";
					when "11011111100010100" => rgb <= "000000";
					when "11011111100010101" => rgb <= "000000";
					when "11011111100010110" => rgb <= "000000";
					when "11011111100010111" => rgb <= "000000";
					when "11011111100011000" => rgb <= "000000";
					when "11011111100011001" => rgb <= "000000";
					when "11011111100011010" => rgb <= "000000";
					when "11011111100011011" => rgb <= "000000";
					when "11011111100011100" => rgb <= "000000";
					when "11011111100011101" => rgb <= "000000";
					when "11011111100011110" => rgb <= "000000";
					when "11011111100011111" => rgb <= "000000";
					when "11011111100100000" => rgb <= "000000";
					when "11011111100100001" => rgb <= "000000";
					when "11011111100100010" => rgb <= "000000";
					when "11011111100100011" => rgb <= "000000";
					when "11011111100100100" => rgb <= "000000";
					when "11011111100100101" => rgb <= "000000";
					when "11011111100100110" => rgb <= "000000";
					when "11011111100100111" => rgb <= "000000";
					when "11011111100101000" => rgb <= "000000";
					when "11011111100101001" => rgb <= "000000";
					when "11011111100101010" => rgb <= "000000";
					when "11011111100101011" => rgb <= "000000";
					when "11011111100101100" => rgb <= "000000";
					when "11011111100101101" => rgb <= "000000";
					when "11011111100101110" => rgb <= "000000";
					when "11011111100101111" => rgb <= "000000";
					when "11011111100110000" => rgb <= "000000";
					when "11011111100110001" => rgb <= "000000";
					when "11011111100110010" => rgb <= "000000";
					when "11011111100110011" => rgb <= "000000";
					when "11011111100110100" => rgb <= "000000";
					when "11011111100110101" => rgb <= "000000";
					when "11011111100110110" => rgb <= "000000";
					when "11011111100110111" => rgb <= "000000";
					when "11011111100111000" => rgb <= "000000";
					when "11011111100111001" => rgb <= "000000";
					when "11011111100111010" => rgb <= "000000";
					when "11011111100111011" => rgb <= "000000";
					when "11011111100111100" => rgb <= "000000";
					when "11011111100111101" => rgb <= "000000";
					when "11011111100111110" => rgb <= "000000";
					when "11011111100111111" => rgb <= "000000";
					when "11100000000000000" => rgb <= "000000";
					when "11100000000000001" => rgb <= "000000";
					when "11100000000000010" => rgb <= "000000";
					when "11100000000000011" => rgb <= "000000";
					when "11100000000000100" => rgb <= "000000";
					when "11100000000000101" => rgb <= "000000";
					when "11100000000000110" => rgb <= "000000";
					when "11100000000000111" => rgb <= "000000";
					when "11100000000001000" => rgb <= "000000";
					when "11100000000001001" => rgb <= "000000";
					when "11100000000001010" => rgb <= "000000";
					when "11100000000001011" => rgb <= "000000";
					when "11100000000001100" => rgb <= "000000";
					when "11100000000001101" => rgb <= "000000";
					when "11100000000001110" => rgb <= "000000";
					when "11100000000001111" => rgb <= "000000";
					when "11100000000010000" => rgb <= "000000";
					when "11100000000010001" => rgb <= "000000";
					when "11100000000010010" => rgb <= "000000";
					when "11100000000010011" => rgb <= "000000";
					when "11100000000010100" => rgb <= "000000";
					when "11100000000010101" => rgb <= "000000";
					when "11100000000010110" => rgb <= "000000";
					when "11100000000010111" => rgb <= "000000";
					when "11100000000011000" => rgb <= "000000";
					when "11100000000011001" => rgb <= "000000";
					when "11100000000011010" => rgb <= "000000";
					when "11100000000011011" => rgb <= "000000";
					when "11100000000011100" => rgb <= "000000";
					when "11100000000011101" => rgb <= "000000";
					when "11100000000011110" => rgb <= "000000";
					when "11100000000011111" => rgb <= "000000";
					when "11100000000100000" => rgb <= "000000";
					when "11100000000100001" => rgb <= "000000";
					when "11100000000100010" => rgb <= "000000";
					when "11100000000100011" => rgb <= "000000";
					when "11100000000100100" => rgb <= "000000";
					when "11100000000100101" => rgb <= "000000";
					when "11100000000100110" => rgb <= "000000";
					when "11100000000100111" => rgb <= "000000";
					when "11100000000101000" => rgb <= "000000";
					when "11100000000101001" => rgb <= "000000";
					when "11100000000101010" => rgb <= "000000";
					when "11100000000101011" => rgb <= "000000";
					when "11100000000101100" => rgb <= "000000";
					when "11100000000101101" => rgb <= "000000";
					when "11100000000101110" => rgb <= "000000";
					when "11100000000101111" => rgb <= "000000";
					when "11100000000110000" => rgb <= "000000";
					when "11100000000110001" => rgb <= "000000";
					when "11100000000110010" => rgb <= "000000";
					when "11100000000110011" => rgb <= "000000";
					when "11100000000110100" => rgb <= "000000";
					when "11100000000110101" => rgb <= "000000";
					when "11100000000110110" => rgb <= "000000";
					when "11100000000110111" => rgb <= "000000";
					when "11100000000111000" => rgb <= "000000";
					when "11100000000111001" => rgb <= "000000";
					when "11100000000111010" => rgb <= "000000";
					when "11100000000111011" => rgb <= "000000";
					when "11100000000111100" => rgb <= "000000";
					when "11100000000111101" => rgb <= "000000";
					when "11100000000111110" => rgb <= "000000";
					when "11100000000111111" => rgb <= "000000";
					when "11100000001000000" => rgb <= "000000";
					when "11100000001000001" => rgb <= "000000";
					when "11100000001000010" => rgb <= "000000";
					when "11100000001000011" => rgb <= "000000";
					when "11100000001000100" => rgb <= "000000";
					when "11100000001000101" => rgb <= "000000";
					when "11100000001000110" => rgb <= "000000";
					when "11100000001000111" => rgb <= "000000";
					when "11100000001001000" => rgb <= "000000";
					when "11100000001001001" => rgb <= "000000";
					when "11100000001001010" => rgb <= "000000";
					when "11100000001001011" => rgb <= "000000";
					when "11100000001001100" => rgb <= "000000";
					when "11100000001001101" => rgb <= "000000";
					when "11100000001001110" => rgb <= "000000";
					when "11100000001001111" => rgb <= "000000";
					when "11100000001010000" => rgb <= "000000";
					when "11100000001010001" => rgb <= "000000";
					when "11100000001010010" => rgb <= "000000";
					when "11100000001010011" => rgb <= "000000";
					when "11100000001010100" => rgb <= "000000";
					when "11100000001010101" => rgb <= "000000";
					when "11100000001010110" => rgb <= "000000";
					when "11100000001010111" => rgb <= "000000";
					when "11100000001011000" => rgb <= "000000";
					when "11100000001011001" => rgb <= "000000";
					when "11100000001011010" => rgb <= "000000";
					when "11100000001011011" => rgb <= "000000";
					when "11100000001011100" => rgb <= "000000";
					when "11100000001011101" => rgb <= "000000";
					when "11100000001011110" => rgb <= "000000";
					when "11100000001011111" => rgb <= "000000";
					when "11100000001100000" => rgb <= "000000";
					when "11100000001100001" => rgb <= "000000";
					when "11100000001100010" => rgb <= "000000";
					when "11100000001100011" => rgb <= "000000";
					when "11100000001100100" => rgb <= "000000";
					when "11100000001100101" => rgb <= "000000";
					when "11100000001100110" => rgb <= "000000";
					when "11100000001100111" => rgb <= "000000";
					when "11100000001101000" => rgb <= "000000";
					when "11100000001101001" => rgb <= "000000";
					when "11100000001101010" => rgb <= "000000";
					when "11100000001101011" => rgb <= "000000";
					when "11100000001101100" => rgb <= "000000";
					when "11100000001101101" => rgb <= "000000";
					when "11100000001101110" => rgb <= "000000";
					when "11100000001101111" => rgb <= "000000";
					when "11100000001110000" => rgb <= "000000";
					when "11100000001110001" => rgb <= "000000";
					when "11100000001110010" => rgb <= "000000";
					when "11100000001110011" => rgb <= "000000";
					when "11100000001110100" => rgb <= "000000";
					when "11100000001110101" => rgb <= "000000";
					when "11100000001110110" => rgb <= "000000";
					when "11100000001110111" => rgb <= "000000";
					when "11100000001111000" => rgb <= "000000";
					when "11100000001111001" => rgb <= "000000";
					when "11100000001111010" => rgb <= "000000";
					when "11100000001111011" => rgb <= "000000";
					when "11100000001111100" => rgb <= "000000";
					when "11100000001111101" => rgb <= "000000";
					when "11100000001111110" => rgb <= "000000";
					when "11100000001111111" => rgb <= "000000";
					when "11100000010000000" => rgb <= "000000";
					when "11100000010000001" => rgb <= "000000";
					when "11100000010000010" => rgb <= "000000";
					when "11100000010000011" => rgb <= "000000";
					when "11100000010000100" => rgb <= "000000";
					when "11100000010000101" => rgb <= "000000";
					when "11100000010000110" => rgb <= "000000";
					when "11100000010000111" => rgb <= "000000";
					when "11100000010001000" => rgb <= "000000";
					when "11100000010001001" => rgb <= "000000";
					when "11100000010001010" => rgb <= "000000";
					when "11100000010001011" => rgb <= "000000";
					when "11100000010001100" => rgb <= "000000";
					when "11100000010001101" => rgb <= "000000";
					when "11100000010001110" => rgb <= "000000";
					when "11100000010001111" => rgb <= "000000";
					when "11100000010010000" => rgb <= "000000";
					when "11100000010010001" => rgb <= "000000";
					when "11100000010010010" => rgb <= "000000";
					when "11100000010010011" => rgb <= "000000";
					when "11100000010010100" => rgb <= "000000";
					when "11100000010010101" => rgb <= "000000";
					when "11100000010010110" => rgb <= "000000";
					when "11100000010010111" => rgb <= "000000";
					when "11100000010011000" => rgb <= "000000";
					when "11100000010011001" => rgb <= "000000";
					when "11100000010011010" => rgb <= "000000";
					when "11100000010011011" => rgb <= "000000";
					when "11100000010011100" => rgb <= "000000";
					when "11100000010011101" => rgb <= "000000";
					when "11100000010011110" => rgb <= "000000";
					when "11100000010011111" => rgb <= "000000";
					when "11100000010100000" => rgb <= "000000";
					when "11100000010100001" => rgb <= "000000";
					when "11100000010100010" => rgb <= "000000";
					when "11100000010100011" => rgb <= "000000";
					when "11100000010100100" => rgb <= "000000";
					when "11100000010100101" => rgb <= "000000";
					when "11100000010100110" => rgb <= "000000";
					when "11100000010100111" => rgb <= "000000";
					when "11100000010101000" => rgb <= "000000";
					when "11100000010101001" => rgb <= "000000";
					when "11100000010101010" => rgb <= "000000";
					when "11100000010101011" => rgb <= "000000";
					when "11100000010101100" => rgb <= "000000";
					when "11100000010101101" => rgb <= "000000";
					when "11100000010101110" => rgb <= "000000";
					when "11100000010101111" => rgb <= "000000";
					when "11100000010110000" => rgb <= "000000";
					when "11100000010110001" => rgb <= "000000";
					when "11100000010110010" => rgb <= "000000";
					when "11100000010110011" => rgb <= "000000";
					when "11100000010110100" => rgb <= "000000";
					when "11100000010110101" => rgb <= "000000";
					when "11100000010110110" => rgb <= "000000";
					when "11100000010110111" => rgb <= "000000";
					when "11100000010111000" => rgb <= "000000";
					when "11100000010111001" => rgb <= "000000";
					when "11100000010111010" => rgb <= "000000";
					when "11100000010111011" => rgb <= "000000";
					when "11100000010111100" => rgb <= "000000";
					when "11100000010111101" => rgb <= "000000";
					when "11100000010111110" => rgb <= "000000";
					when "11100000010111111" => rgb <= "000000";
					when "11100000011000000" => rgb <= "000000";
					when "11100000011000001" => rgb <= "000000";
					when "11100000011000010" => rgb <= "000000";
					when "11100000011000011" => rgb <= "000000";
					when "11100000011000100" => rgb <= "000000";
					when "11100000011000101" => rgb <= "000000";
					when "11100000011000110" => rgb <= "000000";
					when "11100000011000111" => rgb <= "000000";
					when "11100000011001000" => rgb <= "000000";
					when "11100000011001001" => rgb <= "000000";
					when "11100000011001010" => rgb <= "000000";
					when "11100000011001011" => rgb <= "000000";
					when "11100000011001100" => rgb <= "000000";
					when "11100000011001101" => rgb <= "000000";
					when "11100000011001110" => rgb <= "000000";
					when "11100000011001111" => rgb <= "000000";
					when "11100000011010000" => rgb <= "000000";
					when "11100000011010001" => rgb <= "000000";
					when "11100000011010010" => rgb <= "000000";
					when "11100000011010011" => rgb <= "000000";
					when "11100000011010100" => rgb <= "000000";
					when "11100000011010101" => rgb <= "000000";
					when "11100000011010110" => rgb <= "000000";
					when "11100000011010111" => rgb <= "000000";
					when "11100000011011000" => rgb <= "000000";
					when "11100000011011001" => rgb <= "000000";
					when "11100000011011010" => rgb <= "000000";
					when "11100000011011011" => rgb <= "000000";
					when "11100000011011100" => rgb <= "000000";
					when "11100000011011101" => rgb <= "000000";
					when "11100000011011110" => rgb <= "000000";
					when "11100000011011111" => rgb <= "000000";
					when "11100000011100000" => rgb <= "000000";
					when "11100000011100001" => rgb <= "000000";
					when "11100000011100010" => rgb <= "000000";
					when "11100000011100011" => rgb <= "000000";
					when "11100000011100100" => rgb <= "000000";
					when "11100000011100101" => rgb <= "000000";
					when "11100000011100110" => rgb <= "000000";
					when "11100000011100111" => rgb <= "000000";
					when "11100000011101000" => rgb <= "000000";
					when "11100000011101001" => rgb <= "000000";
					when "11100000011101010" => rgb <= "000000";
					when "11100000011101011" => rgb <= "000000";
					when "11100000011101100" => rgb <= "000000";
					when "11100000011101101" => rgb <= "000000";
					when "11100000011101110" => rgb <= "000000";
					when "11100000011101111" => rgb <= "000000";
					when "11100000011110000" => rgb <= "000000";
					when "11100000011110001" => rgb <= "000000";
					when "11100000011110010" => rgb <= "000000";
					when "11100000011110011" => rgb <= "000000";
					when "11100000011110100" => rgb <= "000000";
					when "11100000011110101" => rgb <= "000000";
					when "11100000011110110" => rgb <= "000000";
					when "11100000011110111" => rgb <= "000000";
					when "11100000011111000" => rgb <= "000000";
					when "11100000011111001" => rgb <= "000000";
					when "11100000011111010" => rgb <= "000000";
					when "11100000011111011" => rgb <= "000000";
					when "11100000011111100" => rgb <= "000000";
					when "11100000011111101" => rgb <= "000000";
					when "11100000011111110" => rgb <= "000000";
					when "11100000011111111" => rgb <= "000000";
					when "11100000100000000" => rgb <= "000000";
					when "11100000100000001" => rgb <= "000000";
					when "11100000100000010" => rgb <= "000000";
					when "11100000100000011" => rgb <= "000000";
					when "11100000100000100" => rgb <= "000000";
					when "11100000100000101" => rgb <= "000000";
					when "11100000100000110" => rgb <= "000000";
					when "11100000100000111" => rgb <= "000000";
					when "11100000100001000" => rgb <= "000000";
					when "11100000100001001" => rgb <= "000000";
					when "11100000100001010" => rgb <= "000000";
					when "11100000100001011" => rgb <= "000000";
					when "11100000100001100" => rgb <= "000000";
					when "11100000100001101" => rgb <= "000000";
					when "11100000100001110" => rgb <= "000000";
					when "11100000100001111" => rgb <= "000000";
					when "11100000100010000" => rgb <= "000000";
					when "11100000100010001" => rgb <= "000000";
					when "11100000100010010" => rgb <= "000000";
					when "11100000100010011" => rgb <= "000000";
					when "11100000100010100" => rgb <= "000000";
					when "11100000100010101" => rgb <= "000000";
					when "11100000100010110" => rgb <= "000000";
					when "11100000100010111" => rgb <= "000000";
					when "11100000100011000" => rgb <= "000000";
					when "11100000100011001" => rgb <= "000000";
					when "11100000100011010" => rgb <= "000000";
					when "11100000100011011" => rgb <= "000000";
					when "11100000100011100" => rgb <= "000000";
					when "11100000100011101" => rgb <= "000000";
					when "11100000100011110" => rgb <= "000000";
					when "11100000100011111" => rgb <= "000000";
					when "11100000100100000" => rgb <= "000000";
					when "11100000100100001" => rgb <= "000000";
					when "11100000100100010" => rgb <= "000000";
					when "11100000100100011" => rgb <= "000000";
					when "11100000100100100" => rgb <= "000000";
					when "11100000100100101" => rgb <= "000000";
					when "11100000100100110" => rgb <= "000000";
					when "11100000100100111" => rgb <= "000000";
					when "11100000100101000" => rgb <= "000000";
					when "11100000100101001" => rgb <= "000000";
					when "11100000100101010" => rgb <= "000000";
					when "11100000100101011" => rgb <= "000000";
					when "11100000100101100" => rgb <= "000000";
					when "11100000100101101" => rgb <= "000000";
					when "11100000100101110" => rgb <= "000000";
					when "11100000100101111" => rgb <= "000000";
					when "11100000100110000" => rgb <= "000000";
					when "11100000100110001" => rgb <= "000000";
					when "11100000100110010" => rgb <= "000000";
					when "11100000100110011" => rgb <= "000000";
					when "11100000100110100" => rgb <= "000000";
					when "11100000100110101" => rgb <= "000000";
					when "11100000100110110" => rgb <= "000000";
					when "11100000100110111" => rgb <= "000000";
					when "11100000100111000" => rgb <= "000000";
					when "11100000100111001" => rgb <= "000000";
					when "11100000100111010" => rgb <= "000000";
					when "11100000100111011" => rgb <= "000000";
					when "11100000100111100" => rgb <= "000000";
					when "11100000100111101" => rgb <= "000000";
					when "11100000100111110" => rgb <= "000000";
					when "11100000100111111" => rgb <= "000000";
					when "11100001000000000" => rgb <= "000000";
					when "11100001000000001" => rgb <= "000000";
					when "11100001000000010" => rgb <= "000000";
					when "11100001000000011" => rgb <= "000000";
					when "11100001000000100" => rgb <= "000000";
					when "11100001000000101" => rgb <= "000000";
					when "11100001000000110" => rgb <= "000000";
					when "11100001000000111" => rgb <= "000000";
					when "11100001000001000" => rgb <= "000000";
					when "11100001000001001" => rgb <= "000000";
					when "11100001000001010" => rgb <= "000000";
					when "11100001000001011" => rgb <= "000000";
					when "11100001000001100" => rgb <= "000000";
					when "11100001000001101" => rgb <= "000000";
					when "11100001000001110" => rgb <= "000000";
					when "11100001000001111" => rgb <= "000000";
					when "11100001000010000" => rgb <= "000000";
					when "11100001000010001" => rgb <= "000000";
					when "11100001000010010" => rgb <= "000000";
					when "11100001000010011" => rgb <= "000000";
					when "11100001000010100" => rgb <= "000000";
					when "11100001000010101" => rgb <= "000000";
					when "11100001000010110" => rgb <= "000000";
					when "11100001000010111" => rgb <= "000000";
					when "11100001000011000" => rgb <= "000000";
					when "11100001000011001" => rgb <= "000000";
					when "11100001000011010" => rgb <= "000000";
					when "11100001000011011" => rgb <= "000000";
					when "11100001000011100" => rgb <= "000000";
					when "11100001000011101" => rgb <= "000000";
					when "11100001000011110" => rgb <= "000000";
					when "11100001000011111" => rgb <= "000000";
					when "11100001000100000" => rgb <= "000000";
					when "11100001000100001" => rgb <= "000000";
					when "11100001000100010" => rgb <= "000000";
					when "11100001000100011" => rgb <= "000000";
					when "11100001000100100" => rgb <= "000000";
					when "11100001000100101" => rgb <= "000000";
					when "11100001000100110" => rgb <= "000000";
					when "11100001000100111" => rgb <= "000000";
					when "11100001000101000" => rgb <= "000000";
					when "11100001000101001" => rgb <= "000000";
					when "11100001000101010" => rgb <= "000000";
					when "11100001000101011" => rgb <= "000000";
					when "11100001000101100" => rgb <= "000000";
					when "11100001000101101" => rgb <= "000000";
					when "11100001000101110" => rgb <= "000000";
					when "11100001000101111" => rgb <= "000000";
					when "11100001000110000" => rgb <= "000000";
					when "11100001000110001" => rgb <= "000000";
					when "11100001000110010" => rgb <= "000000";
					when "11100001000110011" => rgb <= "000000";
					when "11100001000110100" => rgb <= "000000";
					when "11100001000110101" => rgb <= "000000";
					when "11100001000110110" => rgb <= "000000";
					when "11100001000110111" => rgb <= "000000";
					when "11100001000111000" => rgb <= "000000";
					when "11100001000111001" => rgb <= "000000";
					when "11100001000111010" => rgb <= "000000";
					when "11100001000111011" => rgb <= "000000";
					when "11100001000111100" => rgb <= "000000";
					when "11100001000111101" => rgb <= "000000";
					when "11100001000111110" => rgb <= "000000";
					when "11100001000111111" => rgb <= "000000";
					when "11100001001000000" => rgb <= "000000";
					when "11100001001000001" => rgb <= "000000";
					when "11100001001000010" => rgb <= "000000";
					when "11100001001000011" => rgb <= "000000";
					when "11100001001000100" => rgb <= "000000";
					when "11100001001000101" => rgb <= "000000";
					when "11100001001000110" => rgb <= "000000";
					when "11100001001000111" => rgb <= "000000";
					when "11100001001001000" => rgb <= "000000";
					when "11100001001001001" => rgb <= "000000";
					when "11100001001001010" => rgb <= "000000";
					when "11100001001001011" => rgb <= "000000";
					when "11100001001001100" => rgb <= "000000";
					when "11100001001001101" => rgb <= "000000";
					when "11100001001001110" => rgb <= "000000";
					when "11100001001001111" => rgb <= "000000";
					when "11100001001010000" => rgb <= "000000";
					when "11100001001010001" => rgb <= "000000";
					when "11100001001010010" => rgb <= "000000";
					when "11100001001010011" => rgb <= "000000";
					when "11100001001010100" => rgb <= "000000";
					when "11100001001010101" => rgb <= "000000";
					when "11100001001010110" => rgb <= "000000";
					when "11100001001010111" => rgb <= "000000";
					when "11100001001011000" => rgb <= "000000";
					when "11100001001011001" => rgb <= "000000";
					when "11100001001011010" => rgb <= "000000";
					when "11100001001011011" => rgb <= "000000";
					when "11100001001011100" => rgb <= "000000";
					when "11100001001011101" => rgb <= "000000";
					when "11100001001011110" => rgb <= "000000";
					when "11100001001011111" => rgb <= "000000";
					when "11100001001100000" => rgb <= "000000";
					when "11100001001100001" => rgb <= "000000";
					when "11100001001100010" => rgb <= "000000";
					when "11100001001100011" => rgb <= "000000";
					when "11100001001100100" => rgb <= "000000";
					when "11100001001100101" => rgb <= "000000";
					when "11100001001100110" => rgb <= "000000";
					when "11100001001100111" => rgb <= "000000";
					when "11100001001101000" => rgb <= "000000";
					when "11100001001101001" => rgb <= "000000";
					when "11100001001101010" => rgb <= "000000";
					when "11100001001101011" => rgb <= "000000";
					when "11100001001101100" => rgb <= "000000";
					when "11100001001101101" => rgb <= "000000";
					when "11100001001101110" => rgb <= "000000";
					when "11100001001101111" => rgb <= "000000";
					when "11100001001110000" => rgb <= "000000";
					when "11100001001110001" => rgb <= "000000";
					when "11100001001110010" => rgb <= "000000";
					when "11100001001110011" => rgb <= "000000";
					when "11100001001110100" => rgb <= "000000";
					when "11100001001110101" => rgb <= "000000";
					when "11100001001110110" => rgb <= "000000";
					when "11100001001110111" => rgb <= "000000";
					when "11100001001111000" => rgb <= "000000";
					when "11100001001111001" => rgb <= "000000";
					when "11100001001111010" => rgb <= "000000";
					when "11100001001111011" => rgb <= "000000";
					when "11100001001111100" => rgb <= "000000";
					when "11100001001111101" => rgb <= "000000";
					when "11100001001111110" => rgb <= "000000";
					when "11100001001111111" => rgb <= "000000";
					when "11100001010000000" => rgb <= "000000";
					when "11100001010000001" => rgb <= "000000";
					when "11100001010000010" => rgb <= "000000";
					when "11100001010000011" => rgb <= "000000";
					when "11100001010000100" => rgb <= "000000";
					when "11100001010000101" => rgb <= "000000";
					when "11100001010000110" => rgb <= "000000";
					when "11100001010000111" => rgb <= "000000";
					when "11100001010001000" => rgb <= "000000";
					when "11100001010001001" => rgb <= "000000";
					when "11100001010001010" => rgb <= "000000";
					when "11100001010001011" => rgb <= "000000";
					when "11100001010001100" => rgb <= "000000";
					when "11100001010001101" => rgb <= "000000";
					when "11100001010001110" => rgb <= "000000";
					when "11100001010001111" => rgb <= "000000";
					when "11100001010010000" => rgb <= "000000";
					when "11100001010010001" => rgb <= "000000";
					when "11100001010010010" => rgb <= "000000";
					when "11100001010010011" => rgb <= "000000";
					when "11100001010010100" => rgb <= "000000";
					when "11100001010010101" => rgb <= "000000";
					when "11100001010010110" => rgb <= "000000";
					when "11100001010010111" => rgb <= "000000";
					when "11100001010011000" => rgb <= "000000";
					when "11100001010011001" => rgb <= "000000";
					when "11100001010011010" => rgb <= "000000";
					when "11100001010011011" => rgb <= "000000";
					when "11100001010011100" => rgb <= "000000";
					when "11100001010011101" => rgb <= "000000";
					when "11100001010011110" => rgb <= "000000";
					when "11100001010011111" => rgb <= "000000";
					when "11100001010100000" => rgb <= "000000";
					when "11100001010100001" => rgb <= "000000";
					when "11100001010100010" => rgb <= "000000";
					when "11100001010100011" => rgb <= "000000";
					when "11100001010100100" => rgb <= "000000";
					when "11100001010100101" => rgb <= "000000";
					when "11100001010100110" => rgb <= "000000";
					when "11100001010100111" => rgb <= "000000";
					when "11100001010101000" => rgb <= "000000";
					when "11100001010101001" => rgb <= "000000";
					when "11100001010101010" => rgb <= "000000";
					when "11100001010101011" => rgb <= "000000";
					when "11100001010101100" => rgb <= "000000";
					when "11100001010101101" => rgb <= "000000";
					when "11100001010101110" => rgb <= "000000";
					when "11100001010101111" => rgb <= "000000";
					when "11100001010110000" => rgb <= "000000";
					when "11100001010110001" => rgb <= "000000";
					when "11100001010110010" => rgb <= "000000";
					when "11100001010110011" => rgb <= "000000";
					when "11100001010110100" => rgb <= "000000";
					when "11100001010110101" => rgb <= "000000";
					when "11100001010110110" => rgb <= "000000";
					when "11100001010110111" => rgb <= "000000";
					when "11100001010111000" => rgb <= "000000";
					when "11100001010111001" => rgb <= "000000";
					when "11100001010111010" => rgb <= "000000";
					when "11100001010111011" => rgb <= "000000";
					when "11100001010111100" => rgb <= "000000";
					when "11100001010111101" => rgb <= "000000";
					when "11100001010111110" => rgb <= "000000";
					when "11100001010111111" => rgb <= "000000";
					when "11100001011000000" => rgb <= "000000";
					when "11100001011000001" => rgb <= "000000";
					when "11100001011000010" => rgb <= "000000";
					when "11100001011000011" => rgb <= "000000";
					when "11100001011000100" => rgb <= "000000";
					when "11100001011000101" => rgb <= "000000";
					when "11100001011000110" => rgb <= "000000";
					when "11100001011000111" => rgb <= "000000";
					when "11100001011001000" => rgb <= "000000";
					when "11100001011001001" => rgb <= "000000";
					when "11100001011001010" => rgb <= "000000";
					when "11100001011001011" => rgb <= "000000";
					when "11100001011001100" => rgb <= "000000";
					when "11100001011001101" => rgb <= "000000";
					when "11100001011001110" => rgb <= "000000";
					when "11100001011001111" => rgb <= "000000";
					when "11100001011010000" => rgb <= "000000";
					when "11100001011010001" => rgb <= "000000";
					when "11100001011010010" => rgb <= "000000";
					when "11100001011010011" => rgb <= "000000";
					when "11100001011010100" => rgb <= "000000";
					when "11100001011010101" => rgb <= "000000";
					when "11100001011010110" => rgb <= "000000";
					when "11100001011010111" => rgb <= "000000";
					when "11100001011011000" => rgb <= "000000";
					when "11100001011011001" => rgb <= "000000";
					when "11100001011011010" => rgb <= "000000";
					when "11100001011011011" => rgb <= "000000";
					when "11100001011011100" => rgb <= "000000";
					when "11100001011011101" => rgb <= "000000";
					when "11100001011011110" => rgb <= "000000";
					when "11100001011011111" => rgb <= "000000";
					when "11100001011100000" => rgb <= "000000";
					when "11100001011100001" => rgb <= "000000";
					when "11100001011100010" => rgb <= "000000";
					when "11100001011100011" => rgb <= "000000";
					when "11100001011100100" => rgb <= "000000";
					when "11100001011100101" => rgb <= "000000";
					when "11100001011100110" => rgb <= "000000";
					when "11100001011100111" => rgb <= "000000";
					when "11100001011101000" => rgb <= "000000";
					when "11100001011101001" => rgb <= "000000";
					when "11100001011101010" => rgb <= "000000";
					when "11100001011101011" => rgb <= "000000";
					when "11100001011101100" => rgb <= "000000";
					when "11100001011101101" => rgb <= "000000";
					when "11100001011101110" => rgb <= "000000";
					when "11100001011101111" => rgb <= "000000";
					when "11100001011110000" => rgb <= "000000";
					when "11100001011110001" => rgb <= "000000";
					when "11100001011110010" => rgb <= "000000";
					when "11100001011110011" => rgb <= "000000";
					when "11100001011110100" => rgb <= "000000";
					when "11100001011110101" => rgb <= "000000";
					when "11100001011110110" => rgb <= "000000";
					when "11100001011110111" => rgb <= "000000";
					when "11100001011111000" => rgb <= "000000";
					when "11100001011111001" => rgb <= "000000";
					when "11100001011111010" => rgb <= "000000";
					when "11100001011111011" => rgb <= "000000";
					when "11100001011111100" => rgb <= "000000";
					when "11100001011111101" => rgb <= "000000";
					when "11100001011111110" => rgb <= "000000";
					when "11100001011111111" => rgb <= "000000";
					when "11100001100000000" => rgb <= "000000";
					when "11100001100000001" => rgb <= "000000";
					when "11100001100000010" => rgb <= "000000";
					when "11100001100000011" => rgb <= "000000";
					when "11100001100000100" => rgb <= "000000";
					when "11100001100000101" => rgb <= "000000";
					when "11100001100000110" => rgb <= "000000";
					when "11100001100000111" => rgb <= "000000";
					when "11100001100001000" => rgb <= "000000";
					when "11100001100001001" => rgb <= "000000";
					when "11100001100001010" => rgb <= "000000";
					when "11100001100001011" => rgb <= "000000";
					when "11100001100001100" => rgb <= "000000";
					when "11100001100001101" => rgb <= "000000";
					when "11100001100001110" => rgb <= "000000";
					when "11100001100001111" => rgb <= "000000";
					when "11100001100010000" => rgb <= "000000";
					when "11100001100010001" => rgb <= "000000";
					when "11100001100010010" => rgb <= "000000";
					when "11100001100010011" => rgb <= "000000";
					when "11100001100010100" => rgb <= "000000";
					when "11100001100010101" => rgb <= "000000";
					when "11100001100010110" => rgb <= "000000";
					when "11100001100010111" => rgb <= "000000";
					when "11100001100011000" => rgb <= "000000";
					when "11100001100011001" => rgb <= "000000";
					when "11100001100011010" => rgb <= "000000";
					when "11100001100011011" => rgb <= "000000";
					when "11100001100011100" => rgb <= "000000";
					when "11100001100011101" => rgb <= "000000";
					when "11100001100011110" => rgb <= "000000";
					when "11100001100011111" => rgb <= "000000";
					when "11100001100100000" => rgb <= "000000";
					when "11100001100100001" => rgb <= "000000";
					when "11100001100100010" => rgb <= "000000";
					when "11100001100100011" => rgb <= "000000";
					when "11100001100100100" => rgb <= "000000";
					when "11100001100100101" => rgb <= "000000";
					when "11100001100100110" => rgb <= "000000";
					when "11100001100100111" => rgb <= "000000";
					when "11100001100101000" => rgb <= "000000";
					when "11100001100101001" => rgb <= "000000";
					when "11100001100101010" => rgb <= "000000";
					when "11100001100101011" => rgb <= "000000";
					when "11100001100101100" => rgb <= "000000";
					when "11100001100101101" => rgb <= "000000";
					when "11100001100101110" => rgb <= "000000";
					when "11100001100101111" => rgb <= "000000";
					when "11100001100110000" => rgb <= "000000";
					when "11100001100110001" => rgb <= "000000";
					when "11100001100110010" => rgb <= "000000";
					when "11100001100110011" => rgb <= "000000";
					when "11100001100110100" => rgb <= "000000";
					when "11100001100110101" => rgb <= "000000";
					when "11100001100110110" => rgb <= "000000";
					when "11100001100110111" => rgb <= "000000";
					when "11100001100111000" => rgb <= "000000";
					when "11100001100111001" => rgb <= "000000";
					when "11100001100111010" => rgb <= "000000";
					when "11100001100111011" => rgb <= "000000";
					when "11100001100111100" => rgb <= "000000";
					when "11100001100111101" => rgb <= "000000";
					when "11100001100111110" => rgb <= "000000";
					when "11100001100111111" => rgb <= "000000";
					when "11100010000000000" => rgb <= "000000";
					when "11100010000000001" => rgb <= "000000";
					when "11100010000000010" => rgb <= "000000";
					when "11100010000000011" => rgb <= "000000";
					when "11100010000000100" => rgb <= "000000";
					when "11100010000000101" => rgb <= "000000";
					when "11100010000000110" => rgb <= "000000";
					when "11100010000000111" => rgb <= "000000";
					when "11100010000001000" => rgb <= "000000";
					when "11100010000001001" => rgb <= "000000";
					when "11100010000001010" => rgb <= "000000";
					when "11100010000001011" => rgb <= "000000";
					when "11100010000001100" => rgb <= "000000";
					when "11100010000001101" => rgb <= "000000";
					when "11100010000001110" => rgb <= "000000";
					when "11100010000001111" => rgb <= "000000";
					when "11100010000010000" => rgb <= "000000";
					when "11100010000010001" => rgb <= "000000";
					when "11100010000010010" => rgb <= "000000";
					when "11100010000010011" => rgb <= "000000";
					when "11100010000010100" => rgb <= "000000";
					when "11100010000010101" => rgb <= "000000";
					when "11100010000010110" => rgb <= "000000";
					when "11100010000010111" => rgb <= "000000";
					when "11100010000011000" => rgb <= "000000";
					when "11100010000011001" => rgb <= "000000";
					when "11100010000011010" => rgb <= "000000";
					when "11100010000011011" => rgb <= "000000";
					when "11100010000011100" => rgb <= "000000";
					when "11100010000011101" => rgb <= "000000";
					when "11100010000011110" => rgb <= "000000";
					when "11100010000011111" => rgb <= "000000";
					when "11100010000100000" => rgb <= "000000";
					when "11100010000100001" => rgb <= "000000";
					when "11100010000100010" => rgb <= "000000";
					when "11100010000100011" => rgb <= "000000";
					when "11100010000100100" => rgb <= "000000";
					when "11100010000100101" => rgb <= "000000";
					when "11100010000100110" => rgb <= "000000";
					when "11100010000100111" => rgb <= "000000";
					when "11100010000101000" => rgb <= "000000";
					when "11100010000101001" => rgb <= "000000";
					when "11100010000101010" => rgb <= "000000";
					when "11100010000101011" => rgb <= "000000";
					when "11100010000101100" => rgb <= "000000";
					when "11100010000101101" => rgb <= "000000";
					when "11100010000101110" => rgb <= "000000";
					when "11100010000101111" => rgb <= "000000";
					when "11100010000110000" => rgb <= "000000";
					when "11100010000110001" => rgb <= "000000";
					when "11100010000110010" => rgb <= "000000";
					when "11100010000110011" => rgb <= "000000";
					when "11100010000110100" => rgb <= "000000";
					when "11100010000110101" => rgb <= "000000";
					when "11100010000110110" => rgb <= "000000";
					when "11100010000110111" => rgb <= "000000";
					when "11100010000111000" => rgb <= "000000";
					when "11100010000111001" => rgb <= "000000";
					when "11100010000111010" => rgb <= "000000";
					when "11100010000111011" => rgb <= "000000";
					when "11100010000111100" => rgb <= "000000";
					when "11100010000111101" => rgb <= "000000";
					when "11100010000111110" => rgb <= "000000";
					when "11100010000111111" => rgb <= "000000";
					when "11100010001000000" => rgb <= "000000";
					when "11100010001000001" => rgb <= "000000";
					when "11100010001000010" => rgb <= "000000";
					when "11100010001000011" => rgb <= "000000";
					when "11100010001000100" => rgb <= "000000";
					when "11100010001000101" => rgb <= "000000";
					when "11100010001000110" => rgb <= "000000";
					when "11100010001000111" => rgb <= "000000";
					when "11100010001001000" => rgb <= "000000";
					when "11100010001001001" => rgb <= "000000";
					when "11100010001001010" => rgb <= "000000";
					when "11100010001001011" => rgb <= "000000";
					when "11100010001001100" => rgb <= "000000";
					when "11100010001001101" => rgb <= "000000";
					when "11100010001001110" => rgb <= "000000";
					when "11100010001001111" => rgb <= "000000";
					when "11100010001010000" => rgb <= "000000";
					when "11100010001010001" => rgb <= "000000";
					when "11100010001010010" => rgb <= "000000";
					when "11100010001010011" => rgb <= "000000";
					when "11100010001010100" => rgb <= "000000";
					when "11100010001010101" => rgb <= "000000";
					when "11100010001010110" => rgb <= "000000";
					when "11100010001010111" => rgb <= "000000";
					when "11100010001011000" => rgb <= "000000";
					when "11100010001011001" => rgb <= "000000";
					when "11100010001011010" => rgb <= "000000";
					when "11100010001011011" => rgb <= "000000";
					when "11100010001011100" => rgb <= "000000";
					when "11100010001011101" => rgb <= "000000";
					when "11100010001011110" => rgb <= "000000";
					when "11100010001011111" => rgb <= "000000";
					when "11100010001100000" => rgb <= "000000";
					when "11100010001100001" => rgb <= "000000";
					when "11100010001100010" => rgb <= "000000";
					when "11100010001100011" => rgb <= "000000";
					when "11100010001100100" => rgb <= "000000";
					when "11100010001100101" => rgb <= "000000";
					when "11100010001100110" => rgb <= "000000";
					when "11100010001100111" => rgb <= "000000";
					when "11100010001101000" => rgb <= "000000";
					when "11100010001101001" => rgb <= "000000";
					when "11100010001101010" => rgb <= "000000";
					when "11100010001101011" => rgb <= "000000";
					when "11100010001101100" => rgb <= "000000";
					when "11100010001101101" => rgb <= "000000";
					when "11100010001101110" => rgb <= "000000";
					when "11100010001101111" => rgb <= "000000";
					when "11100010001110000" => rgb <= "000000";
					when "11100010001110001" => rgb <= "000000";
					when "11100010001110010" => rgb <= "000000";
					when "11100010001110011" => rgb <= "000000";
					when "11100010001110100" => rgb <= "000000";
					when "11100010001110101" => rgb <= "000000";
					when "11100010001110110" => rgb <= "000000";
					when "11100010001110111" => rgb <= "000000";
					when "11100010001111000" => rgb <= "000000";
					when "11100010001111001" => rgb <= "000000";
					when "11100010001111010" => rgb <= "000000";
					when "11100010001111011" => rgb <= "000000";
					when "11100010001111100" => rgb <= "000000";
					when "11100010001111101" => rgb <= "000000";
					when "11100010001111110" => rgb <= "000000";
					when "11100010001111111" => rgb <= "000000";
					when "11100010010000000" => rgb <= "000000";
					when "11100010010000001" => rgb <= "000000";
					when "11100010010000010" => rgb <= "000000";
					when "11100010010000011" => rgb <= "000000";
					when "11100010010000100" => rgb <= "000000";
					when "11100010010000101" => rgb <= "000000";
					when "11100010010000110" => rgb <= "000000";
					when "11100010010000111" => rgb <= "000000";
					when "11100010010001000" => rgb <= "000000";
					when "11100010010001001" => rgb <= "000000";
					when "11100010010001010" => rgb <= "000000";
					when "11100010010001011" => rgb <= "000000";
					when "11100010010001100" => rgb <= "000000";
					when "11100010010001101" => rgb <= "000000";
					when "11100010010001110" => rgb <= "000000";
					when "11100010010001111" => rgb <= "000000";
					when "11100010010010000" => rgb <= "000000";
					when "11100010010010001" => rgb <= "000000";
					when "11100010010010010" => rgb <= "000000";
					when "11100010010010011" => rgb <= "000000";
					when "11100010010010100" => rgb <= "000000";
					when "11100010010010101" => rgb <= "000000";
					when "11100010010010110" => rgb <= "000000";
					when "11100010010010111" => rgb <= "000000";
					when "11100010010011000" => rgb <= "000000";
					when "11100010010011001" => rgb <= "000000";
					when "11100010010011010" => rgb <= "000000";
					when "11100010010011011" => rgb <= "000000";
					when "11100010010011100" => rgb <= "000000";
					when "11100010010011101" => rgb <= "000000";
					when "11100010010011110" => rgb <= "000000";
					when "11100010010011111" => rgb <= "000000";
					when "11100010010100000" => rgb <= "000000";
					when "11100010010100001" => rgb <= "000000";
					when "11100010010100010" => rgb <= "000000";
					when "11100010010100011" => rgb <= "000000";
					when "11100010010100100" => rgb <= "000000";
					when "11100010010100101" => rgb <= "000000";
					when "11100010010100110" => rgb <= "000000";
					when "11100010010100111" => rgb <= "000000";
					when "11100010010101000" => rgb <= "000000";
					when "11100010010101001" => rgb <= "000000";
					when "11100010010101010" => rgb <= "000000";
					when "11100010010101011" => rgb <= "000000";
					when "11100010010101100" => rgb <= "000000";
					when "11100010010101101" => rgb <= "000000";
					when "11100010010101110" => rgb <= "000000";
					when "11100010010101111" => rgb <= "000000";
					when "11100010010110000" => rgb <= "000000";
					when "11100010010110001" => rgb <= "000000";
					when "11100010010110010" => rgb <= "000000";
					when "11100010010110011" => rgb <= "000000";
					when "11100010010110100" => rgb <= "000000";
					when "11100010010110101" => rgb <= "000000";
					when "11100010010110110" => rgb <= "000000";
					when "11100010010110111" => rgb <= "000000";
					when "11100010010111000" => rgb <= "000000";
					when "11100010010111001" => rgb <= "000000";
					when "11100010010111010" => rgb <= "000000";
					when "11100010010111011" => rgb <= "000000";
					when "11100010010111100" => rgb <= "000000";
					when "11100010010111101" => rgb <= "000000";
					when "11100010010111110" => rgb <= "000000";
					when "11100010010111111" => rgb <= "000000";
					when "11100010011000000" => rgb <= "000000";
					when "11100010011000001" => rgb <= "000000";
					when "11100010011000010" => rgb <= "000000";
					when "11100010011000011" => rgb <= "000000";
					when "11100010011000100" => rgb <= "000000";
					when "11100010011000101" => rgb <= "000000";
					when "11100010011000110" => rgb <= "000000";
					when "11100010011000111" => rgb <= "000000";
					when "11100010011001000" => rgb <= "000000";
					when "11100010011001001" => rgb <= "000000";
					when "11100010011001010" => rgb <= "000000";
					when "11100010011001011" => rgb <= "000000";
					when "11100010011001100" => rgb <= "000000";
					when "11100010011001101" => rgb <= "000000";
					when "11100010011001110" => rgb <= "000000";
					when "11100010011001111" => rgb <= "000000";
					when "11100010011010000" => rgb <= "000000";
					when "11100010011010001" => rgb <= "000000";
					when "11100010011010010" => rgb <= "000000";
					when "11100010011010011" => rgb <= "000000";
					when "11100010011010100" => rgb <= "000000";
					when "11100010011010101" => rgb <= "000000";
					when "11100010011010110" => rgb <= "000000";
					when "11100010011010111" => rgb <= "000000";
					when "11100010011011000" => rgb <= "000000";
					when "11100010011011001" => rgb <= "000000";
					when "11100010011011010" => rgb <= "000000";
					when "11100010011011011" => rgb <= "000000";
					when "11100010011011100" => rgb <= "000000";
					when "11100010011011101" => rgb <= "000000";
					when "11100010011011110" => rgb <= "000000";
					when "11100010011011111" => rgb <= "000000";
					when "11100010011100000" => rgb <= "000000";
					when "11100010011100001" => rgb <= "000000";
					when "11100010011100010" => rgb <= "000000";
					when "11100010011100011" => rgb <= "000000";
					when "11100010011100100" => rgb <= "000000";
					when "11100010011100101" => rgb <= "000000";
					when "11100010011100110" => rgb <= "000000";
					when "11100010011100111" => rgb <= "000000";
					when "11100010011101000" => rgb <= "000000";
					when "11100010011101001" => rgb <= "000000";
					when "11100010011101010" => rgb <= "000000";
					when "11100010011101011" => rgb <= "000000";
					when "11100010011101100" => rgb <= "000000";
					when "11100010011101101" => rgb <= "000000";
					when "11100010011101110" => rgb <= "000000";
					when "11100010011101111" => rgb <= "000000";
					when "11100010011110000" => rgb <= "000000";
					when "11100010011110001" => rgb <= "000000";
					when "11100010011110010" => rgb <= "000000";
					when "11100010011110011" => rgb <= "000000";
					when "11100010011110100" => rgb <= "000000";
					when "11100010011110101" => rgb <= "000000";
					when "11100010011110110" => rgb <= "000000";
					when "11100010011110111" => rgb <= "000000";
					when "11100010011111000" => rgb <= "000000";
					when "11100010011111001" => rgb <= "000000";
					when "11100010011111010" => rgb <= "000000";
					when "11100010011111011" => rgb <= "000000";
					when "11100010011111100" => rgb <= "000000";
					when "11100010011111101" => rgb <= "000000";
					when "11100010011111110" => rgb <= "000000";
					when "11100010011111111" => rgb <= "000000";
					when "11100010100000000" => rgb <= "000000";
					when "11100010100000001" => rgb <= "000000";
					when "11100010100000010" => rgb <= "000000";
					when "11100010100000011" => rgb <= "000000";
					when "11100010100000100" => rgb <= "000000";
					when "11100010100000101" => rgb <= "000000";
					when "11100010100000110" => rgb <= "000000";
					when "11100010100000111" => rgb <= "000000";
					when "11100010100001000" => rgb <= "000000";
					when "11100010100001001" => rgb <= "000000";
					when "11100010100001010" => rgb <= "000000";
					when "11100010100001011" => rgb <= "000000";
					when "11100010100001100" => rgb <= "000000";
					when "11100010100001101" => rgb <= "000000";
					when "11100010100001110" => rgb <= "000000";
					when "11100010100001111" => rgb <= "000000";
					when "11100010100010000" => rgb <= "000000";
					when "11100010100010001" => rgb <= "000000";
					when "11100010100010010" => rgb <= "000000";
					when "11100010100010011" => rgb <= "000000";
					when "11100010100010100" => rgb <= "000000";
					when "11100010100010101" => rgb <= "000000";
					when "11100010100010110" => rgb <= "000000";
					when "11100010100010111" => rgb <= "000000";
					when "11100010100011000" => rgb <= "000000";
					when "11100010100011001" => rgb <= "000000";
					when "11100010100011010" => rgb <= "000000";
					when "11100010100011011" => rgb <= "000000";
					when "11100010100011100" => rgb <= "000000";
					when "11100010100011101" => rgb <= "000000";
					when "11100010100011110" => rgb <= "000000";
					when "11100010100011111" => rgb <= "000000";
					when "11100010100100000" => rgb <= "000000";
					when "11100010100100001" => rgb <= "000000";
					when "11100010100100010" => rgb <= "000000";
					when "11100010100100011" => rgb <= "000000";
					when "11100010100100100" => rgb <= "000000";
					when "11100010100100101" => rgb <= "000000";
					when "11100010100100110" => rgb <= "000000";
					when "11100010100100111" => rgb <= "000000";
					when "11100010100101000" => rgb <= "000000";
					when "11100010100101001" => rgb <= "000000";
					when "11100010100101010" => rgb <= "000000";
					when "11100010100101011" => rgb <= "000000";
					when "11100010100101100" => rgb <= "000000";
					when "11100010100101101" => rgb <= "000000";
					when "11100010100101110" => rgb <= "000000";
					when "11100010100101111" => rgb <= "000000";
					when "11100010100110000" => rgb <= "000000";
					when "11100010100110001" => rgb <= "000000";
					when "11100010100110010" => rgb <= "000000";
					when "11100010100110011" => rgb <= "000000";
					when "11100010100110100" => rgb <= "000000";
					when "11100010100110101" => rgb <= "000000";
					when "11100010100110110" => rgb <= "000000";
					when "11100010100110111" => rgb <= "000000";
					when "11100010100111000" => rgb <= "000000";
					when "11100010100111001" => rgb <= "000000";
					when "11100010100111010" => rgb <= "000000";
					when "11100010100111011" => rgb <= "000000";
					when "11100010100111100" => rgb <= "000000";
					when "11100010100111101" => rgb <= "000000";
					when "11100010100111110" => rgb <= "000000";
					when "11100010100111111" => rgb <= "000000";
					when "11100011000000000" => rgb <= "000000";
					when "11100011000000001" => rgb <= "000000";
					when "11100011000000010" => rgb <= "000000";
					when "11100011000000011" => rgb <= "000000";
					when "11100011000000100" => rgb <= "000000";
					when "11100011000000101" => rgb <= "000000";
					when "11100011000000110" => rgb <= "000000";
					when "11100011000000111" => rgb <= "000000";
					when "11100011000001000" => rgb <= "000000";
					when "11100011000001001" => rgb <= "000000";
					when "11100011000001010" => rgb <= "000000";
					when "11100011000001011" => rgb <= "000000";
					when "11100011000001100" => rgb <= "000000";
					when "11100011000001101" => rgb <= "000000";
					when "11100011000001110" => rgb <= "000000";
					when "11100011000001111" => rgb <= "000000";
					when "11100011000010000" => rgb <= "000000";
					when "11100011000010001" => rgb <= "000000";
					when "11100011000010010" => rgb <= "000000";
					when "11100011000010011" => rgb <= "000000";
					when "11100011000010100" => rgb <= "000000";
					when "11100011000010101" => rgb <= "000000";
					when "11100011000010110" => rgb <= "000000";
					when "11100011000010111" => rgb <= "000000";
					when "11100011000011000" => rgb <= "000000";
					when "11100011000011001" => rgb <= "000000";
					when "11100011000011010" => rgb <= "000000";
					when "11100011000011011" => rgb <= "000000";
					when "11100011000011100" => rgb <= "000000";
					when "11100011000011101" => rgb <= "000000";
					when "11100011000011110" => rgb <= "000000";
					when "11100011000011111" => rgb <= "000000";
					when "11100011000100000" => rgb <= "000000";
					when "11100011000100001" => rgb <= "000000";
					when "11100011000100010" => rgb <= "000000";
					when "11100011000100011" => rgb <= "000000";
					when "11100011000100100" => rgb <= "000000";
					when "11100011000100101" => rgb <= "000000";
					when "11100011000100110" => rgb <= "000000";
					when "11100011000100111" => rgb <= "000000";
					when "11100011000101000" => rgb <= "000000";
					when "11100011000101001" => rgb <= "000000";
					when "11100011000101010" => rgb <= "000000";
					when "11100011000101011" => rgb <= "000000";
					when "11100011000101100" => rgb <= "000000";
					when "11100011000101101" => rgb <= "000000";
					when "11100011000101110" => rgb <= "000000";
					when "11100011000101111" => rgb <= "000000";
					when "11100011000110000" => rgb <= "000000";
					when "11100011000110001" => rgb <= "000000";
					when "11100011000110010" => rgb <= "000000";
					when "11100011000110011" => rgb <= "000000";
					when "11100011000110100" => rgb <= "000000";
					when "11100011000110101" => rgb <= "000000";
					when "11100011000110110" => rgb <= "000000";
					when "11100011000110111" => rgb <= "000000";
					when "11100011000111000" => rgb <= "000000";
					when "11100011000111001" => rgb <= "000000";
					when "11100011000111010" => rgb <= "000000";
					when "11100011000111011" => rgb <= "000000";
					when "11100011000111100" => rgb <= "000000";
					when "11100011000111101" => rgb <= "000000";
					when "11100011000111110" => rgb <= "000000";
					when "11100011000111111" => rgb <= "000000";
					when "11100011001000000" => rgb <= "000000";
					when "11100011001000001" => rgb <= "000000";
					when "11100011001000010" => rgb <= "000000";
					when "11100011001000011" => rgb <= "000000";
					when "11100011001000100" => rgb <= "000000";
					when "11100011001000101" => rgb <= "000000";
					when "11100011001000110" => rgb <= "000000";
					when "11100011001000111" => rgb <= "000000";
					when "11100011001001000" => rgb <= "000000";
					when "11100011001001001" => rgb <= "000000";
					when "11100011001001010" => rgb <= "000000";
					when "11100011001001011" => rgb <= "000000";
					when "11100011001001100" => rgb <= "000000";
					when "11100011001001101" => rgb <= "000000";
					when "11100011001001110" => rgb <= "000000";
					when "11100011001001111" => rgb <= "000000";
					when "11100011001010000" => rgb <= "000000";
					when "11100011001010001" => rgb <= "000000";
					when "11100011001010010" => rgb <= "000000";
					when "11100011001010011" => rgb <= "000000";
					when "11100011001010100" => rgb <= "000000";
					when "11100011001010101" => rgb <= "000000";
					when "11100011001010110" => rgb <= "000000";
					when "11100011001010111" => rgb <= "000000";
					when "11100011001011000" => rgb <= "000000";
					when "11100011001011001" => rgb <= "000000";
					when "11100011001011010" => rgb <= "000000";
					when "11100011001011011" => rgb <= "000000";
					when "11100011001011100" => rgb <= "000000";
					when "11100011001011101" => rgb <= "000000";
					when "11100011001011110" => rgb <= "000000";
					when "11100011001011111" => rgb <= "000000";
					when "11100011001100000" => rgb <= "000000";
					when "11100011001100001" => rgb <= "000000";
					when "11100011001100010" => rgb <= "000000";
					when "11100011001100011" => rgb <= "000000";
					when "11100011001100100" => rgb <= "000000";
					when "11100011001100101" => rgb <= "000000";
					when "11100011001100110" => rgb <= "000000";
					when "11100011001100111" => rgb <= "000000";
					when "11100011001101000" => rgb <= "000000";
					when "11100011001101001" => rgb <= "000000";
					when "11100011001101010" => rgb <= "000000";
					when "11100011001101011" => rgb <= "000000";
					when "11100011001101100" => rgb <= "000000";
					when "11100011001101101" => rgb <= "000000";
					when "11100011001101110" => rgb <= "000000";
					when "11100011001101111" => rgb <= "000000";
					when "11100011001110000" => rgb <= "000000";
					when "11100011001110001" => rgb <= "000000";
					when "11100011001110010" => rgb <= "000000";
					when "11100011001110011" => rgb <= "000000";
					when "11100011001110100" => rgb <= "000000";
					when "11100011001110101" => rgb <= "000000";
					when "11100011001110110" => rgb <= "000000";
					when "11100011001110111" => rgb <= "000000";
					when "11100011001111000" => rgb <= "000000";
					when "11100011001111001" => rgb <= "000000";
					when "11100011001111010" => rgb <= "000000";
					when "11100011001111011" => rgb <= "000000";
					when "11100011001111100" => rgb <= "000000";
					when "11100011001111101" => rgb <= "000000";
					when "11100011001111110" => rgb <= "000000";
					when "11100011001111111" => rgb <= "000000";
					when "11100011010000000" => rgb <= "000000";
					when "11100011010000001" => rgb <= "000000";
					when "11100011010000010" => rgb <= "000000";
					when "11100011010000011" => rgb <= "000000";
					when "11100011010000100" => rgb <= "000000";
					when "11100011010000101" => rgb <= "000000";
					when "11100011010000110" => rgb <= "000000";
					when "11100011010000111" => rgb <= "000000";
					when "11100011010001000" => rgb <= "000000";
					when "11100011010001001" => rgb <= "000000";
					when "11100011010001010" => rgb <= "000000";
					when "11100011010001011" => rgb <= "000000";
					when "11100011010001100" => rgb <= "000000";
					when "11100011010001101" => rgb <= "000000";
					when "11100011010001110" => rgb <= "000000";
					when "11100011010001111" => rgb <= "000000";
					when "11100011010010000" => rgb <= "000000";
					when "11100011010010001" => rgb <= "000000";
					when "11100011010010010" => rgb <= "000000";
					when "11100011010010011" => rgb <= "000000";
					when "11100011010010100" => rgb <= "000000";
					when "11100011010010101" => rgb <= "000000";
					when "11100011010010110" => rgb <= "000000";
					when "11100011010010111" => rgb <= "000000";
					when "11100011010011000" => rgb <= "000000";
					when "11100011010011001" => rgb <= "000000";
					when "11100011010011010" => rgb <= "000000";
					when "11100011010011011" => rgb <= "000000";
					when "11100011010011100" => rgb <= "000000";
					when "11100011010011101" => rgb <= "000000";
					when "11100011010011110" => rgb <= "000000";
					when "11100011010011111" => rgb <= "000000";
					when "11100011010100000" => rgb <= "000000";
					when "11100011010100001" => rgb <= "000000";
					when "11100011010100010" => rgb <= "000000";
					when "11100011010100011" => rgb <= "000000";
					when "11100011010100100" => rgb <= "000000";
					when "11100011010100101" => rgb <= "000000";
					when "11100011010100110" => rgb <= "000000";
					when "11100011010100111" => rgb <= "000000";
					when "11100011010101000" => rgb <= "000000";
					when "11100011010101001" => rgb <= "000000";
					when "11100011010101010" => rgb <= "000000";
					when "11100011010101011" => rgb <= "000000";
					when "11100011010101100" => rgb <= "000000";
					when "11100011010101101" => rgb <= "000000";
					when "11100011010101110" => rgb <= "000000";
					when "11100011010101111" => rgb <= "000000";
					when "11100011010110000" => rgb <= "000000";
					when "11100011010110001" => rgb <= "000000";
					when "11100011010110010" => rgb <= "000000";
					when "11100011010110011" => rgb <= "000000";
					when "11100011010110100" => rgb <= "000000";
					when "11100011010110101" => rgb <= "000000";
					when "11100011010110110" => rgb <= "000000";
					when "11100011010110111" => rgb <= "000000";
					when "11100011010111000" => rgb <= "000000";
					when "11100011010111001" => rgb <= "000000";
					when "11100011010111010" => rgb <= "000000";
					when "11100011010111011" => rgb <= "000000";
					when "11100011010111100" => rgb <= "000000";
					when "11100011010111101" => rgb <= "000000";
					when "11100011010111110" => rgb <= "000000";
					when "11100011010111111" => rgb <= "000000";
					when "11100011011000000" => rgb <= "000000";
					when "11100011011000001" => rgb <= "000000";
					when "11100011011000010" => rgb <= "000000";
					when "11100011011000011" => rgb <= "000000";
					when "11100011011000100" => rgb <= "000000";
					when "11100011011000101" => rgb <= "000000";
					when "11100011011000110" => rgb <= "000000";
					when "11100011011000111" => rgb <= "000000";
					when "11100011011001000" => rgb <= "000000";
					when "11100011011001001" => rgb <= "000000";
					when "11100011011001010" => rgb <= "000000";
					when "11100011011001011" => rgb <= "000000";
					when "11100011011001100" => rgb <= "000000";
					when "11100011011001101" => rgb <= "000000";
					when "11100011011001110" => rgb <= "000000";
					when "11100011011001111" => rgb <= "000000";
					when "11100011011010000" => rgb <= "000000";
					when "11100011011010001" => rgb <= "000000";
					when "11100011011010010" => rgb <= "000000";
					when "11100011011010011" => rgb <= "000000";
					when "11100011011010100" => rgb <= "000000";
					when "11100011011010101" => rgb <= "000000";
					when "11100011011010110" => rgb <= "000000";
					when "11100011011010111" => rgb <= "000000";
					when "11100011011011000" => rgb <= "000000";
					when "11100011011011001" => rgb <= "000000";
					when "11100011011011010" => rgb <= "000000";
					when "11100011011011011" => rgb <= "000000";
					when "11100011011011100" => rgb <= "000000";
					when "11100011011011101" => rgb <= "000000";
					when "11100011011011110" => rgb <= "000000";
					when "11100011011011111" => rgb <= "000000";
					when "11100011011100000" => rgb <= "000000";
					when "11100011011100001" => rgb <= "000000";
					when "11100011011100010" => rgb <= "000000";
					when "11100011011100011" => rgb <= "000000";
					when "11100011011100100" => rgb <= "000000";
					when "11100011011100101" => rgb <= "000000";
					when "11100011011100110" => rgb <= "000000";
					when "11100011011100111" => rgb <= "000000";
					when "11100011011101000" => rgb <= "000000";
					when "11100011011101001" => rgb <= "000000";
					when "11100011011101010" => rgb <= "000000";
					when "11100011011101011" => rgb <= "000000";
					when "11100011011101100" => rgb <= "000000";
					when "11100011011101101" => rgb <= "000000";
					when "11100011011101110" => rgb <= "000000";
					when "11100011011101111" => rgb <= "000000";
					when "11100011011110000" => rgb <= "000000";
					when "11100011011110001" => rgb <= "000000";
					when "11100011011110010" => rgb <= "000000";
					when "11100011011110011" => rgb <= "000000";
					when "11100011011110100" => rgb <= "000000";
					when "11100011011110101" => rgb <= "000000";
					when "11100011011110110" => rgb <= "000000";
					when "11100011011110111" => rgb <= "000000";
					when "11100011011111000" => rgb <= "000000";
					when "11100011011111001" => rgb <= "000000";
					when "11100011011111010" => rgb <= "000000";
					when "11100011011111011" => rgb <= "000000";
					when "11100011011111100" => rgb <= "000000";
					when "11100011011111101" => rgb <= "000000";
					when "11100011011111110" => rgb <= "000000";
					when "11100011011111111" => rgb <= "000000";
					when "11100011100000000" => rgb <= "000000";
					when "11100011100000001" => rgb <= "000000";
					when "11100011100000010" => rgb <= "000000";
					when "11100011100000011" => rgb <= "000000";
					when "11100011100000100" => rgb <= "000000";
					when "11100011100000101" => rgb <= "000000";
					when "11100011100000110" => rgb <= "000000";
					when "11100011100000111" => rgb <= "000000";
					when "11100011100001000" => rgb <= "000000";
					when "11100011100001001" => rgb <= "000000";
					when "11100011100001010" => rgb <= "000000";
					when "11100011100001011" => rgb <= "000000";
					when "11100011100001100" => rgb <= "000000";
					when "11100011100001101" => rgb <= "000000";
					when "11100011100001110" => rgb <= "000000";
					when "11100011100001111" => rgb <= "000000";
					when "11100011100010000" => rgb <= "000000";
					when "11100011100010001" => rgb <= "000000";
					when "11100011100010010" => rgb <= "000000";
					when "11100011100010011" => rgb <= "000000";
					when "11100011100010100" => rgb <= "000000";
					when "11100011100010101" => rgb <= "000000";
					when "11100011100010110" => rgb <= "000000";
					when "11100011100010111" => rgb <= "000000";
					when "11100011100011000" => rgb <= "000000";
					when "11100011100011001" => rgb <= "000000";
					when "11100011100011010" => rgb <= "000000";
					when "11100011100011011" => rgb <= "000000";
					when "11100011100011100" => rgb <= "000000";
					when "11100011100011101" => rgb <= "000000";
					when "11100011100011110" => rgb <= "000000";
					when "11100011100011111" => rgb <= "000000";
					when "11100011100100000" => rgb <= "000000";
					when "11100011100100001" => rgb <= "000000";
					when "11100011100100010" => rgb <= "000000";
					when "11100011100100011" => rgb <= "000000";
					when "11100011100100100" => rgb <= "000000";
					when "11100011100100101" => rgb <= "000000";
					when "11100011100100110" => rgb <= "000000";
					when "11100011100100111" => rgb <= "000000";
					when "11100011100101000" => rgb <= "000000";
					when "11100011100101001" => rgb <= "000000";
					when "11100011100101010" => rgb <= "000000";
					when "11100011100101011" => rgb <= "000000";
					when "11100011100101100" => rgb <= "000000";
					when "11100011100101101" => rgb <= "000000";
					when "11100011100101110" => rgb <= "000000";
					when "11100011100101111" => rgb <= "000000";
					when "11100011100110000" => rgb <= "000000";
					when "11100011100110001" => rgb <= "000000";
					when "11100011100110010" => rgb <= "000000";
					when "11100011100110011" => rgb <= "000000";
					when "11100011100110100" => rgb <= "000000";
					when "11100011100110101" => rgb <= "000000";
					when "11100011100110110" => rgb <= "000000";
					when "11100011100110111" => rgb <= "000000";
					when "11100011100111000" => rgb <= "000000";
					when "11100011100111001" => rgb <= "000000";
					when "11100011100111010" => rgb <= "000000";
					when "11100011100111011" => rgb <= "000000";
					when "11100011100111100" => rgb <= "000000";
					when "11100011100111101" => rgb <= "000000";
					when "11100011100111110" => rgb <= "000000";
					when "11100011100111111" => rgb <= "000000";
					when "11100100000000000" => rgb <= "000000";
					when "11100100000000001" => rgb <= "000000";
					when "11100100000000010" => rgb <= "000000";
					when "11100100000000011" => rgb <= "000000";
					when "11100100000000100" => rgb <= "000000";
					when "11100100000000101" => rgb <= "000000";
					when "11100100000000110" => rgb <= "000000";
					when "11100100000000111" => rgb <= "000000";
					when "11100100000001000" => rgb <= "000000";
					when "11100100000001001" => rgb <= "000000";
					when "11100100000001010" => rgb <= "000000";
					when "11100100000001011" => rgb <= "000000";
					when "11100100000001100" => rgb <= "000000";
					when "11100100000001101" => rgb <= "000000";
					when "11100100000001110" => rgb <= "000000";
					when "11100100000001111" => rgb <= "000000";
					when "11100100000010000" => rgb <= "000000";
					when "11100100000010001" => rgb <= "000000";
					when "11100100000010010" => rgb <= "000000";
					when "11100100000010011" => rgb <= "000000";
					when "11100100000010100" => rgb <= "000000";
					when "11100100000010101" => rgb <= "000000";
					when "11100100000010110" => rgb <= "000000";
					when "11100100000010111" => rgb <= "000000";
					when "11100100000011000" => rgb <= "000000";
					when "11100100000011001" => rgb <= "000000";
					when "11100100000011010" => rgb <= "000000";
					when "11100100000011011" => rgb <= "000000";
					when "11100100000011100" => rgb <= "000000";
					when "11100100000011101" => rgb <= "000000";
					when "11100100000011110" => rgb <= "000000";
					when "11100100000011111" => rgb <= "000000";
					when "11100100000100000" => rgb <= "000000";
					when "11100100000100001" => rgb <= "000000";
					when "11100100000100010" => rgb <= "000000";
					when "11100100000100011" => rgb <= "000000";
					when "11100100000100100" => rgb <= "000000";
					when "11100100000100101" => rgb <= "000000";
					when "11100100000100110" => rgb <= "000000";
					when "11100100000100111" => rgb <= "000000";
					when "11100100000101000" => rgb <= "000000";
					when "11100100000101001" => rgb <= "000000";
					when "11100100000101010" => rgb <= "000000";
					when "11100100000101011" => rgb <= "000000";
					when "11100100000101100" => rgb <= "000000";
					when "11100100000101101" => rgb <= "000000";
					when "11100100000101110" => rgb <= "000000";
					when "11100100000101111" => rgb <= "000000";
					when "11100100000110000" => rgb <= "000000";
					when "11100100000110001" => rgb <= "000000";
					when "11100100000110010" => rgb <= "000000";
					when "11100100000110011" => rgb <= "000000";
					when "11100100000110100" => rgb <= "000000";
					when "11100100000110101" => rgb <= "000000";
					when "11100100000110110" => rgb <= "000000";
					when "11100100000110111" => rgb <= "000000";
					when "11100100000111000" => rgb <= "000000";
					when "11100100000111001" => rgb <= "000000";
					when "11100100000111010" => rgb <= "000000";
					when "11100100000111011" => rgb <= "000000";
					when "11100100000111100" => rgb <= "000000";
					when "11100100000111101" => rgb <= "000000";
					when "11100100000111110" => rgb <= "000000";
					when "11100100000111111" => rgb <= "000000";
					when "11100100001000000" => rgb <= "000000";
					when "11100100001000001" => rgb <= "000000";
					when "11100100001000010" => rgb <= "000000";
					when "11100100001000011" => rgb <= "000000";
					when "11100100001000100" => rgb <= "000000";
					when "11100100001000101" => rgb <= "000000";
					when "11100100001000110" => rgb <= "000000";
					when "11100100001000111" => rgb <= "000000";
					when "11100100001001000" => rgb <= "000000";
					when "11100100001001001" => rgb <= "000000";
					when "11100100001001010" => rgb <= "000000";
					when "11100100001001011" => rgb <= "000000";
					when "11100100001001100" => rgb <= "000000";
					when "11100100001001101" => rgb <= "000000";
					when "11100100001001110" => rgb <= "000000";
					when "11100100001001111" => rgb <= "000000";
					when "11100100001010000" => rgb <= "000000";
					when "11100100001010001" => rgb <= "000000";
					when "11100100001010010" => rgb <= "000000";
					when "11100100001010011" => rgb <= "000000";
					when "11100100001010100" => rgb <= "000000";
					when "11100100001010101" => rgb <= "000000";
					when "11100100001010110" => rgb <= "000000";
					when "11100100001010111" => rgb <= "000000";
					when "11100100001011000" => rgb <= "000000";
					when "11100100001011001" => rgb <= "000000";
					when "11100100001011010" => rgb <= "000000";
					when "11100100001011011" => rgb <= "000000";
					when "11100100001011100" => rgb <= "000000";
					when "11100100001011101" => rgb <= "000000";
					when "11100100001011110" => rgb <= "000000";
					when "11100100001011111" => rgb <= "000000";
					when "11100100001100000" => rgb <= "000000";
					when "11100100001100001" => rgb <= "000000";
					when "11100100001100010" => rgb <= "000000";
					when "11100100001100011" => rgb <= "000000";
					when "11100100001100100" => rgb <= "000000";
					when "11100100001100101" => rgb <= "000000";
					when "11100100001100110" => rgb <= "000000";
					when "11100100001100111" => rgb <= "000000";
					when "11100100001101000" => rgb <= "000000";
					when "11100100001101001" => rgb <= "000000";
					when "11100100001101010" => rgb <= "000000";
					when "11100100001101011" => rgb <= "000000";
					when "11100100001101100" => rgb <= "000000";
					when "11100100001101101" => rgb <= "000000";
					when "11100100001101110" => rgb <= "000000";
					when "11100100001101111" => rgb <= "000000";
					when "11100100001110000" => rgb <= "000000";
					when "11100100001110001" => rgb <= "000000";
					when "11100100001110010" => rgb <= "000000";
					when "11100100001110011" => rgb <= "000000";
					when "11100100001110100" => rgb <= "000000";
					when "11100100001110101" => rgb <= "000000";
					when "11100100001110110" => rgb <= "000000";
					when "11100100001110111" => rgb <= "000000";
					when "11100100001111000" => rgb <= "000000";
					when "11100100001111001" => rgb <= "000000";
					when "11100100001111010" => rgb <= "000000";
					when "11100100001111011" => rgb <= "000000";
					when "11100100001111100" => rgb <= "000000";
					when "11100100001111101" => rgb <= "000000";
					when "11100100001111110" => rgb <= "000000";
					when "11100100001111111" => rgb <= "000000";
					when "11100100010000000" => rgb <= "000000";
					when "11100100010000001" => rgb <= "000000";
					when "11100100010000010" => rgb <= "000000";
					when "11100100010000011" => rgb <= "000000";
					when "11100100010000100" => rgb <= "000000";
					when "11100100010000101" => rgb <= "000000";
					when "11100100010000110" => rgb <= "000000";
					when "11100100010000111" => rgb <= "000000";
					when "11100100010001000" => rgb <= "000000";
					when "11100100010001001" => rgb <= "000000";
					when "11100100010001010" => rgb <= "000000";
					when "11100100010001011" => rgb <= "000000";
					when "11100100010001100" => rgb <= "000000";
					when "11100100010001101" => rgb <= "000000";
					when "11100100010001110" => rgb <= "000000";
					when "11100100010001111" => rgb <= "000000";
					when "11100100010010000" => rgb <= "000000";
					when "11100100010010001" => rgb <= "000000";
					when "11100100010010010" => rgb <= "000000";
					when "11100100010010011" => rgb <= "000000";
					when "11100100010010100" => rgb <= "000000";
					when "11100100010010101" => rgb <= "000000";
					when "11100100010010110" => rgb <= "000000";
					when "11100100010010111" => rgb <= "000000";
					when "11100100010011000" => rgb <= "000000";
					when "11100100010011001" => rgb <= "000000";
					when "11100100010011010" => rgb <= "000000";
					when "11100100010011011" => rgb <= "000000";
					when "11100100010011100" => rgb <= "000000";
					when "11100100010011101" => rgb <= "000000";
					when "11100100010011110" => rgb <= "000000";
					when "11100100010011111" => rgb <= "000000";
					when "11100100010100000" => rgb <= "000000";
					when "11100100010100001" => rgb <= "000000";
					when "11100100010100010" => rgb <= "000000";
					when "11100100010100011" => rgb <= "000000";
					when "11100100010100100" => rgb <= "000000";
					when "11100100010100101" => rgb <= "000000";
					when "11100100010100110" => rgb <= "000000";
					when "11100100010100111" => rgb <= "000000";
					when "11100100010101000" => rgb <= "000000";
					when "11100100010101001" => rgb <= "000000";
					when "11100100010101010" => rgb <= "000000";
					when "11100100010101011" => rgb <= "000000";
					when "11100100010101100" => rgb <= "000000";
					when "11100100010101101" => rgb <= "000000";
					when "11100100010101110" => rgb <= "000000";
					when "11100100010101111" => rgb <= "000000";
					when "11100100010110000" => rgb <= "000000";
					when "11100100010110001" => rgb <= "000000";
					when "11100100010110010" => rgb <= "000000";
					when "11100100010110011" => rgb <= "000000";
					when "11100100010110100" => rgb <= "000000";
					when "11100100010110101" => rgb <= "000000";
					when "11100100010110110" => rgb <= "000000";
					when "11100100010110111" => rgb <= "000000";
					when "11100100010111000" => rgb <= "000000";
					when "11100100010111001" => rgb <= "000000";
					when "11100100010111010" => rgb <= "000000";
					when "11100100010111011" => rgb <= "000000";
					when "11100100010111100" => rgb <= "000000";
					when "11100100010111101" => rgb <= "000000";
					when "11100100010111110" => rgb <= "000000";
					when "11100100010111111" => rgb <= "000000";
					when "11100100011000000" => rgb <= "000000";
					when "11100100011000001" => rgb <= "000000";
					when "11100100011000010" => rgb <= "000000";
					when "11100100011000011" => rgb <= "000000";
					when "11100100011000100" => rgb <= "000000";
					when "11100100011000101" => rgb <= "000000";
					when "11100100011000110" => rgb <= "000000";
					when "11100100011000111" => rgb <= "000000";
					when "11100100011001000" => rgb <= "000000";
					when "11100100011001001" => rgb <= "000000";
					when "11100100011001010" => rgb <= "000000";
					when "11100100011001011" => rgb <= "000000";
					when "11100100011001100" => rgb <= "000000";
					when "11100100011001101" => rgb <= "000000";
					when "11100100011001110" => rgb <= "000000";
					when "11100100011001111" => rgb <= "000000";
					when "11100100011010000" => rgb <= "000000";
					when "11100100011010001" => rgb <= "000000";
					when "11100100011010010" => rgb <= "000000";
					when "11100100011010011" => rgb <= "000000";
					when "11100100011010100" => rgb <= "000000";
					when "11100100011010101" => rgb <= "000000";
					when "11100100011010110" => rgb <= "000000";
					when "11100100011010111" => rgb <= "000000";
					when "11100100011011000" => rgb <= "000000";
					when "11100100011011001" => rgb <= "000000";
					when "11100100011011010" => rgb <= "000000";
					when "11100100011011011" => rgb <= "000000";
					when "11100100011011100" => rgb <= "000000";
					when "11100100011011101" => rgb <= "000000";
					when "11100100011011110" => rgb <= "000000";
					when "11100100011011111" => rgb <= "000000";
					when "11100100011100000" => rgb <= "000000";
					when "11100100011100001" => rgb <= "000000";
					when "11100100011100010" => rgb <= "000000";
					when "11100100011100011" => rgb <= "000000";
					when "11100100011100100" => rgb <= "000000";
					when "11100100011100101" => rgb <= "000000";
					when "11100100011100110" => rgb <= "000000";
					when "11100100011100111" => rgb <= "000000";
					when "11100100011101000" => rgb <= "000000";
					when "11100100011101001" => rgb <= "000000";
					when "11100100011101010" => rgb <= "000000";
					when "11100100011101011" => rgb <= "000000";
					when "11100100011101100" => rgb <= "000000";
					when "11100100011101101" => rgb <= "000000";
					when "11100100011101110" => rgb <= "000000";
					when "11100100011101111" => rgb <= "000000";
					when "11100100011110000" => rgb <= "000000";
					when "11100100011110001" => rgb <= "000000";
					when "11100100011110010" => rgb <= "000000";
					when "11100100011110011" => rgb <= "000000";
					when "11100100011110100" => rgb <= "000000";
					when "11100100011110101" => rgb <= "000000";
					when "11100100011110110" => rgb <= "000000";
					when "11100100011110111" => rgb <= "000000";
					when "11100100011111000" => rgb <= "000000";
					when "11100100011111001" => rgb <= "000000";
					when "11100100011111010" => rgb <= "000000";
					when "11100100011111011" => rgb <= "000000";
					when "11100100011111100" => rgb <= "000000";
					when "11100100011111101" => rgb <= "000000";
					when "11100100011111110" => rgb <= "000000";
					when "11100100011111111" => rgb <= "000000";
					when "11100100100000000" => rgb <= "000000";
					when "11100100100000001" => rgb <= "000000";
					when "11100100100000010" => rgb <= "000000";
					when "11100100100000011" => rgb <= "000000";
					when "11100100100000100" => rgb <= "000000";
					when "11100100100000101" => rgb <= "000000";
					when "11100100100000110" => rgb <= "000000";
					when "11100100100000111" => rgb <= "000000";
					when "11100100100001000" => rgb <= "000000";
					when "11100100100001001" => rgb <= "000000";
					when "11100100100001010" => rgb <= "000000";
					when "11100100100001011" => rgb <= "000000";
					when "11100100100001100" => rgb <= "000000";
					when "11100100100001101" => rgb <= "000000";
					when "11100100100001110" => rgb <= "000000";
					when "11100100100001111" => rgb <= "000000";
					when "11100100100010000" => rgb <= "000000";
					when "11100100100010001" => rgb <= "000000";
					when "11100100100010010" => rgb <= "000000";
					when "11100100100010011" => rgb <= "000000";
					when "11100100100010100" => rgb <= "000000";
					when "11100100100010101" => rgb <= "000000";
					when "11100100100010110" => rgb <= "000000";
					when "11100100100010111" => rgb <= "000000";
					when "11100100100011000" => rgb <= "000000";
					when "11100100100011001" => rgb <= "000000";
					when "11100100100011010" => rgb <= "000000";
					when "11100100100011011" => rgb <= "000000";
					when "11100100100011100" => rgb <= "000000";
					when "11100100100011101" => rgb <= "000000";
					when "11100100100011110" => rgb <= "000000";
					when "11100100100011111" => rgb <= "000000";
					when "11100100100100000" => rgb <= "000000";
					when "11100100100100001" => rgb <= "000000";
					when "11100100100100010" => rgb <= "000000";
					when "11100100100100011" => rgb <= "000000";
					when "11100100100100100" => rgb <= "000000";
					when "11100100100100101" => rgb <= "000000";
					when "11100100100100110" => rgb <= "000000";
					when "11100100100100111" => rgb <= "000000";
					when "11100100100101000" => rgb <= "000000";
					when "11100100100101001" => rgb <= "000000";
					when "11100100100101010" => rgb <= "000000";
					when "11100100100101011" => rgb <= "000000";
					when "11100100100101100" => rgb <= "000000";
					when "11100100100101101" => rgb <= "000000";
					when "11100100100101110" => rgb <= "000000";
					when "11100100100101111" => rgb <= "000000";
					when "11100100100110000" => rgb <= "000000";
					when "11100100100110001" => rgb <= "000000";
					when "11100100100110010" => rgb <= "000000";
					when "11100100100110011" => rgb <= "000000";
					when "11100100100110100" => rgb <= "000000";
					when "11100100100110101" => rgb <= "000000";
					when "11100100100110110" => rgb <= "000000";
					when "11100100100110111" => rgb <= "000000";
					when "11100100100111000" => rgb <= "000000";
					when "11100100100111001" => rgb <= "000000";
					when "11100100100111010" => rgb <= "000000";
					when "11100100100111011" => rgb <= "000000";
					when "11100100100111100" => rgb <= "000000";
					when "11100100100111101" => rgb <= "000000";
					when "11100100100111110" => rgb <= "000000";
					when "11100100100111111" => rgb <= "000000";
					when others => rgb <= "000000";
                end case;
            end if;
        end process;   
        addr <=  std_logic_vector(yaddr) & std_logic_vector(xaddr);   
    end;
