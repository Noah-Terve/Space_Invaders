library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alien_sprite is
  port(
    clk : in std_logic;
    xaddr : in unsigned(3 downto 0);
    yaddr : in unsigned(2 downto 0);
	rgb : out std_logic_vector(5 downto 0)
  );
end alien_sprite;

architecture synth of alien_sprite is
    signal addr : std_logic_vector(6 downto 0);         
    begin
        process(clk) is begin
            if rising_edge(clk) then
                case addr is
					when "0000000" => rgb <= "000000";
					when "0000001" => rgb <= "000000";
					when "0000010" => rgb <= "001100";
					when "0000011" => rgb <= "000000";
					when "0000100" => rgb <= "000000";
					when "0000101" => rgb <= "000000";
					when "0000110" => rgb <= "000000";
					when "0000111" => rgb <= "000000";
					when "0001000" => rgb <= "001100";
					when "0001001" => rgb <= "000000";
					when "0001010" => rgb <= "000000";
					when "0010000" => rgb <= "000000";
					when "0010001" => rgb <= "000000";
					when "0010010" => rgb <= "000000";
					when "0010011" => rgb <= "001100";
					when "0010100" => rgb <= "000000";
					when "0010101" => rgb <= "000000";
					when "0010110" => rgb <= "000000";
					when "0010111" => rgb <= "001100";
					when "0011000" => rgb <= "000000";
					when "0011001" => rgb <= "000000";
					when "0011010" => rgb <= "000000";
					when "0100000" => rgb <= "000000";
					when "0100001" => rgb <= "000000";
					when "0100010" => rgb <= "001100";
					when "0100011" => rgb <= "001100";
					when "0100100" => rgb <= "001100";
					when "0100101" => rgb <= "001100";
					when "0100110" => rgb <= "001100";
					when "0100111" => rgb <= "001100";
					when "0101000" => rgb <= "001100";
					when "0101001" => rgb <= "000000";
					when "0101010" => rgb <= "000000";
					when "0110000" => rgb <= "000000";
					when "0110001" => rgb <= "001100";
					when "0110010" => rgb <= "001100";
					when "0110011" => rgb <= "000000";
					when "0110100" => rgb <= "001100";
					when "0110101" => rgb <= "001100";
					when "0110110" => rgb <= "001100";
					when "0110111" => rgb <= "000000";
					when "0111000" => rgb <= "001100";
					when "0111001" => rgb <= "001100";
					when "0111010" => rgb <= "000000";
					when "1000000" => rgb <= "001100";
					when "1000001" => rgb <= "001100";
					when "1000010" => rgb <= "001100";
					when "1000011" => rgb <= "001100";
					when "1000100" => rgb <= "001100";
					when "1000101" => rgb <= "001100";
					when "1000110" => rgb <= "001100";
					when "1000111" => rgb <= "001100";
					when "1001000" => rgb <= "001100";
					when "1001001" => rgb <= "001100";
					when "1001010" => rgb <= "001100";
					when "1010000" => rgb <= "001100";
					when "1010001" => rgb <= "000000";
					when "1010010" => rgb <= "001100";
					when "1010011" => rgb <= "001100";
					when "1010100" => rgb <= "001100";
					when "1010101" => rgb <= "001100";
					when "1010110" => rgb <= "001100";
					when "1010111" => rgb <= "001100";
					when "1011000" => rgb <= "001100";
					when "1011001" => rgb <= "000000";
					when "1011010" => rgb <= "001100";
					when "1100000" => rgb <= "001100";
					when "1100001" => rgb <= "000000";
					when "1100010" => rgb <= "001100";
					when "1100011" => rgb <= "000000";
					when "1100100" => rgb <= "000000";
					when "1100101" => rgb <= "000000";
					when "1100110" => rgb <= "000000";
					when "1100111" => rgb <= "000000";
					when "1101000" => rgb <= "001100";
					when "1101001" => rgb <= "000000";
					when "1101010" => rgb <= "001100";
					when "1110000" => rgb <= "000000";
					when "1110001" => rgb <= "000000";
					when "1110010" => rgb <= "000000";
					when "1110011" => rgb <= "001100";
					when "1110100" => rgb <= "001100";
					when "1110101" => rgb <= "000000";
					when "1110110" => rgb <= "001100";
					when "1110111" => rgb <= "001100";
					when "1111000" => rgb <= "000000";
					when "1111001" => rgb <= "000000";
					when "1111010" => rgb <= "000000";
					when others => rgb <= "000000";
                end case;
            end if;
        end process;   
        addr <=  std_logic_vector(yaddr) & std_logic_vector(xaddr);   
    end;
