library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity alien_sprite is
  port(
    clk : in std_logic;
    xaddr : in unsigned(4 downto 0);
    yaddr : in unsigned(5 downto 0);
	rgb : out std_logic_vector(5 downto 0)
  );
end alien_sprite;

architecture synth of alien_sprite is
    signal addr : std_logic_vector(10 downto 0);         
    begin
        process(clk) is begin
            if rising_edge(clk) then
                case addr is
                    when "0000000000" => rgb <= "000000";
					when "0000000001" => rgb <= "000000";
					when "0000000010" => rgb <= "001100";
					when "0000000011" => rgb <= "000000";
					when "0000000100" => rgb <= "000000";
					when "0000000101" => rgb <= "000000";
					when "0000000110" => rgb <= "000000";
					when "0000000111" => rgb <= "000000";
					when "0000001000" => rgb <= "001100";
					when "0000001001" => rgb <= "000000";
					when "0000001010" => rgb <= "000000";
					when "0001000000" => rgb <= "000000";
					when "0001000001" => rgb <= "000000";
					when "0001000010" => rgb <= "000000";
					when "0001000011" => rgb <= "001100";
					when "0001000100" => rgb <= "000000";
					when "0001000101" => rgb <= "000000";
					when "0001000110" => rgb <= "000000";
					when "0001000111" => rgb <= "001100";
					when "0001001000" => rgb <= "000000";
					when "0001001001" => rgb <= "000000";
					when "0001001010" => rgb <= "000000";
					when "0010000000" => rgb <= "000000";
					when "0010000001" => rgb <= "000000";
					when "0010000010" => rgb <= "001100";
					when "0010000011" => rgb <= "001100";
					when "0010000100" => rgb <= "001100";
					when "0010000101" => rgb <= "001100";
					when "0010000110" => rgb <= "001100";
					when "0010000111" => rgb <= "001100";
					when "0010001000" => rgb <= "001100";
					when "0010001001" => rgb <= "000000";
					when "0010001010" => rgb <= "000000";
					when "0011000000" => rgb <= "000000";
					when "0011000001" => rgb <= "001100";
					when "0011000010" => rgb <= "001100";
					when "0011000011" => rgb <= "000000";
					when "0011000100" => rgb <= "001100";
					when "0011000101" => rgb <= "001100";
					when "0011000110" => rgb <= "001100";
					when "0011000111" => rgb <= "000000";
					when "0011001000" => rgb <= "001100";
					when "0011001001" => rgb <= "001100";
					when "0011001010" => rgb <= "000000";
					when "0100000000" => rgb <= "001100";
					when "0100000001" => rgb <= "001100";
					when "0100000010" => rgb <= "001100";
					when "0100000011" => rgb <= "001100";
					when "0100000100" => rgb <= "001100";
					when "0100000101" => rgb <= "001100";
					when "0100000110" => rgb <= "001100";
					when "0100000111" => rgb <= "001100";
					when "0100001000" => rgb <= "001100";
					when "0100001001" => rgb <= "001100";
					when "0100001010" => rgb <= "001100";
					when "0101000000" => rgb <= "001100";
					when "0101000001" => rgb <= "000000";
					when "0101000010" => rgb <= "001100";
					when "0101000011" => rgb <= "001100";
					when "0101000100" => rgb <= "001100";
					when "0101000101" => rgb <= "001100";
					when "0101000110" => rgb <= "001100";
					when "0101000111" => rgb <= "001100";
					when "0101001000" => rgb <= "001100";
					when "0101001001" => rgb <= "000000";
					when "0101001010" => rgb <= "001100";
					when "0110000000" => rgb <= "001100";
					when "0110000001" => rgb <= "000000";
					when "0110000010" => rgb <= "001100";
					when "0110000011" => rgb <= "000000";
					when "0110000100" => rgb <= "000000";
					when "0110000101" => rgb <= "000000";
					when "0110000110" => rgb <= "000000";
					when "0110000111" => rgb <= "000000";
					when "0110001000" => rgb <= "001100";
					when "0110001001" => rgb <= "000000";
					when "0110001010" => rgb <= "001100";
					when "0111000000" => rgb <= "000000";
					when "0111000001" => rgb <= "000000";
					when "0111000010" => rgb <= "000000";
					when "0111000011" => rgb <= "001100";
					when "0111000100" => rgb <= "001100";
					when "0111000101" => rgb <= "000000";
					when "0111000110" => rgb <= "001100";
					when "0111000111" => rgb <= "001100";
					when "0111001000" => rgb <= "000000";
					when "0111001001" => rgb <= "000000";
					when "0111001010" => rgb <= "000000";
					when others => rgb <= "000000";
                end case;
            end if;
        end process;   
        addr <=  std_logic_vector(yaddr) & std_logic_vector(xaddr);   
    end;
